//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n445, new_n447, new_n451, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n565, new_n566, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n630,
    new_n633, new_n635, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1199, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g023(.A(G452), .Z(G391));
  AND2_X1   g024(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g027(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR4_X1   g032(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  AOI22_X1  g036(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(G319));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OR2_X1    g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(KEYINPUT66), .A3(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n469), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n463), .A2(new_n471), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n472), .A2(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n476), .A2(KEYINPUT67), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n463), .A2(new_n481), .A3(new_n471), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT68), .Z(new_n487));
  INV_X1    g062(.A(G112), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n473), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n471), .B1(new_n466), .B2(new_n467), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n487), .A2(new_n489), .B1(G124), .B2(new_n490), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n485), .A2(new_n491), .ZN(G162));
  NAND4_X1  g067(.A1(new_n465), .A2(G138), .A3(new_n471), .A4(new_n468), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n463), .A2(KEYINPUT4), .A3(G138), .A4(new_n471), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n463), .A2(G126), .A3(G2105), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G114), .C2(new_n471), .ZN(new_n499));
  AND3_X1   g074(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(G75), .A2(G543), .ZN(new_n504));
  XOR2_X1   g079(.A(new_n504), .B(KEYINPUT71), .Z(new_n505));
  OR2_X1    g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n505), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT70), .B1(new_n508), .B2(new_n509), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n503), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n503), .A2(KEYINPUT69), .A3(KEYINPUT6), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n506), .A2(new_n507), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n517), .A2(G651), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n503), .A2(KEYINPUT69), .A3(KEYINPUT6), .ZN(new_n525));
  AOI21_X1  g100(.A(KEYINPUT69), .B1(new_n503), .B2(KEYINPUT6), .ZN(new_n526));
  OAI211_X1 g101(.A(G543), .B(new_n524), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G50), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n522), .A2(new_n523), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n514), .A2(new_n529), .ZN(G166));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XOR2_X1   g106(.A(new_n531), .B(KEYINPUT7), .Z(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n520), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n534), .B2(new_n508), .ZN(new_n535));
  INV_X1    g110(.A(G51), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT72), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n527), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n520), .A2(KEYINPUT72), .A3(G543), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n535), .A2(new_n540), .ZN(G168));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n542), .B1(new_n538), .B2(new_n539), .ZN(new_n543));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n522), .A2(new_n544), .B1(new_n545), .B2(new_n503), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(G171));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n538), .A2(new_n539), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G43), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n520), .A2(G81), .A3(new_n521), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(new_n506), .B2(new_n507), .ZN(new_n553));
  AND2_X1   g128(.A1(G68), .A2(G543), .ZN(new_n554));
  OAI21_X1  g129(.A(G651), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n548), .B1(new_n550), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(G43), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n559), .B1(new_n538), .B2(new_n539), .ZN(new_n560));
  NOR3_X1   g135(.A1(new_n560), .A2(new_n556), .A3(KEYINPUT73), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  XNOR2_X1  g142(.A(KEYINPUT75), .B(G65), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n521), .A2(new_n568), .B1(G78), .B2(G543), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT76), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n503), .B1(new_n569), .B2(new_n570), .ZN(new_n572));
  INV_X1    g147(.A(new_n522), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n571), .A2(new_n572), .B1(G91), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT9), .B1(new_n527), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT9), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n520), .A2(new_n578), .A3(G53), .A4(G543), .ZN(new_n579));
  AND3_X1   g154(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n577), .B1(new_n576), .B2(new_n579), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n574), .B1(new_n580), .B2(new_n581), .ZN(G299));
  INV_X1    g157(.A(G171), .ZN(G301));
  INV_X1    g158(.A(G168), .ZN(G286));
  OR2_X1    g159(.A1(new_n514), .A2(new_n529), .ZN(G303));
  NAND2_X1  g160(.A1(new_n573), .A2(G87), .ZN(new_n586));
  INV_X1    g161(.A(new_n527), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G49), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(G288));
  NAND2_X1  g165(.A1(new_n521), .A2(G61), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n591), .A2(new_n592), .B1(G73), .B2(G543), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n521), .A2(KEYINPUT77), .A3(G61), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n503), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(G48), .B2(new_n587), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n573), .A2(G86), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(KEYINPUT78), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n597), .A2(KEYINPUT78), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(new_n549), .A2(G47), .ZN(new_n601));
  NAND2_X1  g176(.A1(G72), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G60), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n508), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G651), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n573), .A2(G85), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n601), .A2(new_n605), .A3(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n573), .A2(G92), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT79), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n527), .A2(new_n537), .ZN(new_n613));
  AOI21_X1  g188(.A(KEYINPUT72), .B1(new_n520), .B2(G543), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n538), .A2(KEYINPUT79), .A3(new_n539), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n615), .A2(G54), .A3(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n618));
  AND2_X1   g193(.A1(new_n521), .A2(G66), .ZN(new_n619));
  NAND2_X1  g194(.A1(G79), .A2(G543), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT80), .Z(new_n621));
  OAI21_X1  g196(.A(G651), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  AND3_X1   g197(.A1(new_n617), .A2(new_n618), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n618), .B1(new_n617), .B2(new_n622), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n611), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n608), .B1(new_n626), .B2(G868), .ZN(G284));
  OAI21_X1  g202(.A(new_n608), .B1(new_n626), .B2(G868), .ZN(G321));
  NAND2_X1  g203(.A1(G286), .A2(G868), .ZN(new_n629));
  INV_X1    g204(.A(G299), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G868), .ZN(G280));
  XNOR2_X1  g206(.A(G280), .B(KEYINPUT82), .ZN(G297));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n626), .B1(new_n633), .B2(G860), .ZN(G148));
  NOR2_X1   g209(.A1(new_n562), .A2(G868), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n626), .A2(new_n633), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(G868), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT83), .Z(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n490), .A2(G123), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n471), .A2(G111), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  INV_X1    g217(.A(G135), .ZN(new_n643));
  OAI221_X1 g218(.A(new_n640), .B1(new_n641), .B2(new_n642), .C1(new_n483), .C2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT85), .B(G2096), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n469), .A2(new_n474), .A3(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n647), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n465), .A2(new_n468), .ZN(new_n650));
  INV_X1    g225(.A(new_n474), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(KEYINPUT13), .B(G2100), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n646), .A2(new_n655), .ZN(G156));
  INV_X1    g231(.A(KEYINPUT14), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2435), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n661), .B1(new_n660), .B2(new_n659), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2451), .B(G2454), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT16), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1341), .B(G1348), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n662), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2443), .B(G2446), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(G14), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(G401));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT86), .ZN(new_n674));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2072), .B(G2078), .Z(new_n677));
  NOR3_X1   g252(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT18), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n677), .B(KEYINPUT17), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n680), .A2(new_n675), .A3(new_n674), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n675), .B1(new_n674), .B2(new_n677), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n682), .A2(KEYINPUT87), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(KEYINPUT87), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(new_n674), .B2(new_n680), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n679), .B(new_n681), .C1(new_n683), .C2(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G2096), .B(G2100), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G227));
  XNOR2_X1  g263(.A(G1971), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1956), .B(G2474), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT88), .ZN(new_n693));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  NAND3_X1  g269(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT20), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n693), .A2(new_n694), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n693), .A2(new_n694), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n697), .A2(new_n690), .A3(new_n698), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n696), .B(new_n699), .C1(new_n690), .C2(new_n697), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1991), .B(G1996), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(G229));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  NAND2_X1  g282(.A1(G115), .A2(G2104), .ZN(new_n708));
  INV_X1    g283(.A(G127), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n650), .B2(new_n709), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n710), .A2(G2105), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(KEYINPUT92), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(KEYINPUT92), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT91), .B(KEYINPUT25), .Z(new_n714));
  NAND3_X1  g289(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n714), .B(new_n715), .Z(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G139), .B2(new_n484), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n712), .A2(new_n713), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(KEYINPUT93), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT93), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n707), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n707), .B2(G33), .ZN(new_n724));
  OR3_X1    g299(.A1(new_n724), .A2(KEYINPUT94), .A3(new_n442), .ZN(new_n725));
  OAI21_X1  g300(.A(KEYINPUT94), .B1(new_n724), .B2(new_n442), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n484), .A2(G141), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT95), .B(KEYINPUT26), .ZN(new_n728));
  NAND3_X1  g303(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n728), .B(new_n729), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n490), .A2(G129), .ZN(new_n731));
  INV_X1    g306(.A(G105), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n730), .B(new_n731), .C1(new_n732), .C2(new_n651), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n727), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(new_n707), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n707), .B2(G32), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT27), .B(G1996), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT24), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n707), .B1(new_n739), .B2(G34), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n739), .B2(G34), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G160), .B2(G29), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G2084), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n724), .B2(new_n442), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n725), .A2(KEYINPUT96), .A3(new_n726), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n626), .A2(G16), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G4), .B2(G16), .ZN(new_n748));
  INV_X1    g323(.A(G1348), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  INV_X1    g326(.A(G16), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G19), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n562), .B2(new_n752), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(G1341), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n707), .A2(G35), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G162), .B2(new_n707), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT29), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n758), .A2(G2090), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(G2090), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n752), .A2(G21), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G168), .B2(new_n752), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G1966), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n752), .A2(G5), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G171), .B2(new_n752), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n763), .B1(G1961), .B2(new_n765), .ZN(new_n766));
  NOR3_X1   g341(.A1(new_n759), .A2(new_n760), .A3(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G28), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n768), .A2(KEYINPUT30), .ZN(new_n769));
  AOI21_X1  g344(.A(G29), .B1(new_n768), .B2(KEYINPUT30), .ZN(new_n770));
  OR2_X1    g345(.A1(KEYINPUT31), .A2(G11), .ZN(new_n771));
  NAND2_X1  g346(.A1(KEYINPUT31), .A2(G11), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n769), .A2(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n644), .B2(new_n707), .ZN(new_n774));
  NOR2_X1   g349(.A1(G164), .A2(new_n707), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G27), .B2(new_n707), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n774), .B1(new_n776), .B2(new_n443), .ZN(new_n777));
  OAI221_X1 g352(.A(new_n777), .B1(new_n443), .B2(new_n776), .C1(new_n736), .C2(new_n737), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n707), .A2(G26), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT28), .Z(new_n780));
  NAND3_X1  g355(.A1(new_n480), .A2(G140), .A3(new_n482), .ZN(new_n781));
  OAI21_X1  g356(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n782));
  INV_X1    g357(.A(G116), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(G2105), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n490), .B2(G128), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n780), .B1(new_n786), .B2(G29), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G2067), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n742), .B2(G2084), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n765), .A2(G1961), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G1966), .B2(new_n762), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n778), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n752), .A2(G20), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT23), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n630), .B2(new_n752), .ZN(new_n795));
  INV_X1    g370(.A(G1956), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  AND4_X1   g372(.A1(new_n755), .A2(new_n767), .A3(new_n792), .A4(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n746), .A2(new_n750), .A3(new_n751), .A4(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT96), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n725), .A2(new_n726), .A3(new_n745), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n707), .A2(G25), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n484), .A2(G131), .ZN(new_n804));
  OAI21_X1  g379(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n805));
  INV_X1    g380(.A(G107), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(G2105), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n490), .B2(G119), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n803), .B1(new_n810), .B2(new_n707), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT35), .B(G1991), .Z(new_n812));
  XOR2_X1   g387(.A(new_n811), .B(new_n812), .Z(new_n813));
  NOR2_X1   g388(.A1(G16), .A2(G24), .ZN(new_n814));
  XOR2_X1   g389(.A(G290), .B(KEYINPUT89), .Z(new_n815));
  AOI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(G16), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G1986), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT34), .ZN(new_n818));
  NOR2_X1   g393(.A1(G166), .A2(new_n752), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n752), .B2(G22), .ZN(new_n820));
  INV_X1    g395(.A(G1971), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n752), .A2(G23), .ZN(new_n823));
  INV_X1    g398(.A(G288), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n824), .B2(new_n752), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT33), .B(G1976), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n820), .A2(new_n821), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n822), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n752), .A2(G6), .ZN(new_n830));
  INV_X1    g405(.A(G305), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(new_n752), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT32), .B(G1981), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  AOI211_X1 g410(.A(new_n813), .B(new_n817), .C1(new_n818), .C2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT90), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n835), .B2(new_n818), .ZN(new_n838));
  OAI211_X1 g413(.A(KEYINPUT90), .B(KEYINPUT34), .C1(new_n829), .C2(new_n834), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n836), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT36), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT36), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n836), .A2(new_n842), .A3(new_n838), .A4(new_n839), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n802), .A2(KEYINPUT97), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(KEYINPUT97), .B1(new_n802), .B2(new_n844), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(G311));
  NAND2_X1  g422(.A1(new_n802), .A2(new_n844), .ZN(G150));
  INV_X1    g423(.A(G93), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n850));
  OAI22_X1  g425(.A1(new_n522), .A2(new_n849), .B1(new_n850), .B2(new_n503), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(G55), .B2(new_n549), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(new_n558), .B2(new_n561), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n560), .A2(new_n556), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT38), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n626), .A2(G559), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n861));
  AOI21_X1  g436(.A(G860), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(new_n861), .B2(new_n860), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n853), .A2(G860), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT37), .Z(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT98), .ZN(G145));
  INV_X1    g442(.A(new_n786), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n495), .A2(new_n500), .A3(KEYINPUT99), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT99), .B1(new_n495), .B2(new_n500), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n501), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n874), .A2(new_n786), .A3(new_n869), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n727), .A2(new_n733), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT100), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n872), .A2(new_n734), .A3(new_n875), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n721), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n719), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n884));
  AOI22_X1  g459(.A1(new_n879), .A2(new_n722), .B1(new_n878), .B2(new_n880), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n480), .A2(G142), .A3(new_n482), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n890));
  INV_X1    g465(.A(G118), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n890), .B1(new_n891), .B2(G2105), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n892), .B1(new_n490), .B2(G130), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n653), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n648), .A2(new_n652), .A3(new_n889), .A4(new_n893), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n809), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n895), .A2(new_n809), .A3(new_n896), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n888), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  INV_X1    g476(.A(new_n888), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n901), .A2(new_n897), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n718), .B1(new_n881), .B2(new_n721), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT104), .B1(new_n905), .B2(new_n885), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n887), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT105), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n887), .A2(new_n906), .A3(KEYINPUT105), .A4(new_n904), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n883), .A2(new_n886), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n900), .B2(new_n903), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n898), .A2(new_n888), .A3(new_n899), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n902), .B1(new_n901), .B2(new_n897), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(new_n916), .A3(KEYINPUT103), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n912), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g495(.A1(G160), .A2(new_n644), .ZN(new_n921));
  NAND2_X1  g496(.A1(G160), .A2(new_n644), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n921), .A2(G162), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(G162), .B1(new_n921), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT106), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OR3_X1    g500(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT106), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n920), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n911), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n923), .A2(new_n924), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n912), .A2(new_n919), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n918), .B1(new_n883), .B2(new_n886), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(G37), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n929), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g512(.A(new_n636), .B(new_n857), .Z(new_n938));
  INV_X1    g513(.A(KEYINPUT41), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n616), .A2(G54), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT79), .B1(new_n538), .B2(new_n539), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n622), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT81), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n617), .A2(new_n618), .A3(new_n622), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n630), .B1(new_n945), .B2(new_n611), .ZN(new_n946));
  AOI211_X1 g521(.A(G299), .B(new_n610), .C1(new_n943), .C2(new_n944), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n939), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n625), .A2(G299), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n945), .A2(new_n630), .A3(new_n611), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(KEYINPUT41), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n938), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n946), .A2(new_n947), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n953), .B1(new_n954), .B2(new_n938), .ZN(new_n955));
  NAND2_X1  g530(.A1(G166), .A2(KEYINPUT107), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(G166), .A2(KEYINPUT107), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n831), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(G290), .B(G288), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n961));
  NAND2_X1  g536(.A1(G303), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n962), .A2(G305), .A3(new_n956), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n959), .A2(new_n960), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n960), .B1(new_n959), .B2(new_n963), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT42), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n955), .B(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(G868), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(G868), .B2(new_n852), .ZN(G295));
  OAI21_X1  g545(.A(new_n969), .B1(G868), .B2(new_n852), .ZN(G331));
  INV_X1    g546(.A(new_n543), .ZN(new_n972));
  INV_X1    g547(.A(new_n546), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n972), .B(new_n973), .C1(new_n540), .C2(new_n535), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n549), .A2(G51), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n520), .A2(G89), .ZN(new_n976));
  NAND2_X1  g551(.A1(G63), .A2(G651), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n532), .B1(new_n978), .B2(new_n521), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n975), .B(new_n979), .C1(new_n543), .C2(new_n546), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n854), .A2(new_n856), .A3(new_n974), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n974), .A2(new_n980), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n550), .A2(new_n548), .A3(new_n557), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT73), .B1(new_n560), .B2(new_n556), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n852), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n852), .A2(new_n855), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n982), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n981), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n948), .A2(new_n951), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n988), .A2(new_n949), .A3(new_n950), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(new_n966), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n934), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n991), .B(KEYINPUT111), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n948), .A2(new_n951), .A3(KEYINPUT110), .A4(new_n989), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n990), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n994), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n966), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n993), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n1000), .A2(KEYINPUT43), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n990), .A2(new_n991), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n966), .B1(new_n1002), .B2(KEYINPUT108), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT108), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n990), .A2(new_n1004), .A3(new_n991), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n993), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(KEYINPUT43), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT44), .B1(new_n1001), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n998), .A2(new_n999), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n1010));
  INV_X1    g585(.A(new_n993), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT112), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1000), .A2(new_n1014), .A3(new_n1010), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT109), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT109), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n990), .A2(new_n1004), .A3(new_n991), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1004), .B1(new_n990), .B2(new_n991), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1018), .A2(new_n1019), .A3(new_n966), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1017), .B(KEYINPUT43), .C1(new_n1020), .C2(new_n993), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n1013), .A2(new_n1015), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1008), .B1(new_n1022), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g598(.A(KEYINPUT45), .ZN(new_n1024));
  INV_X1    g599(.A(G1384), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n501), .A2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(KEYINPUT113), .B(G40), .ZN(new_n1027));
  AND4_X1   g602(.A1(new_n1024), .A2(G160), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1996), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  XOR2_X1   g607(.A(new_n1032), .B(KEYINPUT125), .Z(new_n1033));
  INV_X1    g608(.A(G2067), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n786), .B(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n734), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1030), .A2(new_n1031), .B1(new_n1028), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1033), .A2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1038), .B(KEYINPUT47), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n734), .B(G1996), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1040), .A2(new_n1035), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n810), .A2(new_n812), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n810), .A2(new_n812), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1044), .A2(new_n1028), .ZN(new_n1045));
  NOR2_X1   g620(.A1(G290), .A2(G1986), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT48), .B1(new_n1028), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1028), .A2(KEYINPUT48), .A3(new_n1046), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1041), .ZN(new_n1050));
  XOR2_X1   g625(.A(new_n1042), .B(KEYINPUT124), .Z(new_n1051));
  OAI22_X1  g626(.A1(new_n1050), .A2(new_n1051), .B1(G2067), .B2(new_n786), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1048), .A2(new_n1049), .B1(new_n1028), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1039), .A2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1054), .B(KEYINPUT126), .ZN(new_n1055));
  OR2_X1    g630(.A1(G305), .A2(G1981), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n596), .A2(new_n597), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G1981), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT49), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1061), .B(KEYINPUT115), .ZN(new_n1062));
  INV_X1    g637(.A(G8), .ZN(new_n1063));
  AND4_X1   g638(.A1(new_n1025), .A2(G160), .A3(new_n501), .A4(new_n1027), .ZN(new_n1064));
  AOI211_X1 g639(.A(new_n1063), .B(new_n1064), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1976), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n824), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1056), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1064), .A2(new_n1063), .ZN(new_n1070));
  AND2_X1   g645(.A1(G160), .A2(new_n1027), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n1026), .A2(KEYINPUT50), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1026), .A2(KEYINPUT50), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G2090), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1026), .B(KEYINPUT45), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1071), .A2(new_n1077), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1075), .A2(new_n1076), .B1(new_n1078), .B2(new_n821), .ZN(new_n1079));
  NAND2_X1  g654(.A1(G303), .A2(G8), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n1080), .B(KEYINPUT55), .ZN(new_n1081));
  OR3_X1    g656(.A1(new_n1079), .A2(new_n1063), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT52), .B1(G288), .B2(new_n1067), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1070), .B(new_n1084), .C1(new_n1067), .C2(G288), .ZN(new_n1085));
  AOI211_X1 g660(.A(new_n1063), .B(new_n1064), .C1(G1976), .C2(new_n824), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT52), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1088), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1069), .A2(new_n1070), .B1(new_n1083), .B2(new_n1089), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1079), .A2(new_n1063), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n1081), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1078), .ZN(new_n1093));
  OAI22_X1  g668(.A1(new_n1093), .A2(G1966), .B1(new_n1074), .B2(G2084), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G8), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1095), .A2(G286), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1089), .A2(new_n1092), .A3(new_n1082), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT63), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1091), .A2(KEYINPUT116), .ZN(new_n1100));
  OR3_X1    g675(.A1(new_n1079), .A2(KEYINPUT116), .A3(new_n1063), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1100), .A2(new_n1081), .A3(new_n1101), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1095), .A2(new_n1098), .A3(G286), .ZN(new_n1103));
  AND4_X1   g678(.A1(new_n1082), .A2(new_n1102), .A3(new_n1089), .A4(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1090), .B1(new_n1099), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1078), .A2(G2078), .ZN(new_n1107));
  OAI22_X1  g682(.A1(new_n1107), .A2(KEYINPUT53), .B1(new_n1075), .B2(G1961), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1107), .A2(KEYINPUT53), .ZN(new_n1109));
  OAI21_X1  g684(.A(G171), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT122), .B(G2078), .Z(new_n1111));
  AND3_X1   g686(.A1(new_n1111), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1077), .A2(G160), .A3(new_n1112), .ZN(new_n1113));
  XOR2_X1   g688(.A(new_n1113), .B(KEYINPUT123), .Z(new_n1114));
  OR2_X1    g689(.A1(new_n1114), .A2(new_n1108), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1110), .B1(new_n1115), .B2(G171), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1106), .B1(new_n1115), .B2(G171), .ZN(new_n1117));
  OR3_X1    g692(.A1(new_n1108), .A2(new_n1109), .A3(G171), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1106), .A2(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n630), .A2(KEYINPUT57), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n576), .A2(new_n579), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n574), .A2(new_n1121), .ZN(new_n1122));
  XOR2_X1   g697(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT56), .B(G2072), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1071), .A2(new_n1077), .A3(new_n1125), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n1126), .A2(KEYINPUT118), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1074), .A2(new_n796), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1126), .A2(KEYINPUT118), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1120), .B(new_n1124), .C1(new_n1129), .C2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1127), .A2(new_n1130), .A3(new_n1128), .A4(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT61), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(KEYINPUT61), .ZN(new_n1136));
  XNOR2_X1  g711(.A(KEYINPUT58), .B(G1341), .ZN(new_n1137));
  OAI22_X1  g712(.A1(new_n1078), .A2(G1996), .B1(new_n1064), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1138), .A2(KEYINPUT59), .A3(new_n562), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1074), .A2(new_n749), .B1(new_n1034), .B2(new_n1064), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT60), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1140), .A2(new_n1141), .A3(new_n626), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1138), .A2(new_n562), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT59), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1136), .A2(new_n1139), .A3(new_n1142), .A4(new_n1145), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n1140), .A2(new_n625), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1140), .A2(new_n625), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1141), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1135), .A2(new_n1146), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1134), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1133), .B(KEYINPUT119), .ZN(new_n1153));
  OAI22_X1  g728(.A1(new_n1151), .A2(new_n1147), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1119), .B1(new_n1150), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1110), .A2(KEYINPUT62), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1094), .A2(KEYINPUT120), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT120), .ZN(new_n1158));
  OAI221_X1 g733(.A(new_n1158), .B1(new_n1074), .B2(G2084), .C1(new_n1093), .C2(G1966), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1157), .A2(new_n1159), .A3(G8), .ZN(new_n1160));
  NAND2_X1  g735(.A1(G286), .A2(G8), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT121), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT51), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT51), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1095), .A2(new_n1165), .A3(new_n1162), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1157), .A2(new_n1159), .A3(new_n1163), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1156), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1155), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1089), .A2(new_n1092), .A3(new_n1082), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1172));
  OAI211_X1 g747(.A(KEYINPUT62), .B(G171), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1105), .B1(new_n1170), .B2(new_n1174), .ZN(new_n1175));
  AND2_X1   g750(.A1(G290), .A2(G1986), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1028), .B1(new_n1046), .B2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT114), .ZN(new_n1178));
  OR2_X1    g753(.A1(new_n1045), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1055), .B1(new_n1175), .B2(new_n1179), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n1182));
  NAND2_X1  g756(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1183));
  NAND2_X1  g757(.A1(new_n1016), .A2(new_n1021), .ZN(new_n1184));
  NAND2_X1  g758(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g759(.A(G319), .B1(new_n670), .B2(new_n671), .ZN(new_n1186));
  OR2_X1    g760(.A1(new_n1186), .A2(G227), .ZN(new_n1187));
  INV_X1    g761(.A(new_n705), .ZN(new_n1188));
  OR2_X1    g762(.A1(new_n704), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g763(.A1(new_n704), .A2(new_n1188), .ZN(new_n1190));
  AOI21_X1  g764(.A(new_n1187), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g765(.A(new_n927), .B1(new_n909), .B2(new_n910), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n933), .A2(new_n934), .ZN(new_n1193));
  OAI21_X1  g767(.A(new_n1191), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g768(.A(new_n1194), .ZN(new_n1195));
  AOI21_X1  g769(.A(new_n1182), .B1(new_n1185), .B2(new_n1195), .ZN(new_n1196));
  AOI211_X1 g770(.A(KEYINPUT127), .B(new_n1194), .C1(new_n1183), .C2(new_n1184), .ZN(new_n1197));
  NOR2_X1   g771(.A1(new_n1196), .A2(new_n1197), .ZN(G308));
  OAI21_X1  g772(.A(KEYINPUT127), .B1(new_n1022), .B2(new_n1194), .ZN(new_n1199));
  NAND3_X1  g773(.A1(new_n1185), .A2(new_n1195), .A3(new_n1182), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n1199), .A2(new_n1200), .ZN(G225));
endmodule


