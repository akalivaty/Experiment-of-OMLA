

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763;

  AND2_X1 U375 ( .A1(n732), .A2(n618), .ZN(n365) );
  OR2_X1 U376 ( .A1(n748), .A2(n370), .ZN(n363) );
  BUF_X1 U377 ( .A(n579), .Z(n594) );
  XNOR2_X1 U378 ( .A(n375), .B(n374), .ZN(n703) );
  XNOR2_X1 U379 ( .A(n398), .B(n397), .ZN(n681) );
  OR2_X1 U380 ( .A1(n703), .A2(n521), .ZN(n373) );
  XNOR2_X1 U381 ( .A(n453), .B(n419), .ZN(n432) );
  XNOR2_X1 U382 ( .A(G131), .B(KEYINPUT4), .ZN(n419) );
  XNOR2_X1 U383 ( .A(G146), .B(G125), .ZN(n479) );
  NAND2_X1 U384 ( .A1(n618), .A2(KEYINPUT2), .ZN(n372) );
  NOR2_X1 U385 ( .A1(n757), .A2(n762), .ZN(n509) );
  AND2_X1 U386 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U387 ( .A1(n662), .A2(n373), .ZN(n528) );
  INV_X1 U388 ( .A(G210), .ZN(n493) );
  XNOR2_X1 U389 ( .A(G128), .B(KEYINPUT24), .ZN(n383) );
  XOR2_X1 U390 ( .A(G137), .B(G140), .Z(n430) );
  INV_X1 U391 ( .A(G902), .ZN(n472) );
  XNOR2_X1 U392 ( .A(n367), .B(n432), .ZN(n631) );
  INV_X1 U393 ( .A(n488), .ZN(n368) );
  XOR2_X1 U394 ( .A(G146), .B(G110), .Z(n434) );
  OR2_X1 U395 ( .A1(n369), .A2(n592), .ZN(n429) );
  XNOR2_X1 U396 ( .A(n379), .B(KEYINPUT41), .ZN(n712) );
  AND2_X1 U397 ( .A1(n698), .A2(n377), .ZN(n379) );
  NOR2_X1 U398 ( .A1(n700), .A2(n378), .ZN(n377) );
  XNOR2_X1 U399 ( .A(n457), .B(n456), .ZN(n458) );
  NOR2_X1 U400 ( .A1(n728), .A2(G902), .ZN(n459) );
  INV_X1 U401 ( .A(KEYINPUT99), .ZN(n456) );
  XNOR2_X1 U402 ( .A(G104), .B(G101), .ZN(n439) );
  XNOR2_X1 U403 ( .A(n471), .B(n470), .ZN(n722) );
  AND2_X1 U404 ( .A1(n544), .A2(n669), .ZN(n375) );
  XNOR2_X1 U405 ( .A(KEYINPUT87), .B(KEYINPUT15), .ZN(n391) );
  NOR2_X1 U406 ( .A1(G902), .A2(G237), .ZN(n492) );
  XNOR2_X1 U407 ( .A(n401), .B(KEYINPUT91), .ZN(n558) );
  XNOR2_X1 U408 ( .A(G146), .B(G119), .ZN(n422) );
  NOR2_X1 U409 ( .A1(G953), .A2(G237), .ZN(n466) );
  AND2_X1 U410 ( .A1(n606), .A2(n605), .ZN(n607) );
  AND2_X1 U411 ( .A1(n604), .A2(KEYINPUT44), .ZN(n606) );
  NOR2_X1 U412 ( .A1(n542), .A2(n353), .ZN(n543) );
  XNOR2_X1 U413 ( .A(n400), .B(n399), .ZN(n405) );
  NAND2_X1 U414 ( .A1(G234), .A2(G237), .ZN(n399) );
  XNOR2_X1 U415 ( .A(KEYINPUT76), .B(KEYINPUT14), .ZN(n400) );
  XNOR2_X1 U416 ( .A(n413), .B(KEYINPUT67), .ZN(n369) );
  AND2_X1 U417 ( .A1(n681), .A2(n412), .ZN(n413) );
  XOR2_X1 U418 ( .A(G113), .B(G116), .Z(n426) );
  XNOR2_X1 U419 ( .A(n390), .B(n389), .ZN(n623) );
  XOR2_X1 U420 ( .A(G116), .B(G107), .Z(n448) );
  INV_X1 U421 ( .A(G953), .ZN(n477) );
  BUF_X1 U422 ( .A(n523), .Z(n549) );
  NAND2_X1 U423 ( .A1(n446), .A2(n355), .ZN(n662) );
  AND2_X1 U424 ( .A1(n573), .A2(n684), .ZN(n600) );
  XNOR2_X1 U425 ( .A(n437), .B(n436), .ZN(n441) );
  XNOR2_X1 U426 ( .A(n501), .B(n500), .ZN(n757) );
  NOR2_X1 U427 ( .A1(n522), .A2(n712), .ZN(n501) );
  AND2_X1 U428 ( .A1(n358), .A2(n666), .ZN(n508) );
  XNOR2_X1 U429 ( .A(n572), .B(n571), .ZN(n648) );
  NAND2_X1 U430 ( .A1(n520), .A2(n530), .ZN(n673) );
  XOR2_X1 U431 ( .A(KEYINPUT74), .B(n541), .Z(n353) );
  AND2_X1 U432 ( .A1(n408), .A2(n559), .ZN(n354) );
  AND2_X1 U433 ( .A1(n527), .A2(n445), .ZN(n355) );
  NOR2_X1 U434 ( .A1(n511), .A2(n369), .ZN(n356) );
  XNOR2_X1 U435 ( .A(n391), .B(n472), .ZN(n617) );
  INV_X1 U436 ( .A(n371), .ZN(n370) );
  NAND2_X1 U437 ( .A1(n372), .A2(n376), .ZN(n371) );
  XNOR2_X2 U438 ( .A(n569), .B(n568), .ZN(n573) );
  XNOR2_X2 U439 ( .A(n616), .B(n615), .ZN(n732) );
  AND2_X1 U440 ( .A1(n358), .A2(n357), .ZN(n545) );
  INV_X1 U441 ( .A(n544), .ZN(n357) );
  XNOR2_X1 U442 ( .A(n506), .B(n359), .ZN(n358) );
  INV_X1 U443 ( .A(KEYINPUT39), .ZN(n359) );
  NAND2_X1 U444 ( .A1(n360), .A2(n748), .ZN(n362) );
  NAND2_X1 U445 ( .A1(n732), .A2(n620), .ZN(n360) );
  AND2_X1 U446 ( .A1(n748), .A2(n732), .ZN(n679) );
  NAND2_X2 U447 ( .A1(n364), .A2(n361), .ZN(n622) );
  NAND2_X1 U448 ( .A1(n363), .A2(n362), .ZN(n361) );
  OR2_X2 U449 ( .A1(n365), .A2(n371), .ZN(n364) );
  XNOR2_X1 U450 ( .A(n366), .B(n368), .ZN(n367) );
  XNOR2_X1 U451 ( .A(n425), .B(n424), .ZN(n366) );
  NAND2_X1 U452 ( .A1(n631), .A2(n472), .ZN(n427) );
  NAND2_X1 U453 ( .A1(n446), .A2(n445), .ZN(n522) );
  INV_X1 U454 ( .A(KEYINPUT101), .ZN(n374) );
  INV_X1 U455 ( .A(KEYINPUT83), .ZN(n376) );
  NAND2_X1 U456 ( .A1(n698), .A2(n697), .ZN(n702) );
  INV_X1 U457 ( .A(n697), .ZN(n378) );
  XNOR2_X2 U458 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n474) );
  BUF_X1 U459 ( .A(n721), .Z(n727) );
  INV_X1 U460 ( .A(n562), .ZN(n527) );
  NOR2_X1 U461 ( .A1(n514), .A2(n685), .ZN(n380) );
  INV_X1 U462 ( .A(KEYINPUT82), .ZN(n535) );
  XNOR2_X1 U463 ( .A(n536), .B(n535), .ZN(n538) );
  AND2_X1 U464 ( .A1(n538), .A2(n537), .ZN(n539) );
  INV_X1 U465 ( .A(KEYINPUT102), .ZN(n403) );
  INV_X1 U466 ( .A(KEYINPUT79), .ZN(n435) );
  XNOR2_X1 U467 ( .A(n435), .B(KEYINPUT92), .ZN(n436) );
  XNOR2_X1 U468 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U469 ( .A(n469), .B(n744), .ZN(n470) );
  BUF_X1 U470 ( .A(n639), .Z(n642) );
  NOR2_X1 U471 ( .A1(n531), .A2(n505), .ZN(n506) );
  XNOR2_X1 U472 ( .A(n497), .B(n496), .ZN(n523) );
  INV_X1 U473 ( .A(n731), .ZN(n635) );
  BUF_X2 U474 ( .A(n477), .Z(n749) );
  NAND2_X1 U475 ( .A1(G234), .A2(n749), .ZN(n381) );
  XOR2_X1 U476 ( .A(KEYINPUT8), .B(n381), .Z(n447) );
  NAND2_X1 U477 ( .A1(G221), .A2(n447), .ZN(n382) );
  XOR2_X2 U478 ( .A(G119), .B(G110), .Z(n485) );
  XNOR2_X1 U479 ( .A(n382), .B(n485), .ZN(n390) );
  XOR2_X1 U480 ( .A(KEYINPUT23), .B(KEYINPUT68), .Z(n384) );
  XNOR2_X1 U481 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U482 ( .A(n430), .B(n385), .ZN(n388) );
  INV_X1 U483 ( .A(KEYINPUT10), .ZN(n386) );
  XNOR2_X1 U484 ( .A(n479), .B(n386), .ZN(n744) );
  INV_X1 U485 ( .A(n744), .ZN(n387) );
  NAND2_X1 U486 ( .A1(n623), .A2(n472), .ZN(n398) );
  XNOR2_X1 U487 ( .A(KEYINPUT25), .B(KEYINPUT93), .ZN(n394) );
  NAND2_X1 U488 ( .A1(n617), .A2(G234), .ZN(n392) );
  XNOR2_X1 U489 ( .A(n392), .B(KEYINPUT20), .ZN(n409) );
  NAND2_X1 U490 ( .A1(n409), .A2(G217), .ZN(n393) );
  XNOR2_X1 U491 ( .A(n394), .B(n393), .ZN(n396) );
  XOR2_X1 U492 ( .A(KEYINPUT78), .B(KEYINPUT94), .Z(n395) );
  XNOR2_X1 U493 ( .A(n396), .B(n395), .ZN(n397) );
  NAND2_X1 U494 ( .A1(n405), .A2(G902), .ZN(n401) );
  NAND2_X1 U495 ( .A1(G953), .A2(n558), .ZN(n402) );
  NOR2_X1 U496 ( .A1(G900), .A2(n402), .ZN(n404) );
  XNOR2_X1 U497 ( .A(n404), .B(n403), .ZN(n408) );
  NAND2_X1 U498 ( .A1(G952), .A2(n405), .ZN(n711) );
  NOR2_X1 U499 ( .A1(G953), .A2(n711), .ZN(n407) );
  INV_X1 U500 ( .A(KEYINPUT90), .ZN(n406) );
  XNOR2_X1 U501 ( .A(n407), .B(n406), .ZN(n559) );
  AND2_X1 U502 ( .A1(n409), .A2(G221), .ZN(n411) );
  INV_X1 U503 ( .A(KEYINPUT21), .ZN(n410) );
  XNOR2_X1 U504 ( .A(n411), .B(n410), .ZN(n680) );
  NOR2_X1 U505 ( .A1(n354), .A2(n680), .ZN(n412) );
  INV_X1 U506 ( .A(G143), .ZN(n414) );
  XNOR2_X1 U507 ( .A(n414), .B(G128), .ZN(n475) );
  INV_X1 U508 ( .A(n475), .ZN(n415) );
  NAND2_X1 U509 ( .A1(G134), .A2(n415), .ZN(n418) );
  INV_X1 U510 ( .A(G134), .ZN(n416) );
  NAND2_X1 U511 ( .A1(n416), .A2(n475), .ZN(n417) );
  NAND2_X1 U512 ( .A1(n418), .A2(n417), .ZN(n453) );
  XOR2_X1 U513 ( .A(KEYINPUT5), .B(KEYINPUT95), .Z(n421) );
  NAND2_X1 U514 ( .A1(n466), .A2(G210), .ZN(n420) );
  XNOR2_X1 U515 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U516 ( .A(G137), .B(G101), .Z(n423) );
  XNOR2_X1 U517 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U518 ( .A(n426), .B(KEYINPUT3), .ZN(n488) );
  XNOR2_X2 U519 ( .A(n427), .B(G472), .ZN(n691) );
  INV_X1 U520 ( .A(n691), .ZN(n592) );
  XNOR2_X1 U521 ( .A(KEYINPUT105), .B(KEYINPUT28), .ZN(n428) );
  XNOR2_X1 U522 ( .A(n429), .B(n428), .ZN(n446) );
  INV_X1 U523 ( .A(n430), .ZN(n431) );
  XNOR2_X1 U524 ( .A(n432), .B(n431), .ZN(n745) );
  NAND2_X1 U525 ( .A1(G227), .A2(n477), .ZN(n433) );
  XNOR2_X1 U526 ( .A(n434), .B(n433), .ZN(n437) );
  XNOR2_X1 U527 ( .A(KEYINPUT88), .B(G107), .ZN(n438) );
  XNOR2_X1 U528 ( .A(n439), .B(n438), .ZN(n738) );
  XNOR2_X1 U529 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n440) );
  XNOR2_X1 U530 ( .A(n738), .B(n440), .ZN(n483) );
  XNOR2_X1 U531 ( .A(n441), .B(n483), .ZN(n442) );
  XNOR2_X1 U532 ( .A(n745), .B(n442), .ZN(n652) );
  NAND2_X1 U533 ( .A1(n652), .A2(n472), .ZN(n444) );
  INV_X1 U534 ( .A(G469), .ZN(n443) );
  XNOR2_X2 U535 ( .A(n444), .B(n443), .ZN(n514) );
  INV_X1 U536 ( .A(n514), .ZN(n445) );
  NAND2_X1 U537 ( .A1(n447), .A2(G217), .ZN(n449) );
  XNOR2_X1 U538 ( .A(n449), .B(n448), .ZN(n455) );
  XOR2_X1 U539 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n451) );
  XNOR2_X1 U540 ( .A(G122), .B(KEYINPUT98), .ZN(n450) );
  XNOR2_X1 U541 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U542 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U543 ( .A(n455), .B(n454), .ZN(n728) );
  INV_X1 U544 ( .A(G478), .ZN(n457) );
  XNOR2_X2 U545 ( .A(n459), .B(n458), .ZN(n530) );
  XOR2_X1 U546 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n461) );
  XNOR2_X1 U547 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n460) );
  XNOR2_X1 U548 ( .A(n461), .B(n460), .ZN(n465) );
  XOR2_X1 U549 ( .A(G140), .B(G122), .Z(n463) );
  XNOR2_X1 U550 ( .A(G113), .B(G131), .ZN(n462) );
  XNOR2_X1 U551 ( .A(n463), .B(n462), .ZN(n464) );
  XOR2_X1 U552 ( .A(n465), .B(n464), .Z(n471) );
  XOR2_X1 U553 ( .A(G143), .B(G104), .Z(n468) );
  NAND2_X1 U554 ( .A1(G214), .A2(n466), .ZN(n467) );
  XNOR2_X1 U555 ( .A(n468), .B(n467), .ZN(n469) );
  NAND2_X1 U556 ( .A1(n722), .A2(n472), .ZN(n519) );
  XOR2_X1 U557 ( .A(KEYINPUT13), .B(G475), .Z(n518) );
  XNOR2_X1 U558 ( .A(n519), .B(n518), .ZN(n529) );
  NOR2_X1 U559 ( .A1(n530), .A2(n529), .ZN(n565) );
  INV_X1 U560 ( .A(n565), .ZN(n700) );
  XNOR2_X2 U561 ( .A(KEYINPUT18), .B(KEYINPUT81), .ZN(n473) );
  XNOR2_X1 U562 ( .A(n474), .B(n473), .ZN(n476) );
  XNOR2_X1 U563 ( .A(n476), .B(n475), .ZN(n482) );
  NAND2_X1 U564 ( .A1(n477), .A2(G224), .ZN(n478) );
  XNOR2_X1 U565 ( .A(n478), .B(KEYINPUT80), .ZN(n480) );
  XNOR2_X1 U566 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U567 ( .A(n482), .B(n481), .ZN(n484) );
  XNOR2_X1 U568 ( .A(n484), .B(n483), .ZN(n490) );
  XNOR2_X1 U569 ( .A(G122), .B(n485), .ZN(n487) );
  XOR2_X1 U570 ( .A(KEYINPUT73), .B(KEYINPUT16), .Z(n486) );
  XNOR2_X1 U571 ( .A(n487), .B(n486), .ZN(n489) );
  XNOR2_X1 U572 ( .A(n489), .B(n488), .ZN(n739) );
  XNOR2_X1 U573 ( .A(n490), .B(n739), .ZN(n639) );
  NAND2_X1 U574 ( .A1(n639), .A2(n617), .ZN(n497) );
  INV_X1 U575 ( .A(KEYINPUT77), .ZN(n491) );
  XNOR2_X1 U576 ( .A(n492), .B(n491), .ZN(n499) );
  OR2_X1 U577 ( .A1(n499), .A2(n493), .ZN(n495) );
  INV_X1 U578 ( .A(KEYINPUT89), .ZN(n494) );
  XNOR2_X1 U579 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U580 ( .A(KEYINPUT38), .B(n549), .Z(n505) );
  INV_X1 U581 ( .A(n505), .ZN(n698) );
  INV_X1 U582 ( .A(G214), .ZN(n498) );
  OR2_X1 U583 ( .A1(n499), .A2(n498), .ZN(n697) );
  XNOR2_X1 U584 ( .A(KEYINPUT106), .B(KEYINPUT42), .ZN(n500) );
  OR2_X1 U585 ( .A1(n680), .A2(n681), .ZN(n685) );
  NAND2_X1 U586 ( .A1(n691), .A2(n697), .ZN(n502) );
  XNOR2_X1 U587 ( .A(KEYINPUT30), .B(n502), .ZN(n503) );
  NOR2_X1 U588 ( .A1(n354), .A2(n503), .ZN(n504) );
  NAND2_X1 U589 ( .A1(n380), .A2(n504), .ZN(n531) );
  INV_X1 U590 ( .A(n530), .ZN(n507) );
  AND2_X1 U591 ( .A1(n507), .A2(n529), .ZN(n666) );
  INV_X1 U592 ( .A(n666), .ZN(n669) );
  XNOR2_X1 U593 ( .A(KEYINPUT40), .B(n508), .ZN(n762) );
  XNOR2_X1 U594 ( .A(n509), .B(KEYINPUT46), .ZN(n517) );
  XNOR2_X1 U595 ( .A(n691), .B(KEYINPUT6), .ZN(n598) );
  INV_X1 U596 ( .A(n598), .ZN(n510) );
  NAND2_X1 U597 ( .A1(n666), .A2(n510), .ZN(n511) );
  AND2_X1 U598 ( .A1(n356), .A2(n697), .ZN(n546) );
  INV_X1 U599 ( .A(n549), .ZN(n533) );
  NAND2_X1 U600 ( .A1(n546), .A2(n533), .ZN(n513) );
  XNOR2_X1 U601 ( .A(KEYINPUT107), .B(KEYINPUT36), .ZN(n512) );
  XNOR2_X1 U602 ( .A(n513), .B(n512), .ZN(n516) );
  XNOR2_X2 U603 ( .A(n514), .B(KEYINPUT1), .ZN(n684) );
  INV_X1 U604 ( .A(KEYINPUT86), .ZN(n515) );
  XNOR2_X1 U605 ( .A(n684), .B(n515), .ZN(n557) );
  NAND2_X1 U606 ( .A1(n516), .A2(n557), .ZN(n675) );
  NAND2_X1 U607 ( .A1(n517), .A2(n675), .ZN(n542) );
  XNOR2_X1 U608 ( .A(KEYINPUT66), .B(KEYINPUT47), .ZN(n521) );
  XOR2_X1 U609 ( .A(n519), .B(n518), .Z(n520) );
  XNOR2_X1 U610 ( .A(KEYINPUT100), .B(n673), .ZN(n544) );
  INV_X1 U611 ( .A(n523), .ZN(n524) );
  NAND2_X1 U612 ( .A1(n524), .A2(n697), .ZN(n526) );
  INV_X1 U613 ( .A(KEYINPUT19), .ZN(n525) );
  XNOR2_X1 U614 ( .A(n526), .B(n525), .ZN(n562) );
  XNOR2_X1 U615 ( .A(n528), .B(KEYINPUT75), .ZN(n540) );
  NAND2_X1 U616 ( .A1(n530), .A2(n529), .ZN(n581) );
  NOR2_X1 U617 ( .A1(n531), .A2(n581), .ZN(n532) );
  NAND2_X1 U618 ( .A1(n533), .A2(n532), .ZN(n638) );
  NAND2_X1 U619 ( .A1(n703), .A2(KEYINPUT47), .ZN(n534) );
  NAND2_X1 U620 ( .A1(n638), .A2(n534), .ZN(n536) );
  NAND2_X1 U621 ( .A1(n662), .A2(KEYINPUT47), .ZN(n537) );
  XNOR2_X1 U622 ( .A(n543), .B(KEYINPUT48), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n545), .B(KEYINPUT108), .ZN(n763) );
  INV_X1 U624 ( .A(n763), .ZN(n553) );
  AND2_X1 U625 ( .A1(n684), .A2(n546), .ZN(n548) );
  XNOR2_X1 U626 ( .A(KEYINPUT103), .B(KEYINPUT43), .ZN(n547) );
  XNOR2_X1 U627 ( .A(n548), .B(n547), .ZN(n550) );
  AND2_X1 U628 ( .A1(n550), .A2(n549), .ZN(n552) );
  INV_X1 U629 ( .A(KEYINPUT104), .ZN(n551) );
  XNOR2_X1 U630 ( .A(n552), .B(n551), .ZN(n758) );
  AND2_X1 U631 ( .A1(n553), .A2(n758), .ZN(n554) );
  AND2_X2 U632 ( .A1(n555), .A2(n554), .ZN(n748) );
  AND2_X1 U633 ( .A1(n598), .A2(n681), .ZN(n556) );
  AND2_X1 U634 ( .A1(n557), .A2(n556), .ZN(n570) );
  NOR2_X1 U635 ( .A1(G898), .A2(n749), .ZN(n740) );
  NAND2_X1 U636 ( .A1(n558), .A2(n740), .ZN(n560) );
  AND2_X1 U637 ( .A1(n560), .A2(n559), .ZN(n561) );
  OR2_X2 U638 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X2 U639 ( .A(n563), .B(KEYINPUT0), .ZN(n579) );
  INV_X1 U640 ( .A(n680), .ZN(n564) );
  NAND2_X1 U641 ( .A1(n565), .A2(n564), .ZN(n566) );
  OR2_X2 U642 ( .A1(n579), .A2(n566), .ZN(n569) );
  XNOR2_X1 U643 ( .A(KEYINPUT72), .B(KEYINPUT22), .ZN(n567) );
  XNOR2_X1 U644 ( .A(n567), .B(KEYINPUT65), .ZN(n568) );
  NAND2_X1 U645 ( .A1(n570), .A2(n573), .ZN(n572) );
  INV_X1 U646 ( .A(KEYINPUT32), .ZN(n571) );
  INV_X1 U647 ( .A(n648), .ZN(n605) );
  INV_X1 U648 ( .A(n681), .ZN(n597) );
  NOR2_X1 U649 ( .A1(n691), .A2(n597), .ZN(n574) );
  NAND2_X1 U650 ( .A1(n600), .A2(n574), .ZN(n604) );
  INV_X1 U651 ( .A(KEYINPUT44), .ZN(n609) );
  AND2_X1 U652 ( .A1(n604), .A2(n609), .ZN(n575) );
  NAND2_X1 U653 ( .A1(n605), .A2(n575), .ZN(n576) );
  INV_X1 U654 ( .A(KEYINPUT85), .ZN(n610) );
  NAND2_X1 U655 ( .A1(n576), .A2(n610), .ZN(n586) );
  OR2_X2 U656 ( .A1(n684), .A2(n685), .ZN(n587) );
  NOR2_X1 U657 ( .A1(n587), .A2(n598), .ZN(n578) );
  XOR2_X1 U658 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n577) );
  XNOR2_X1 U659 ( .A(n578), .B(n577), .ZN(n696) );
  NOR2_X1 U660 ( .A1(n696), .A2(n594), .ZN(n580) );
  XNOR2_X1 U661 ( .A(n580), .B(KEYINPUT34), .ZN(n583) );
  INV_X1 U662 ( .A(n581), .ZN(n582) );
  NAND2_X1 U663 ( .A1(n583), .A2(n582), .ZN(n585) );
  INV_X1 U664 ( .A(KEYINPUT35), .ZN(n584) );
  XNOR2_X2 U665 ( .A(n585), .B(n584), .ZN(n761) );
  NAND2_X1 U666 ( .A1(n586), .A2(n761), .ZN(n603) );
  INV_X1 U667 ( .A(n587), .ZN(n588) );
  AND2_X1 U668 ( .A1(n588), .A2(n691), .ZN(n692) );
  INV_X1 U669 ( .A(n594), .ZN(n589) );
  NAND2_X1 U670 ( .A1(n692), .A2(n589), .ZN(n591) );
  INV_X1 U671 ( .A(KEYINPUT31), .ZN(n590) );
  XNOR2_X1 U672 ( .A(n591), .B(n590), .ZN(n672) );
  NAND2_X1 U673 ( .A1(n380), .A2(n592), .ZN(n593) );
  OR2_X1 U674 ( .A1(n594), .A2(n593), .ZN(n658) );
  NAND2_X1 U675 ( .A1(n672), .A2(n658), .ZN(n596) );
  INV_X1 U676 ( .A(n703), .ZN(n595) );
  NAND2_X1 U677 ( .A1(n596), .A2(n595), .ZN(n601) );
  AND2_X1 U678 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U679 ( .A1(n600), .A2(n599), .ZN(n656) );
  AND2_X1 U680 ( .A1(n601), .A2(n656), .ZN(n602) );
  AND2_X1 U681 ( .A1(n603), .A2(n602), .ZN(n614) );
  OR2_X2 U682 ( .A1(n761), .A2(KEYINPUT85), .ZN(n608) );
  NAND2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U685 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n614), .A2(n613), .ZN(n616) );
  XNOR2_X1 U687 ( .A(KEYINPUT84), .B(KEYINPUT45), .ZN(n615) );
  INV_X1 U688 ( .A(n617), .ZN(n618) );
  NAND2_X1 U689 ( .A1(n618), .A2(KEYINPUT83), .ZN(n619) );
  INV_X1 U690 ( .A(KEYINPUT2), .ZN(n678) );
  NAND2_X1 U691 ( .A1(n619), .A2(n678), .ZN(n620) );
  INV_X1 U692 ( .A(KEYINPUT64), .ZN(n621) );
  XNOR2_X2 U693 ( .A(n622), .B(n621), .ZN(n721) );
  NAND2_X1 U694 ( .A1(n721), .A2(G217), .ZN(n625) );
  XOR2_X1 U695 ( .A(KEYINPUT122), .B(n623), .Z(n624) );
  XNOR2_X1 U696 ( .A(n625), .B(n624), .ZN(n627) );
  INV_X1 U697 ( .A(G952), .ZN(n626) );
  AND2_X1 U698 ( .A1(n626), .A2(G953), .ZN(n731) );
  NOR2_X2 U699 ( .A1(n627), .A2(n731), .ZN(n629) );
  INV_X1 U700 ( .A(KEYINPUT123), .ZN(n628) );
  XNOR2_X1 U701 ( .A(n629), .B(n628), .ZN(G66) );
  NAND2_X1 U702 ( .A1(n721), .A2(G472), .ZN(n633) );
  XNOR2_X1 U703 ( .A(KEYINPUT109), .B(KEYINPUT62), .ZN(n630) );
  XNOR2_X1 U704 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U705 ( .A(n633), .B(n632), .ZN(n634) );
  INV_X1 U706 ( .A(n634), .ZN(n636) );
  NAND2_X1 U707 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U708 ( .A(n637), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U709 ( .A(n638), .B(G143), .ZN(G45) );
  NAND2_X1 U710 ( .A1(n721), .A2(G210), .ZN(n644) );
  XNOR2_X1 U711 ( .A(KEYINPUT118), .B(KEYINPUT54), .ZN(n640) );
  XNOR2_X1 U712 ( .A(n640), .B(KEYINPUT55), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n644), .B(n643), .ZN(n645) );
  NOR2_X2 U715 ( .A1(n645), .A2(n731), .ZN(n647) );
  XOR2_X1 U716 ( .A(KEYINPUT119), .B(KEYINPUT56), .Z(n646) );
  XNOR2_X1 U717 ( .A(n647), .B(n646), .ZN(G51) );
  XNOR2_X1 U718 ( .A(n604), .B(G110), .ZN(G12) );
  XOR2_X1 U719 ( .A(n648), .B(G119), .Z(G21) );
  NAND2_X1 U720 ( .A1(n727), .A2(G469), .ZN(n654) );
  XOR2_X1 U721 ( .A(KEYINPUT121), .B(KEYINPUT57), .Z(n650) );
  XNOR2_X1 U722 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U724 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n654), .B(n653), .ZN(n655) );
  NOR2_X1 U726 ( .A1(n655), .A2(n731), .ZN(G54) );
  XNOR2_X1 U727 ( .A(G101), .B(n656), .ZN(G3) );
  NOR2_X1 U728 ( .A1(n669), .A2(n658), .ZN(n657) );
  XOR2_X1 U729 ( .A(G104), .B(n657), .Z(G6) );
  NOR2_X1 U730 ( .A1(n673), .A2(n658), .ZN(n660) );
  XNOR2_X1 U731 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U733 ( .A(G107), .B(n661), .ZN(G9) );
  XOR2_X1 U734 ( .A(G128), .B(KEYINPUT29), .Z(n665) );
  INV_X1 U735 ( .A(n662), .ZN(n667) );
  INV_X1 U736 ( .A(n673), .ZN(n663) );
  NAND2_X1 U737 ( .A1(n667), .A2(n663), .ZN(n664) );
  XNOR2_X1 U738 ( .A(n665), .B(n664), .ZN(G30) );
  NAND2_X1 U739 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U740 ( .A(n668), .B(G146), .ZN(G48) );
  NOR2_X1 U741 ( .A1(n669), .A2(n672), .ZN(n670) );
  XOR2_X1 U742 ( .A(KEYINPUT110), .B(n670), .Z(n671) );
  XNOR2_X1 U743 ( .A(G113), .B(n671), .ZN(G15) );
  NOR2_X1 U744 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U745 ( .A(G116), .B(n674), .Z(G18) );
  XNOR2_X1 U746 ( .A(KEYINPUT37), .B(KEYINPUT111), .ZN(n676) );
  XNOR2_X1 U747 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U748 ( .A(G125), .B(n677), .ZN(G27) );
  XNOR2_X1 U749 ( .A(n679), .B(n678), .ZN(n717) );
  NAND2_X1 U750 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U751 ( .A(n682), .B(KEYINPUT49), .ZN(n683) );
  XNOR2_X1 U752 ( .A(KEYINPUT113), .B(n683), .ZN(n689) );
  NAND2_X1 U753 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U754 ( .A(n686), .B(KEYINPUT114), .ZN(n687) );
  XNOR2_X1 U755 ( .A(KEYINPUT50), .B(n687), .ZN(n688) );
  NAND2_X1 U756 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U757 ( .A1(n691), .A2(n690), .ZN(n693) );
  NOR2_X1 U758 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U759 ( .A(KEYINPUT51), .B(n694), .Z(n695) );
  NOR2_X1 U760 ( .A1(n712), .A2(n695), .ZN(n708) );
  NOR2_X1 U761 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U762 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U763 ( .A(KEYINPUT115), .B(n701), .Z(n705) );
  NOR2_X1 U764 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U765 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U766 ( .A1(n696), .A2(n706), .ZN(n707) );
  NOR2_X1 U767 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U768 ( .A(n709), .B(KEYINPUT52), .ZN(n710) );
  NOR2_X1 U769 ( .A1(n711), .A2(n710), .ZN(n714) );
  NOR2_X1 U770 ( .A1(n696), .A2(n712), .ZN(n713) );
  NOR2_X1 U771 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U772 ( .A(KEYINPUT116), .B(n715), .Z(n716) );
  NOR2_X1 U773 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U774 ( .A1(n749), .A2(n718), .ZN(n719) );
  XNOR2_X1 U775 ( .A(n719), .B(KEYINPUT53), .ZN(n720) );
  XNOR2_X1 U776 ( .A(KEYINPUT117), .B(n720), .ZN(G75) );
  NAND2_X1 U777 ( .A1(n721), .A2(G475), .ZN(n724) );
  XNOR2_X1 U778 ( .A(n722), .B(KEYINPUT59), .ZN(n723) );
  XNOR2_X1 U779 ( .A(n724), .B(n723), .ZN(n725) );
  NOR2_X2 U780 ( .A1(n725), .A2(n731), .ZN(n726) );
  XNOR2_X1 U781 ( .A(n726), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U782 ( .A1(n727), .A2(G478), .ZN(n729) );
  XNOR2_X1 U783 ( .A(n729), .B(n728), .ZN(n730) );
  NOR2_X1 U784 ( .A1(n731), .A2(n730), .ZN(G63) );
  BUF_X1 U785 ( .A(n732), .Z(n733) );
  NAND2_X1 U786 ( .A1(n733), .A2(n749), .ZN(n737) );
  NAND2_X1 U787 ( .A1(G953), .A2(G224), .ZN(n734) );
  XNOR2_X1 U788 ( .A(KEYINPUT61), .B(n734), .ZN(n735) );
  NAND2_X1 U789 ( .A1(n735), .A2(G898), .ZN(n736) );
  NAND2_X1 U790 ( .A1(n737), .A2(n736), .ZN(n743) );
  XNOR2_X1 U791 ( .A(n739), .B(n738), .ZN(n741) );
  NOR2_X1 U792 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U793 ( .A(n743), .B(n742), .ZN(G69) );
  XNOR2_X1 U794 ( .A(n745), .B(n744), .ZN(n746) );
  XNOR2_X1 U795 ( .A(KEYINPUT124), .B(n746), .ZN(n751) );
  XNOR2_X1 U796 ( .A(KEYINPUT125), .B(n751), .ZN(n747) );
  XNOR2_X1 U797 ( .A(n748), .B(n747), .ZN(n750) );
  NAND2_X1 U798 ( .A1(n750), .A2(n749), .ZN(n755) );
  XNOR2_X1 U799 ( .A(G227), .B(n751), .ZN(n752) );
  NAND2_X1 U800 ( .A1(n752), .A2(G900), .ZN(n753) );
  NAND2_X1 U801 ( .A1(G953), .A2(n753), .ZN(n754) );
  NAND2_X1 U802 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U803 ( .A(KEYINPUT126), .B(n756), .ZN(G72) );
  XOR2_X1 U804 ( .A(G137), .B(n757), .Z(G39) );
  XNOR2_X1 U805 ( .A(G140), .B(n758), .ZN(n759) );
  XNOR2_X1 U806 ( .A(n759), .B(KEYINPUT112), .ZN(G42) );
  XOR2_X1 U807 ( .A(G122), .B(KEYINPUT127), .Z(n760) );
  XNOR2_X1 U808 ( .A(n761), .B(n760), .ZN(G24) );
  XOR2_X1 U809 ( .A(G131), .B(n762), .Z(G33) );
  XOR2_X1 U810 ( .A(G134), .B(n763), .Z(G36) );
endmodule

