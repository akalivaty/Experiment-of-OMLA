

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771;

  NOR2_X1 U375 ( .A1(G953), .A2(G237), .ZN(n513) );
  XNOR2_X1 U376 ( .A(n467), .B(G953), .ZN(n505) );
  NOR2_X1 U377 ( .A1(n553), .A2(n552), .ZN(n359) );
  NAND2_X4 U378 ( .A1(n353), .A2(n352), .ZN(n717) );
  NOR2_X2 U379 ( .A1(n408), .A2(n354), .ZN(n407) );
  XNOR2_X2 U380 ( .A(KEYINPUT3), .B(G119), .ZN(n475) );
  NOR2_X2 U381 ( .A1(n770), .A2(n645), .ZN(n583) );
  XNOR2_X2 U382 ( .A(n389), .B(n364), .ZN(n766) );
  XNOR2_X2 U383 ( .A(n412), .B(n411), .ZN(n738) );
  NOR2_X1 U384 ( .A1(n542), .A2(n768), .ZN(n543) );
  OR2_X1 U385 ( .A1(n579), .A2(KEYINPUT39), .ZN(n425) );
  NAND2_X1 U386 ( .A1(n553), .A2(n551), .ZN(n732) );
  INV_X1 U387 ( .A(n376), .ZN(n367) );
  INV_X1 U388 ( .A(G125), .ZN(n390) );
  XNOR2_X2 U389 ( .A(G110), .B(G104), .ZN(n479) );
  AND2_X1 U390 ( .A1(n378), .A2(n355), .ZN(n418) );
  XNOR2_X1 U391 ( .A(n541), .B(KEYINPUT35), .ZN(n768) );
  XNOR2_X1 U392 ( .A(n442), .B(KEYINPUT34), .ZN(n441) );
  AND2_X1 U393 ( .A1(n386), .A2(n512), .ZN(n354) );
  XNOR2_X1 U394 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U395 ( .A(n461), .B(n460), .ZN(n553) );
  XOR2_X1 U396 ( .A(KEYINPUT59), .B(n653), .Z(n654) );
  XNOR2_X1 U397 ( .A(n520), .B(n477), .ZN(n483) );
  XNOR2_X1 U398 ( .A(n484), .B(KEYINPUT4), .ZN(n503) );
  XNOR2_X1 U399 ( .A(n390), .B(G146), .ZN(n377) );
  AND2_X2 U400 ( .A1(n384), .A2(n598), .ZN(n555) );
  XNOR2_X2 U401 ( .A(n503), .B(n502), .ZN(n403) );
  NAND2_X2 U402 ( .A1(n547), .A2(n500), .ZN(n501) );
  XNOR2_X2 U403 ( .A(n374), .B(n499), .ZN(n547) );
  NOR2_X1 U404 ( .A1(G902), .A2(G237), .ZN(n486) );
  XNOR2_X1 U405 ( .A(G134), .B(G131), .ZN(n502) );
  XNOR2_X1 U406 ( .A(n568), .B(KEYINPUT71), .ZN(n596) );
  NAND2_X1 U407 ( .A1(n635), .A2(G472), .ZN(n401) );
  NAND2_X1 U408 ( .A1(n437), .A2(n431), .ZN(n436) );
  AND2_X1 U409 ( .A1(n588), .A2(KEYINPUT86), .ZN(n393) );
  INV_X1 U410 ( .A(KEYINPUT48), .ZN(n612) );
  XNOR2_X1 U411 ( .A(KEYINPUT73), .B(G469), .ZN(n511) );
  XNOR2_X1 U412 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n421) );
  AND2_X1 U413 ( .A1(n578), .A2(n719), .ZN(n388) );
  INV_X1 U414 ( .A(G472), .ZN(n432) );
  NAND2_X1 U415 ( .A1(G902), .A2(G472), .ZN(n433) );
  XNOR2_X1 U416 ( .A(n403), .B(n402), .ZN(n635) );
  XNOR2_X1 U417 ( .A(n391), .B(G122), .ZN(n476) );
  INV_X1 U418 ( .A(KEYINPUT74), .ZN(n391) );
  NAND2_X1 U419 ( .A1(n524), .A2(G221), .ZN(n382) );
  INV_X1 U420 ( .A(G101), .ZN(n478) );
  INV_X1 U421 ( .A(KEYINPUT33), .ZN(n411) );
  XNOR2_X1 U422 ( .A(n561), .B(n395), .ZN(n747) );
  INV_X1 U423 ( .A(KEYINPUT41), .ZN(n395) );
  OR2_X1 U424 ( .A1(n730), .A2(KEYINPUT39), .ZN(n427) );
  XNOR2_X1 U425 ( .A(KEYINPUT69), .B(KEYINPUT0), .ZN(n499) );
  NOR2_X1 U426 ( .A1(n571), .A2(n570), .ZN(n584) );
  NAND2_X1 U427 ( .A1(n587), .A2(n393), .ZN(n593) );
  INV_X1 U428 ( .A(KEYINPUT92), .ZN(n536) );
  NAND2_X1 U429 ( .A1(n440), .A2(n439), .ZN(n386) );
  NAND2_X1 U430 ( .A1(n511), .A2(G902), .ZN(n439) );
  XNOR2_X1 U431 ( .A(G137), .B(G101), .ZN(n517) );
  INV_X1 U432 ( .A(KEYINPUT5), .ZN(n516) );
  NAND2_X1 U433 ( .A1(G234), .A2(G237), .ZN(n494) );
  INV_X1 U434 ( .A(KEYINPUT90), .ZN(n416) );
  XNOR2_X1 U435 ( .A(n415), .B(n533), .ZN(n714) );
  XNOR2_X1 U436 ( .A(G128), .B(G110), .ZN(n528) );
  XNOR2_X1 U437 ( .A(G140), .B(G137), .ZN(n529) );
  XNOR2_X1 U438 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n526) );
  XNOR2_X1 U439 ( .A(G119), .B(KEYINPUT87), .ZN(n525) );
  XNOR2_X1 U440 ( .A(n468), .B(n414), .ZN(n524) );
  INV_X1 U441 ( .A(KEYINPUT8), .ZN(n414) );
  XNOR2_X1 U442 ( .A(G116), .B(KEYINPUT9), .ZN(n462) );
  XOR2_X1 U443 ( .A(KEYINPUT105), .B(KEYINPUT7), .Z(n463) );
  XNOR2_X1 U444 ( .A(G134), .B(G107), .ZN(n465) );
  XNOR2_X1 U445 ( .A(G113), .B(G143), .ZN(n453) );
  XOR2_X1 U446 ( .A(G131), .B(KEYINPUT12), .Z(n449) );
  XNOR2_X1 U447 ( .A(KEYINPUT77), .B(KEYINPUT98), .ZN(n506) );
  XNOR2_X1 U448 ( .A(n420), .B(n419), .ZN(n485) );
  AND2_X1 U449 ( .A1(n505), .A2(G224), .ZN(n419) );
  XNOR2_X1 U450 ( .A(n377), .B(n421), .ZN(n420) );
  INV_X1 U451 ( .A(n706), .ZN(n404) );
  AND2_X1 U452 ( .A1(n359), .A2(n427), .ZN(n423) );
  NOR2_X2 U453 ( .A1(n738), .A2(n443), .ZN(n442) );
  INV_X1 U454 ( .A(KEYINPUT76), .ZN(n399) );
  NOR2_X1 U455 ( .A1(n410), .A2(n576), .ZN(n577) );
  XNOR2_X1 U456 ( .A(n493), .B(n492), .ZN(n373) );
  INV_X1 U457 ( .A(KEYINPUT22), .ZN(n385) );
  NAND2_X1 U458 ( .A1(n432), .A2(n431), .ZN(n430) );
  XNOR2_X1 U459 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U460 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U461 ( .A(n476), .B(KEYINPUT16), .ZN(n477) );
  AND2_X1 U462 ( .A1(n371), .A2(n405), .ZN(n762) );
  INV_X1 U463 ( .A(G953), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n380), .B(n379), .ZN(n674) );
  XNOR2_X1 U465 ( .A(n382), .B(n381), .ZN(n380) );
  XNOR2_X1 U466 ( .A(n664), .B(n527), .ZN(n379) );
  XNOR2_X1 U467 ( .A(n530), .B(n529), .ZN(n381) );
  AND2_X1 U468 ( .A1(n747), .A2(n584), .ZN(n572) );
  OR2_X1 U469 ( .A1(n635), .A2(n430), .ZN(n352) );
  AND2_X1 U470 ( .A1(n401), .A2(n433), .ZN(n353) );
  AND2_X1 U471 ( .A1(n644), .A2(n630), .ZN(n355) );
  BUF_X1 U472 ( .A(n714), .Z(n397) );
  XNOR2_X1 U473 ( .A(KEYINPUT81), .B(n631), .ZN(n356) );
  XOR2_X2 U474 ( .A(G113), .B(G116), .Z(n357) );
  AND2_X1 U475 ( .A1(n378), .A2(n356), .ZN(n358) );
  AND2_X1 U476 ( .A1(n435), .A2(n409), .ZN(n360) );
  NOR2_X1 U477 ( .A1(n616), .A2(n605), .ZN(n361) );
  AND2_X1 U478 ( .A1(n545), .A2(n522), .ZN(n362) );
  INV_X1 U479 ( .A(G902), .ZN(n431) );
  AND2_X1 U480 ( .A1(n424), .A2(n427), .ZN(n363) );
  INV_X1 U481 ( .A(n512), .ZN(n409) );
  XOR2_X1 U482 ( .A(KEYINPUT32), .B(KEYINPUT78), .Z(n364) );
  NAND2_X1 U483 ( .A1(n626), .A2(n627), .ZN(n365) );
  NAND2_X1 U484 ( .A1(n755), .A2(n376), .ZN(n368) );
  NAND2_X1 U485 ( .A1(n366), .A2(n367), .ZN(n369) );
  NAND2_X1 U486 ( .A1(n368), .A2(n369), .ZN(n383) );
  INV_X1 U487 ( .A(n755), .ZN(n366) );
  XNOR2_X1 U488 ( .A(n485), .B(n503), .ZN(n376) );
  NAND2_X1 U489 ( .A1(n555), .A2(n535), .ZN(n389) );
  BUF_X1 U490 ( .A(n766), .Z(n370) );
  XNOR2_X2 U491 ( .A(n560), .B(KEYINPUT45), .ZN(n371) );
  XNOR2_X1 U492 ( .A(n560), .B(KEYINPUT45), .ZN(n428) );
  NAND2_X1 U493 ( .A1(n579), .A2(n361), .ZN(n607) );
  XNOR2_X1 U494 ( .A(n372), .B(n523), .ZN(n392) );
  NAND2_X1 U495 ( .A1(n384), .A2(n362), .ZN(n372) );
  NAND2_X1 U496 ( .A1(n373), .A2(n498), .ZN(n374) );
  NAND2_X1 U497 ( .A1(n584), .A2(n373), .ZN(n585) );
  NAND2_X1 U498 ( .A1(n383), .A2(n623), .ZN(n375) );
  XNOR2_X2 U499 ( .A(n375), .B(n489), .ZN(n616) );
  XNOR2_X2 U500 ( .A(n483), .B(n482), .ZN(n755) );
  XNOR2_X1 U501 ( .A(n377), .B(KEYINPUT10), .ZN(n664) );
  AND2_X1 U502 ( .A1(n424), .A2(n423), .ZN(n422) );
  NAND2_X1 U503 ( .A1(n579), .A2(n426), .ZN(n424) );
  XNOR2_X2 U504 ( .A(n387), .B(n399), .ZN(n579) );
  NAND2_X1 U505 ( .A1(n378), .A2(n644), .ZN(n400) );
  XNOR2_X2 U506 ( .A(n620), .B(n416), .ZN(n378) );
  NAND2_X1 U507 ( .A1(n674), .A2(n431), .ZN(n415) );
  XNOR2_X1 U508 ( .A(n383), .B(n659), .ZN(n660) );
  XNOR2_X2 U509 ( .A(n501), .B(n385), .ZN(n384) );
  NOR2_X2 U510 ( .A1(n766), .A2(n691), .ZN(n537) );
  AND2_X2 U511 ( .A1(n392), .A2(n397), .ZN(n691) );
  INV_X1 U512 ( .A(n386), .ZN(n438) );
  NAND2_X1 U513 ( .A1(n388), .A2(n577), .ZN(n387) );
  NAND2_X1 U514 ( .A1(n717), .A2(n729), .ZN(n575) );
  NAND2_X2 U515 ( .A1(n407), .A2(n406), .ZN(n720) );
  NAND2_X1 U516 ( .A1(n630), .A2(n365), .ZN(n444) );
  NAND2_X1 U517 ( .A1(n678), .A2(n431), .ZN(n473) );
  XNOR2_X1 U518 ( .A(n470), .B(n471), .ZN(n678) );
  NOR2_X1 U519 ( .A1(n613), .A2(n616), .ZN(n600) );
  NAND2_X1 U520 ( .A1(n524), .A2(G217), .ZN(n469) );
  BUF_X1 U521 ( .A(n505), .Z(n666) );
  XNOR2_X2 U522 ( .A(n357), .B(n475), .ZN(n520) );
  XNOR2_X2 U523 ( .A(n394), .B(KEYINPUT70), .ZN(n719) );
  NOR2_X2 U524 ( .A1(n714), .A2(n713), .ZN(n394) );
  NAND2_X1 U525 ( .A1(n438), .A2(n435), .ZN(n410) );
  XNOR2_X1 U526 ( .A(n396), .B(n612), .ZN(n619) );
  NAND2_X1 U527 ( .A1(n610), .A2(n611), .ZN(n396) );
  XNOR2_X1 U528 ( .A(n398), .B(n569), .ZN(n571) );
  NAND2_X1 U529 ( .A1(n596), .A2(n717), .ZN(n398) );
  NAND2_X1 U530 ( .A1(n696), .A2(n586), .ZN(n587) );
  XNOR2_X2 U531 ( .A(n585), .B(KEYINPUT79), .ZN(n696) );
  NAND2_X1 U532 ( .A1(n371), .A2(n358), .ZN(n711) );
  NAND2_X1 U533 ( .A1(n400), .A2(n706), .ZN(n705) );
  XNOR2_X1 U534 ( .A(n400), .B(n668), .ZN(n667) );
  XNOR2_X1 U535 ( .A(n520), .B(n521), .ZN(n402) );
  XNOR2_X2 U536 ( .A(n403), .B(n529), .ZN(n665) );
  NOR2_X1 U537 ( .A1(n371), .A2(n404), .ZN(n707) );
  NAND2_X1 U538 ( .A1(n360), .A2(n438), .ZN(n406) );
  NOR2_X1 U539 ( .A1(n435), .A2(n409), .ZN(n408) );
  NOR2_X1 U540 ( .A1(n410), .A2(n717), .ZN(n548) );
  XNOR2_X1 U541 ( .A(n410), .B(KEYINPUT110), .ZN(n570) );
  NAND2_X1 U542 ( .A1(n413), .A2(n539), .ZN(n412) );
  XNOR2_X1 U543 ( .A(n538), .B(KEYINPUT107), .ZN(n413) );
  NAND2_X1 U544 ( .A1(n417), .A2(n444), .ZN(n429) );
  NAND2_X1 U545 ( .A1(n428), .A2(n418), .ZN(n417) );
  XNOR2_X2 U546 ( .A(n665), .B(n510), .ZN(n648) );
  INV_X1 U547 ( .A(n504), .ZN(n482) );
  NAND2_X1 U548 ( .A1(n422), .A2(n425), .ZN(n582) );
  NAND2_X1 U549 ( .A1(n363), .A2(n425), .ZN(n622) );
  AND2_X1 U550 ( .A1(n730), .A2(KEYINPUT39), .ZN(n426) );
  NAND2_X1 U551 ( .A1(n429), .A2(n711), .ZN(n632) );
  XNOR2_X2 U552 ( .A(n434), .B(G143), .ZN(n484) );
  XNOR2_X2 U553 ( .A(G128), .B(KEYINPUT80), .ZN(n434) );
  OR2_X1 U554 ( .A1(n648), .A2(n436), .ZN(n435) );
  INV_X1 U555 ( .A(n511), .ZN(n437) );
  NAND2_X1 U556 ( .A1(n648), .A2(n511), .ZN(n440) );
  NAND2_X1 U557 ( .A1(n719), .A2(n720), .ZN(n538) );
  INV_X1 U558 ( .A(n738), .ZN(n746) );
  NAND2_X1 U559 ( .A1(n441), .A2(n540), .ZN(n541) );
  INV_X1 U560 ( .A(n547), .ZN(n443) );
  BUF_X1 U561 ( .A(n673), .Z(n677) );
  XNOR2_X1 U562 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U563 ( .A(n519), .B(n518), .ZN(n521) );
  INV_X1 U564 ( .A(KEYINPUT19), .ZN(n492) );
  XNOR2_X1 U565 ( .A(n457), .B(n456), .ZN(n653) );
  XNOR2_X1 U566 ( .A(n488), .B(n487), .ZN(n489) );
  INV_X1 U567 ( .A(KEYINPUT63), .ZN(n641) );
  INV_X1 U568 ( .A(KEYINPUT66), .ZN(n523) );
  XNOR2_X2 U569 ( .A(G902), .B(KEYINPUT15), .ZN(n623) );
  NAND2_X1 U570 ( .A1(n623), .A2(G234), .ZN(n445) );
  XNOR2_X1 U571 ( .A(n445), .B(KEYINPUT20), .ZN(n446) );
  XNOR2_X1 U572 ( .A(n446), .B(KEYINPUT100), .ZN(n531) );
  NAND2_X1 U573 ( .A1(n531), .A2(G221), .ZN(n447) );
  XNOR2_X1 U574 ( .A(n447), .B(KEYINPUT21), .ZN(n713) );
  NAND2_X1 U575 ( .A1(G214), .A2(n513), .ZN(n448) );
  XNOR2_X1 U576 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U577 ( .A(n450), .B(G140), .Z(n452) );
  XNOR2_X1 U578 ( .A(G104), .B(G122), .ZN(n451) );
  XNOR2_X1 U579 ( .A(n452), .B(n451), .ZN(n457) );
  XOR2_X1 U580 ( .A(KEYINPUT103), .B(KEYINPUT11), .Z(n454) );
  XNOR2_X1 U581 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U582 ( .A(n664), .B(n455), .ZN(n456) );
  NOR2_X1 U583 ( .A1(G902), .A2(n653), .ZN(n461) );
  XNOR2_X1 U584 ( .A(KEYINPUT104), .B(KEYINPUT13), .ZN(n459) );
  INV_X1 U585 ( .A(G475), .ZN(n458) );
  XNOR2_X1 U586 ( .A(n463), .B(n462), .ZN(n464) );
  XOR2_X1 U587 ( .A(n464), .B(G122), .Z(n466) );
  XNOR2_X1 U588 ( .A(n466), .B(n465), .ZN(n471) );
  INV_X2 U589 ( .A(KEYINPUT64), .ZN(n467) );
  NAND2_X1 U590 ( .A1(n505), .A2(G234), .ZN(n468) );
  XNOR2_X1 U591 ( .A(n484), .B(n469), .ZN(n470) );
  INV_X1 U592 ( .A(G478), .ZN(n472) );
  XNOR2_X1 U593 ( .A(n473), .B(n472), .ZN(n551) );
  NOR2_X1 U594 ( .A1(n713), .A2(n732), .ZN(n474) );
  XNOR2_X1 U595 ( .A(KEYINPUT106), .B(n474), .ZN(n500) );
  XNOR2_X1 U596 ( .A(n479), .B(n478), .ZN(n481) );
  XOR2_X1 U597 ( .A(KEYINPUT94), .B(G107), .Z(n480) );
  XNOR2_X1 U598 ( .A(n481), .B(n480), .ZN(n504) );
  XNOR2_X1 U599 ( .A(n486), .B(KEYINPUT75), .ZN(n490) );
  NAND2_X1 U600 ( .A1(n490), .A2(G210), .ZN(n488) );
  INV_X1 U601 ( .A(KEYINPUT95), .ZN(n487) );
  NAND2_X1 U602 ( .A1(G214), .A2(n490), .ZN(n729) );
  INV_X1 U603 ( .A(n729), .ZN(n491) );
  NOR2_X2 U604 ( .A1(n616), .A2(n491), .ZN(n493) );
  XNOR2_X1 U605 ( .A(KEYINPUT14), .B(n494), .ZN(n495) );
  NAND2_X1 U606 ( .A1(G952), .A2(n495), .ZN(n745) );
  NOR2_X1 U607 ( .A1(n745), .A2(G953), .ZN(n565) );
  NAND2_X1 U608 ( .A1(G902), .A2(n495), .ZN(n563) );
  XOR2_X1 U609 ( .A(G898), .B(KEYINPUT96), .Z(n761) );
  NAND2_X1 U610 ( .A1(G953), .A2(n761), .ZN(n757) );
  NOR2_X1 U611 ( .A1(n563), .A2(n757), .ZN(n496) );
  NOR2_X1 U612 ( .A1(n565), .A2(n496), .ZN(n497) );
  XNOR2_X1 U613 ( .A(KEYINPUT97), .B(n497), .ZN(n498) );
  NAND2_X1 U614 ( .A1(n666), .A2(G227), .ZN(n508) );
  XNOR2_X1 U615 ( .A(n506), .B(G146), .ZN(n507) );
  XNOR2_X1 U616 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U617 ( .A(n504), .B(n509), .ZN(n510) );
  XNOR2_X1 U618 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n512) );
  INV_X1 U619 ( .A(n720), .ZN(n545) );
  XOR2_X1 U620 ( .A(G146), .B(KEYINPUT101), .Z(n515) );
  NAND2_X1 U621 ( .A1(n513), .A2(G210), .ZN(n514) );
  XNOR2_X1 U622 ( .A(n515), .B(n514), .ZN(n519) );
  INV_X1 U623 ( .A(n717), .ZN(n522) );
  XNOR2_X1 U624 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U625 ( .A(n528), .B(KEYINPUT99), .ZN(n530) );
  NAND2_X1 U626 ( .A1(n531), .A2(G217), .ZN(n532) );
  XNOR2_X1 U627 ( .A(n532), .B(KEYINPUT25), .ZN(n533) );
  INV_X1 U628 ( .A(n397), .ZN(n534) );
  XOR2_X1 U629 ( .A(n717), .B(KEYINPUT6), .Z(n539) );
  NOR2_X1 U630 ( .A1(n545), .A2(n534), .ZN(n535) );
  XNOR2_X1 U631 ( .A(n537), .B(n536), .ZN(n542) );
  INV_X1 U632 ( .A(n539), .ZN(n598) );
  OR2_X1 U633 ( .A1(n553), .A2(n551), .ZN(n605) );
  INV_X1 U634 ( .A(n605), .ZN(n540) );
  XNOR2_X1 U635 ( .A(n543), .B(KEYINPUT44), .ZN(n559) );
  NAND2_X1 U636 ( .A1(n719), .A2(n717), .ZN(n544) );
  NOR2_X1 U637 ( .A1(n545), .A2(n544), .ZN(n725) );
  NAND2_X1 U638 ( .A1(n547), .A2(n725), .ZN(n546) );
  XNOR2_X1 U639 ( .A(n546), .B(KEYINPUT31), .ZN(n700) );
  NAND2_X1 U640 ( .A1(n548), .A2(n719), .ZN(n549) );
  NOR2_X1 U641 ( .A1(n443), .A2(n549), .ZN(n687) );
  NOR2_X1 U642 ( .A1(n700), .A2(n687), .ZN(n550) );
  XOR2_X1 U643 ( .A(KEYINPUT102), .B(n550), .Z(n554) );
  INV_X1 U644 ( .A(n551), .ZN(n552) );
  AND2_X1 U645 ( .A1(n553), .A2(n552), .ZN(n699) );
  NOR2_X1 U646 ( .A1(n359), .A2(n699), .ZN(n734) );
  INV_X1 U647 ( .A(n734), .ZN(n586) );
  NAND2_X1 U648 ( .A1(n554), .A2(n586), .ZN(n557) );
  XNOR2_X1 U649 ( .A(KEYINPUT91), .B(n555), .ZN(n684) );
  OR2_X1 U650 ( .A1(n720), .A2(n397), .ZN(n683) );
  OR2_X1 U651 ( .A1(n684), .A2(n683), .ZN(n556) );
  AND2_X1 U652 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U653 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U654 ( .A(n616), .B(KEYINPUT38), .ZN(n730) );
  NAND2_X1 U655 ( .A1(n730), .A2(n729), .ZN(n733) );
  NOR2_X1 U656 ( .A1(n733), .A2(n732), .ZN(n561) );
  XOR2_X1 U657 ( .A(KEYINPUT28), .B(KEYINPUT111), .Z(n569) );
  OR2_X1 U658 ( .A1(n666), .A2(G900), .ZN(n562) );
  NOR2_X1 U659 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U660 ( .A1(n565), .A2(n564), .ZN(n576) );
  NOR2_X1 U661 ( .A1(n713), .A2(n576), .ZN(n566) );
  XNOR2_X1 U662 ( .A(KEYINPUT72), .B(n566), .ZN(n567) );
  NAND2_X1 U663 ( .A1(n714), .A2(n567), .ZN(n568) );
  XNOR2_X1 U664 ( .A(n572), .B(KEYINPUT42), .ZN(n770) );
  INV_X1 U665 ( .A(KEYINPUT108), .ZN(n573) );
  XNOR2_X1 U666 ( .A(n573), .B(KEYINPUT30), .ZN(n574) );
  XNOR2_X1 U667 ( .A(n575), .B(n574), .ZN(n578) );
  INV_X1 U668 ( .A(KEYINPUT112), .ZN(n580) );
  XNOR2_X1 U669 ( .A(n580), .B(KEYINPUT40), .ZN(n581) );
  XNOR2_X1 U670 ( .A(n582), .B(n581), .ZN(n645) );
  XNOR2_X1 U671 ( .A(n583), .B(KEYINPUT46), .ZN(n611) );
  NOR2_X1 U672 ( .A1(KEYINPUT85), .A2(KEYINPUT47), .ZN(n588) );
  OR2_X1 U673 ( .A1(n696), .A2(KEYINPUT85), .ZN(n591) );
  NAND2_X1 U674 ( .A1(KEYINPUT86), .A2(n734), .ZN(n589) );
  AND2_X1 U675 ( .A1(n589), .A2(KEYINPUT47), .ZN(n590) );
  NAND2_X1 U676 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U677 ( .A1(n593), .A2(n592), .ZN(n604) );
  NAND2_X1 U678 ( .A1(n696), .A2(KEYINPUT85), .ZN(n595) );
  OR2_X1 U679 ( .A1(KEYINPUT86), .A2(n734), .ZN(n594) );
  AND2_X1 U680 ( .A1(n595), .A2(n594), .ZN(n602) );
  NAND2_X1 U681 ( .A1(n596), .A2(n359), .ZN(n597) );
  NOR2_X1 U682 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U683 ( .A1(n599), .A2(n729), .ZN(n613) );
  XNOR2_X1 U684 ( .A(n600), .B(KEYINPUT36), .ZN(n601) );
  NAND2_X1 U685 ( .A1(n601), .A2(n720), .ZN(n703) );
  AND2_X1 U686 ( .A1(n703), .A2(n602), .ZN(n603) );
  NAND2_X1 U687 ( .A1(n604), .A2(n603), .ZN(n609) );
  INV_X1 U688 ( .A(KEYINPUT109), .ZN(n606) );
  XNOR2_X1 U689 ( .A(n607), .B(n606), .ZN(n767) );
  INV_X1 U690 ( .A(n767), .ZN(n608) );
  NOR2_X1 U691 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U692 ( .A1(n613), .A2(n720), .ZN(n615) );
  INV_X1 U693 ( .A(KEYINPUT43), .ZN(n614) );
  XNOR2_X1 U694 ( .A(n615), .B(n614), .ZN(n617) );
  AND2_X1 U695 ( .A1(n616), .A2(n617), .ZN(n704) );
  INV_X1 U696 ( .A(n704), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n620) );
  INV_X1 U698 ( .A(n699), .ZN(n621) );
  OR2_X1 U699 ( .A1(n622), .A2(n621), .ZN(n644) );
  NAND2_X1 U700 ( .A1(KEYINPUT2), .A2(KEYINPUT68), .ZN(n626) );
  INV_X1 U701 ( .A(n623), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n628), .A2(KEYINPUT2), .ZN(n625) );
  INV_X1 U703 ( .A(KEYINPUT68), .ZN(n624) );
  NAND2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n627) );
  INV_X1 U705 ( .A(n627), .ZN(n629) );
  OR2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n644), .A2(KEYINPUT2), .ZN(n631) );
  XNOR2_X2 U708 ( .A(n632), .B(KEYINPUT65), .ZN(n673) );
  NAND2_X1 U709 ( .A1(n673), .A2(G472), .ZN(n637) );
  XNOR2_X1 U710 ( .A(KEYINPUT93), .B(KEYINPUT113), .ZN(n633) );
  XNOR2_X1 U711 ( .A(n633), .B(KEYINPUT62), .ZN(n634) );
  XNOR2_X1 U712 ( .A(n637), .B(n636), .ZN(n640) );
  INV_X1 U713 ( .A(n666), .ZN(n639) );
  INV_X1 U714 ( .A(G952), .ZN(n638) );
  AND2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n681) );
  NOR2_X2 U716 ( .A1(n640), .A2(n681), .ZN(n642) );
  XNOR2_X1 U717 ( .A(n642), .B(n641), .ZN(G57) );
  XNOR2_X1 U718 ( .A(G134), .B(KEYINPUT116), .ZN(n643) );
  XNOR2_X1 U719 ( .A(n644), .B(n643), .ZN(G36) );
  XOR2_X1 U720 ( .A(n645), .B(G131), .Z(G33) );
  NAND2_X1 U721 ( .A1(n673), .A2(G469), .ZN(n650) );
  XNOR2_X1 U722 ( .A(KEYINPUT121), .B(KEYINPUT57), .ZN(n646) );
  XNOR2_X1 U723 ( .A(n646), .B(KEYINPUT58), .ZN(n647) );
  XNOR2_X1 U724 ( .A(n650), .B(n649), .ZN(n651) );
  NOR2_X2 U725 ( .A1(n651), .A2(n681), .ZN(n652) );
  XNOR2_X1 U726 ( .A(n652), .B(KEYINPUT122), .ZN(G54) );
  NAND2_X1 U727 ( .A1(n673), .A2(G475), .ZN(n655) );
  XNOR2_X1 U728 ( .A(n655), .B(n654), .ZN(n656) );
  NOR2_X2 U729 ( .A1(n656), .A2(n681), .ZN(n657) );
  XNOR2_X1 U730 ( .A(n657), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U731 ( .A1(n673), .A2(G210), .ZN(n661) );
  XOR2_X1 U732 ( .A(KEYINPUT83), .B(KEYINPUT54), .Z(n658) );
  XNOR2_X1 U733 ( .A(n658), .B(KEYINPUT55), .ZN(n659) );
  XNOR2_X1 U734 ( .A(n661), .B(n660), .ZN(n662) );
  NOR2_X2 U735 ( .A1(n662), .A2(n681), .ZN(n663) );
  XNOR2_X1 U736 ( .A(n663), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U737 ( .A(n665), .B(n664), .ZN(n668) );
  NAND2_X1 U738 ( .A1(n667), .A2(n666), .ZN(n672) );
  XNOR2_X1 U739 ( .A(n668), .B(G227), .ZN(n669) );
  NAND2_X1 U740 ( .A1(n669), .A2(G900), .ZN(n670) );
  NAND2_X1 U741 ( .A1(G953), .A2(n670), .ZN(n671) );
  NAND2_X1 U742 ( .A1(n672), .A2(n671), .ZN(G72) );
  NAND2_X1 U743 ( .A1(n677), .A2(G217), .ZN(n675) );
  XOR2_X1 U744 ( .A(n675), .B(n674), .Z(n676) );
  NOR2_X1 U745 ( .A1(n676), .A2(n681), .ZN(G66) );
  NAND2_X1 U746 ( .A1(n677), .A2(G478), .ZN(n680) );
  XNOR2_X1 U747 ( .A(n678), .B(KEYINPUT123), .ZN(n679) );
  XNOR2_X1 U748 ( .A(n680), .B(n679), .ZN(n682) );
  NOR2_X1 U749 ( .A1(n682), .A2(n681), .ZN(G63) );
  NOR2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U751 ( .A(G101), .B(n685), .Z(G3) );
  NAND2_X1 U752 ( .A1(n687), .A2(n359), .ZN(n686) );
  XNOR2_X1 U753 ( .A(n686), .B(G104), .ZN(G6) );
  XOR2_X1 U754 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n689) );
  NAND2_X1 U755 ( .A1(n687), .A2(n699), .ZN(n688) );
  XNOR2_X1 U756 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U757 ( .A(G107), .B(n690), .ZN(G9) );
  XOR2_X1 U758 ( .A(n691), .B(G110), .Z(n692) );
  XNOR2_X1 U759 ( .A(KEYINPUT114), .B(n692), .ZN(G12) );
  XOR2_X1 U760 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n694) );
  NAND2_X1 U761 ( .A1(n699), .A2(n696), .ZN(n693) );
  XNOR2_X1 U762 ( .A(n694), .B(n693), .ZN(n695) );
  XOR2_X1 U763 ( .A(G128), .B(n695), .Z(G30) );
  NAND2_X1 U764 ( .A1(n696), .A2(n359), .ZN(n697) );
  XNOR2_X1 U765 ( .A(n697), .B(G146), .ZN(G48) );
  NAND2_X1 U766 ( .A1(n700), .A2(n359), .ZN(n698) );
  XNOR2_X1 U767 ( .A(n698), .B(G113), .ZN(G15) );
  NAND2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U769 ( .A(n701), .B(G116), .ZN(G18) );
  XOR2_X1 U770 ( .A(G125), .B(KEYINPUT37), .Z(n702) );
  XNOR2_X1 U771 ( .A(n703), .B(n702), .ZN(G27) );
  XOR2_X1 U772 ( .A(G140), .B(n704), .Z(G42) );
  XOR2_X1 U773 ( .A(KEYINPUT2), .B(KEYINPUT84), .Z(n706) );
  XNOR2_X1 U774 ( .A(n705), .B(KEYINPUT89), .ZN(n709) );
  XNOR2_X1 U775 ( .A(n707), .B(KEYINPUT88), .ZN(n708) );
  NOR2_X1 U776 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U777 ( .A(n710), .B(KEYINPUT82), .ZN(n712) );
  NAND2_X1 U778 ( .A1(n712), .A2(n711), .ZN(n752) );
  INV_X1 U779 ( .A(n747), .ZN(n728) );
  NAND2_X1 U780 ( .A1(n397), .A2(n713), .ZN(n715) );
  XNOR2_X1 U781 ( .A(n715), .B(KEYINPUT49), .ZN(n716) );
  NOR2_X1 U782 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U783 ( .A(KEYINPUT117), .B(n718), .ZN(n723) );
  NOR2_X1 U784 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U785 ( .A(n721), .B(KEYINPUT50), .ZN(n722) );
  NOR2_X1 U786 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U787 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U788 ( .A(KEYINPUT51), .B(n726), .Z(n727) );
  NOR2_X1 U789 ( .A1(n728), .A2(n727), .ZN(n741) );
  NOR2_X1 U790 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U791 ( .A1(n732), .A2(n731), .ZN(n737) );
  NOR2_X1 U792 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U793 ( .A(n735), .B(KEYINPUT118), .ZN(n736) );
  NOR2_X1 U794 ( .A1(n737), .A2(n736), .ZN(n739) );
  NOR2_X1 U795 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U796 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U797 ( .A(n742), .B(KEYINPUT119), .Z(n743) );
  XNOR2_X1 U798 ( .A(KEYINPUT52), .B(n743), .ZN(n744) );
  NOR2_X1 U799 ( .A1(n745), .A2(n744), .ZN(n750) );
  NAND2_X1 U800 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U801 ( .A(KEYINPUT120), .B(n748), .Z(n749) );
  NOR2_X1 U802 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U803 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U804 ( .A1(n753), .A2(G953), .ZN(n754) );
  XNOR2_X1 U805 ( .A(n754), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U806 ( .A(n755), .B(KEYINPUT125), .Z(n756) );
  NAND2_X1 U807 ( .A1(n757), .A2(n756), .ZN(n765) );
  XOR2_X1 U808 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n759) );
  NAND2_X1 U809 ( .A1(G224), .A2(G953), .ZN(n758) );
  XNOR2_X1 U810 ( .A(n759), .B(n758), .ZN(n760) );
  NOR2_X1 U811 ( .A1(n761), .A2(n760), .ZN(n763) );
  NOR2_X1 U812 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U813 ( .A(n765), .B(n764), .ZN(G69) );
  XOR2_X1 U814 ( .A(n370), .B(G119), .Z(G21) );
  XNOR2_X1 U815 ( .A(G143), .B(n767), .ZN(G45) );
  XOR2_X1 U816 ( .A(n768), .B(G122), .Z(n769) );
  XNOR2_X1 U817 ( .A(KEYINPUT126), .B(n769), .ZN(G24) );
  XNOR2_X1 U818 ( .A(G137), .B(KEYINPUT127), .ZN(n771) );
  XNOR2_X1 U819 ( .A(n771), .B(n770), .ZN(G39) );
endmodule

