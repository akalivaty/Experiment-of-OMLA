//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n563, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n585, new_n586, new_n587, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n631, new_n634, new_n636, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1170, new_n1171, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  XNOR2_X1  g028(.A(G325), .B(KEYINPUT66), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n459), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n462), .A2(G137), .A3(new_n459), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n468));
  XNOR2_X1  g043(.A(new_n467), .B(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n466), .A2(new_n469), .A3(KEYINPUT68), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n465), .B1(new_n472), .B2(new_n473), .ZN(G160));
  NOR2_X1   g049(.A1(new_n460), .A2(new_n461), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n475), .A2(new_n459), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  OAI211_X1 g058(.A(G138), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT4), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n478), .B2(G126), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G164));
  NAND2_X1  g066(.A1(G75), .A2(G543), .ZN(new_n492));
  INV_X1    g067(.A(G543), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT69), .B1(new_n493), .B2(KEYINPUT5), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT5), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n495), .A2(new_n496), .A3(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n493), .A2(KEYINPUT5), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G62), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n492), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G651), .ZN(new_n503));
  OR2_X1    g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AND3_X1   g081(.A1(new_n498), .A2(new_n499), .A3(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT70), .B(G88), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n493), .B1(new_n504), .B2(new_n505), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n507), .A2(new_n508), .B1(G50), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n503), .A2(new_n510), .A3(KEYINPUT71), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(G166));
  AND2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  OAI21_X1  g092(.A(G543), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT72), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n520));
  OAI211_X1 g095(.A(new_n520), .B(G543), .C1(new_n516), .C2(new_n517), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G51), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n494), .A2(new_n497), .B1(KEYINPUT5), .B2(new_n493), .ZN(new_n524));
  AND2_X1   g099(.A1(G63), .A2(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n524), .A2(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n524), .A2(new_n506), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n523), .B(new_n529), .C1(new_n530), .C2(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  AOI22_X1  g108(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G651), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n538), .B1(new_n519), .B2(new_n521), .ZN(new_n539));
  AND4_X1   g114(.A1(G90), .A2(new_n498), .A3(new_n499), .A4(new_n506), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n520), .B1(new_n506), .B2(G543), .ZN(new_n542));
  INV_X1    g117(.A(new_n521), .ZN(new_n543));
  OAI21_X1  g118(.A(G52), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n524), .A2(G90), .A3(new_n506), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n544), .A2(KEYINPUT73), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n536), .B1(new_n541), .B2(new_n546), .ZN(G171));
  AND2_X1   g122(.A1(G68), .A2(G543), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n548), .B1(new_n524), .B2(G56), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT74), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n549), .A2(new_n550), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n551), .A2(KEYINPUT75), .A3(new_n552), .A4(G651), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT75), .ZN(new_n554));
  OAI21_X1  g129(.A(G651), .B1(new_n549), .B2(new_n550), .ZN(new_n555));
  AOI211_X1 g130(.A(KEYINPUT74), .B(new_n548), .C1(new_n524), .C2(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI22_X1  g132(.A1(G43), .A2(new_n522), .B1(new_n507), .B2(G81), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n553), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(G860), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT76), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT77), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n509), .A2(new_n568), .A3(G53), .ZN(new_n569));
  INV_X1    g144(.A(G53), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT9), .B1(new_n518), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n524), .A2(G91), .A3(new_n506), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n498), .A2(G65), .A3(new_n499), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n535), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NOR3_X1   g152(.A1(new_n574), .A2(KEYINPUT78), .A3(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n507), .A2(G91), .B1(new_n569), .B2(new_n571), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n575), .A2(new_n576), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n579), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n578), .A2(new_n583), .ZN(G299));
  INV_X1    g159(.A(new_n536), .ZN(new_n585));
  NOR3_X1   g160(.A1(new_n539), .A2(new_n540), .A3(new_n537), .ZN(new_n586));
  AOI21_X1  g161(.A(KEYINPUT73), .B1(new_n544), .B2(new_n545), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(G301));
  INV_X1    g163(.A(G166), .ZN(G303));
  NAND2_X1  g164(.A1(new_n507), .A2(G87), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n509), .A2(G49), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G288));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n500), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(G48), .B2(new_n509), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n598));
  INV_X1    g173(.A(G86), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n531), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n531), .A2(new_n599), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(KEYINPUT79), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n597), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT80), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g180(.A1(new_n597), .A2(new_n602), .A3(KEYINPUT80), .A4(new_n600), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(G305));
  NAND2_X1  g183(.A1(new_n522), .A2(G47), .ZN(new_n609));
  INV_X1    g184(.A(G85), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n531), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n612), .A2(new_n535), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(G290));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  INV_X1    g191(.A(G92), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n531), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n507), .A2(KEYINPUT10), .A3(G92), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  INV_X1    g196(.A(G66), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n500), .B2(new_n622), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n623), .A2(G651), .B1(G54), .B2(new_n522), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n626), .B2(G171), .ZN(G284));
  OAI21_X1  g203(.A(new_n627), .B1(new_n626), .B2(G171), .ZN(G321));
  NAND2_X1  g204(.A1(G286), .A2(G868), .ZN(new_n630));
  INV_X1    g205(.A(G299), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(G297));
  OAI21_X1  g207(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(G280));
  AOI21_X1  g208(.A(new_n625), .B1(G559), .B2(new_n560), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT81), .ZN(G148));
  OR2_X1    g210(.A1(new_n625), .A2(G559), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G868), .ZN(new_n637));
  INV_X1    g212(.A(new_n559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(G868), .B2(new_n638), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g215(.A1(new_n459), .A2(G2104), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n462), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT12), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  INV_X1    g220(.A(G2100), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  AOI22_X1  g223(.A1(G123), .A2(new_n478), .B1(new_n476), .B2(G135), .ZN(new_n649));
  OAI21_X1  g224(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT82), .ZN(new_n651));
  INV_X1    g226(.A(G111), .ZN(new_n652));
  AOI22_X1  g227(.A1(new_n650), .A2(new_n651), .B1(new_n652), .B2(G2105), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n651), .B2(new_n650), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(G2096), .Z(new_n656));
  NAND3_X1  g231(.A1(new_n647), .A2(new_n648), .A3(new_n656), .ZN(G156));
  XNOR2_X1  g232(.A(KEYINPUT83), .B(KEYINPUT14), .ZN(new_n658));
  XOR2_X1   g233(.A(KEYINPUT15), .B(G2435), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2438), .ZN(new_n660));
  XOR2_X1   g235(.A(G2427), .B(G2430), .Z(new_n661));
  AOI21_X1  g236(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n660), .B2(new_n661), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2451), .B(G2454), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT16), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1341), .B(G1348), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n663), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2443), .B(G2446), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(G14), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT84), .Z(G401));
  XNOR2_X1  g248(.A(G2072), .B(G2078), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT17), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  XOR2_X1   g251(.A(G2084), .B(G2090), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n675), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT87), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(new_n676), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT85), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n676), .B1(new_n682), .B2(new_n674), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(new_n682), .B2(new_n674), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n681), .A2(new_n684), .A3(new_n678), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT86), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n677), .A2(new_n674), .A3(new_n676), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT18), .Z(new_n688));
  NAND3_X1  g263(.A1(new_n680), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G2096), .B(G2100), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(G227));
  XOR2_X1   g266(.A(G1971), .B(G1976), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  XOR2_X1   g268(.A(G1956), .B(G2474), .Z(new_n694));
  XOR2_X1   g269(.A(G1961), .B(G1966), .Z(new_n695));
  AND2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT20), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n694), .A2(new_n695), .ZN(new_n699));
  NOR3_X1   g274(.A1(new_n693), .A2(new_n696), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n693), .B2(new_n699), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(G1991), .B(G1996), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT88), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1981), .B(G1986), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(G229));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G23), .ZN(new_n711));
  INV_X1    g286(.A(G288), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(new_n710), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT33), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G1976), .ZN(new_n715));
  NAND2_X1  g290(.A1(G305), .A2(G16), .ZN(new_n716));
  INV_X1    g291(.A(G6), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n717), .B2(G16), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT32), .B(G1981), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n719), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n716), .B(new_n721), .C1(new_n717), .C2(G16), .ZN(new_n722));
  AND3_X1   g297(.A1(new_n715), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT93), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT90), .B(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(G166), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G22), .B2(new_n725), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(KEYINPUT92), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(KEYINPUT92), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n728), .A2(G1971), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G1971), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n727), .A2(KEYINPUT92), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n727), .A2(KEYINPUT92), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n723), .A2(new_n724), .A3(new_n730), .A4(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n730), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n715), .A2(new_n720), .A3(new_n722), .ZN(new_n737));
  OAI21_X1  g312(.A(KEYINPUT93), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT34), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n735), .A2(KEYINPUT34), .A3(new_n738), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n476), .A2(G131), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n478), .A2(G119), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n459), .A2(G107), .ZN(new_n745));
  OAI21_X1  g320(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n743), .B(new_n744), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT89), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  MUX2_X1   g326(.A(G25), .B(new_n751), .S(G29), .Z(new_n752));
  XOR2_X1   g327(.A(KEYINPUT35), .B(G1991), .Z(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n752), .B(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n725), .A2(G24), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n614), .B2(new_n725), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT91), .B(G1986), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n741), .A2(new_n742), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n762));
  OR2_X1    g337(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n762), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n741), .A2(new_n765), .A3(new_n742), .A4(new_n760), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT97), .B(KEYINPUT28), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT98), .ZN(new_n768));
  INV_X1    g343(.A(G29), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G26), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n768), .B(new_n770), .Z(new_n771));
  AOI22_X1  g346(.A1(G128), .A2(new_n478), .B1(new_n476), .B2(G140), .ZN(new_n772));
  OAI21_X1  g347(.A(KEYINPUT96), .B1(G104), .B2(G2105), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  NOR3_X1   g349(.A1(KEYINPUT96), .A2(G104), .A3(G2105), .ZN(new_n775));
  OAI221_X1 g350(.A(G2104), .B1(G116), .B2(new_n459), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n771), .B1(G29), .B2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G2067), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n769), .A2(G32), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n478), .A2(G129), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n642), .A2(G105), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G141), .B2(new_n476), .ZN(new_n785));
  NAND3_X1  g360(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT101), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT26), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n781), .B1(new_n789), .B2(G29), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT27), .B(G1996), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n769), .A2(G27), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G164), .B2(new_n769), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(G2078), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT100), .B(KEYINPUT24), .ZN(new_n797));
  AOI21_X1  g372(.A(G29), .B1(new_n797), .B2(G34), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G34), .B2(new_n797), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G160), .B2(new_n769), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G2084), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n790), .A2(new_n791), .ZN(new_n802));
  NOR4_X1   g377(.A1(new_n780), .A2(new_n796), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(G20), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n725), .A2(new_n804), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT23), .Z(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n631), .B2(new_n710), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(G1956), .Z(new_n808));
  XOR2_X1   g383(.A(KEYINPUT31), .B(G11), .Z(new_n809));
  NOR2_X1   g384(.A1(new_n655), .A2(new_n769), .ZN(new_n810));
  INV_X1    g385(.A(G28), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(KEYINPUT30), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT102), .Z(new_n813));
  AOI21_X1  g388(.A(G29), .B1(new_n811), .B2(KEYINPUT30), .ZN(new_n814));
  AOI211_X1 g389(.A(new_n809), .B(new_n810), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n769), .A2(G33), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n817), .A2(new_n459), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(KEYINPUT99), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(KEYINPUT99), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT25), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G139), .B2(new_n476), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n819), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n816), .B1(new_n824), .B2(G29), .ZN(new_n825));
  INV_X1    g400(.A(G2072), .ZN(new_n826));
  OAI221_X1 g401(.A(new_n815), .B1(G2078), .B2(new_n794), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n769), .A2(G35), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G162), .B2(new_n769), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT29), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n710), .A2(G21), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(G168), .B2(new_n710), .ZN(new_n832));
  OAI22_X1  g407(.A1(new_n830), .A2(G2090), .B1(G1966), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n827), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n803), .A2(new_n808), .A3(new_n834), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n832), .A2(G1966), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n825), .A2(new_n826), .ZN(new_n837));
  AOI211_X1 g412(.A(new_n836), .B(new_n837), .C1(G2090), .C2(new_n830), .ZN(new_n838));
  NOR2_X1   g413(.A1(G4), .A2(G16), .ZN(new_n839));
  INV_X1    g414(.A(new_n625), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n839), .B1(new_n840), .B2(G16), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT95), .B(G1348), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n710), .A2(G5), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(G171), .B2(new_n710), .ZN(new_n845));
  INV_X1    g420(.A(G1961), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n838), .A2(new_n843), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n725), .A2(G19), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(new_n638), .B2(new_n725), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(G1341), .ZN(new_n851));
  NOR3_X1   g426(.A1(new_n835), .A2(new_n848), .A3(new_n851), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n764), .A2(new_n766), .A3(new_n852), .ZN(G311));
  NAND3_X1  g428(.A1(new_n764), .A2(new_n766), .A3(new_n852), .ZN(G150));
  NAND2_X1  g429(.A1(new_n522), .A2(G55), .ZN(new_n855));
  XOR2_X1   g430(.A(KEYINPUT103), .B(G93), .Z(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n531), .B2(new_n856), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n858), .A2(new_n535), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(G860), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT37), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n840), .A2(G559), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT38), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n559), .A2(new_n861), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n860), .A2(new_n553), .A3(new_n557), .A4(new_n558), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n865), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT104), .Z(new_n872));
  AOI21_X1  g447(.A(G860), .B1(new_n869), .B2(new_n870), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n863), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n874), .B(KEYINPUT105), .Z(G145));
  INV_X1    g450(.A(KEYINPUT107), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n824), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n789), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n751), .B(new_n644), .Z(new_n879));
  OR2_X1    g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n881));
  INV_X1    g456(.A(G118), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n881), .B1(new_n882), .B2(G2105), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n478), .A2(G130), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n884), .B(KEYINPUT108), .Z(new_n885));
  AOI211_X1 g460(.A(new_n883), .B(new_n885), .C1(G142), .C2(new_n476), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n777), .B(new_n490), .Z(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n878), .A2(new_n879), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n880), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n888), .B1(new_n880), .B2(new_n889), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(G160), .B(KEYINPUT106), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n482), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n655), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(G37), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  NOR3_X1   g473(.A1(new_n893), .A2(KEYINPUT109), .A3(new_n897), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT109), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n900), .B1(new_n892), .B2(new_n896), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n898), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g478(.A1(new_n861), .A2(new_n626), .ZN(new_n904));
  XOR2_X1   g479(.A(new_n868), .B(new_n636), .Z(new_n905));
  OAI21_X1  g480(.A(new_n625), .B1(new_n578), .B2(new_n583), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT78), .B1(new_n574), .B2(new_n577), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n580), .A2(new_n582), .A3(new_n579), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n907), .A2(new_n908), .A3(new_n620), .A4(new_n624), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n910), .B(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n905), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n910), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n913), .B1(new_n905), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(KEYINPUT111), .A2(KEYINPUT42), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n915), .B(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n918));
  XNOR2_X1  g493(.A(G288), .B(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n607), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n605), .A3(new_n606), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(G166), .A2(new_n614), .ZN(new_n924));
  NAND3_X1  g499(.A1(G290), .A2(new_n514), .A3(new_n513), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n921), .A2(new_n925), .A3(new_n924), .A4(new_n922), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n929), .B1(KEYINPUT111), .B2(KEYINPUT42), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n917), .B(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n904), .B1(new_n931), .B2(new_n626), .ZN(G295));
  OAI21_X1  g507(.A(new_n904), .B1(new_n931), .B2(new_n626), .ZN(G331));
  AND2_X1   g508(.A1(new_n927), .A2(new_n928), .ZN(new_n934));
  OAI211_X1 g509(.A(KEYINPUT112), .B(new_n585), .C1(new_n586), .C2(new_n587), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(G168), .ZN(new_n936));
  NOR2_X1   g511(.A1(G171), .A2(KEYINPUT112), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT112), .ZN(new_n939));
  NAND3_X1  g514(.A1(G301), .A2(new_n939), .A3(G286), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n868), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(G286), .B1(G171), .B2(KEYINPUT112), .ZN(new_n943));
  NAND2_X1  g518(.A1(G301), .A2(new_n939), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n945), .A2(new_n866), .A3(new_n867), .A4(new_n940), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n942), .A2(new_n910), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n914), .A2(KEYINPUT41), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n910), .A2(new_n911), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n942), .A2(new_n946), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n934), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  AND4_X1   g526(.A1(new_n866), .A2(new_n945), .A3(new_n867), .A4(new_n940), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n945), .A2(new_n940), .B1(new_n866), .B2(new_n867), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n912), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n942), .A2(new_n910), .A3(new_n946), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(new_n929), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  INV_X1    g532(.A(G37), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n951), .A2(new_n956), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT114), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n956), .A2(new_n958), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n954), .A2(new_n955), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n929), .B1(new_n962), .B2(KEYINPUT113), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT113), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n954), .A2(new_n964), .A3(new_n955), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n961), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n960), .B1(new_n966), .B2(new_n957), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT113), .B1(new_n947), .B2(new_n950), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n968), .A2(new_n934), .A3(new_n965), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n947), .A2(new_n950), .ZN(new_n970));
  AOI21_X1  g545(.A(G37), .B1(new_n970), .B2(new_n929), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n972), .A2(KEYINPUT114), .A3(KEYINPUT43), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT44), .B1(new_n967), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n972), .A2(new_n957), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n971), .A2(KEYINPUT43), .A3(new_n951), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT115), .B1(new_n974), .B2(new_n978), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n972), .A2(KEYINPUT43), .B1(KEYINPUT114), .B2(new_n959), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT114), .ZN(new_n981));
  AOI211_X1 g556(.A(new_n981), .B(new_n957), .C1(new_n969), .C2(new_n971), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n975), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n976), .A2(new_n977), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT44), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n983), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n979), .A2(new_n987), .ZN(G397));
  AOI21_X1  g563(.A(G1384), .B1(new_n485), .B2(new_n489), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n465), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n466), .A2(new_n469), .A3(KEYINPUT68), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT68), .B1(new_n466), .B2(new_n469), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n993), .B(G40), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1996), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n789), .B(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n777), .B(new_n779), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n751), .A2(new_n754), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n751), .A2(new_n754), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  XOR2_X1   g580(.A(new_n614), .B(G1986), .Z(new_n1006));
  OAI21_X1  g581(.A(new_n997), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT62), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n989), .A2(KEYINPUT45), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n992), .A2(new_n1009), .A3(G160), .A4(G40), .ZN(new_n1010));
  INV_X1    g585(.A(G1966), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n989), .A2(new_n1013), .ZN(new_n1014));
  AOI211_X1 g589(.A(KEYINPUT50), .B(G1384), .C1(new_n485), .C2(new_n489), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1014), .A2(new_n1015), .A3(new_n996), .ZN(new_n1016));
  INV_X1    g591(.A(G2084), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1012), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(G286), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1012), .A2(new_n1018), .A3(G168), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1020), .A2(KEYINPUT51), .A3(G8), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(G8), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT123), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1022), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1026), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1008), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1010), .A2(new_n1011), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT51), .B1(new_n1030), .B2(G168), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(new_n1023), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT51), .B1(new_n1021), .B2(G8), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT123), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1022), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(KEYINPUT62), .A3(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1014), .A2(new_n996), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1015), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n989), .A2(KEYINPUT45), .ZN(new_n1040));
  AOI211_X1 g615(.A(new_n991), .B(G1384), .C1(new_n485), .C2(new_n489), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1040), .A2(new_n1041), .A3(new_n996), .ZN(new_n1042));
  OAI22_X1  g617(.A1(new_n1039), .A2(G2090), .B1(new_n1042), .B2(G1971), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n1044));
  INV_X1    g619(.A(G8), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1044), .B1(G166), .B2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n513), .A2(KEYINPUT55), .A3(G8), .A4(new_n514), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1043), .A2(G8), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1048), .B1(new_n1043), .B2(G8), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n1052));
  NAND3_X1  g627(.A1(G160), .A2(G40), .A3(new_n989), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n712), .A2(G1976), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(G8), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT52), .ZN(new_n1056));
  INV_X1    g631(.A(G1976), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT52), .B1(G288), .B2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1053), .A2(G8), .A3(new_n1054), .A4(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G1981), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n597), .A2(new_n602), .A3(new_n1061), .A4(new_n600), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n509), .A2(G48), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n524), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(new_n1064), .B2(new_n535), .ZN(new_n1065));
  OAI21_X1  g640(.A(G1981), .B1(new_n1065), .B2(new_n601), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1062), .A2(KEYINPUT49), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1053), .A2(G8), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT49), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1052), .B1(new_n1060), .B2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n1067), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1074), .A2(KEYINPUT116), .A3(new_n1056), .A4(new_n1059), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT124), .B1(new_n1010), .B2(G2078), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT53), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n1079));
  OAI211_X1 g654(.A(KEYINPUT124), .B(new_n1079), .C1(new_n1010), .C2(G2078), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1039), .A2(new_n846), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  AND4_X1   g657(.A1(G171), .A2(new_n1051), .A3(new_n1076), .A4(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1029), .A2(new_n1036), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT125), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT56), .B(G2072), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1042), .A2(new_n1087), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT118), .B(G1956), .Z(new_n1089));
  OAI21_X1  g664(.A(new_n1088), .B1(new_n1016), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(new_n574), .B2(new_n577), .ZN(new_n1092));
  NOR2_X1   g667(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1093), .B(KEYINPUT120), .ZN(new_n1094));
  XOR2_X1   g669(.A(new_n1092), .B(new_n1094), .Z(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1090), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n1010), .B2(G1996), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1042), .A2(KEYINPUT121), .A3(new_n998), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1053), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT58), .B(G1341), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1099), .B(new_n1100), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1103), .A2(new_n1104), .A3(new_n638), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1104), .B1(new_n1103), .B2(new_n638), .ZN(new_n1106));
  INV_X1    g681(.A(G1348), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1039), .A2(new_n1107), .B1(new_n779), .B2(new_n1101), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1108), .A2(new_n625), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1088), .B(new_n1095), .C1(new_n1016), .C2(new_n1089), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1105), .A2(new_n1106), .A3(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n625), .B(KEYINPUT60), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1108), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1110), .B(new_n1116), .C1(new_n625), .C2(new_n1108), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1115), .B1(new_n1109), .B2(KEYINPUT60), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1114), .B(new_n1117), .C1(new_n1118), .C2(new_n1110), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1097), .B1(new_n1112), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1082), .A2(G171), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1078), .A2(G301), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1121), .A2(KEYINPUT54), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT54), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1051), .A2(new_n1076), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1120), .A2(new_n1125), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1029), .A2(new_n1036), .A3(KEYINPUT125), .A4(new_n1083), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1086), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT117), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1030), .A2(new_n1045), .A3(G286), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1051), .A2(new_n1076), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT63), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1060), .A2(new_n1071), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1051), .A2(KEYINPUT63), .A3(new_n1132), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1049), .A2(new_n1136), .ZN(new_n1139));
  NOR2_X1   g714(.A1(G288), .A2(G1976), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1062), .B1(new_n1071), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1142), .A2(G8), .A3(new_n1053), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1131), .B1(new_n1138), .B2(new_n1145), .ZN(new_n1146));
  AOI211_X1 g721(.A(KEYINPUT117), .B(new_n1144), .C1(new_n1135), .C2(new_n1137), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1007), .B1(new_n1130), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1000), .A2(new_n785), .A3(new_n788), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n997), .ZN(new_n1151));
  XOR2_X1   g726(.A(new_n1151), .B(KEYINPUT126), .Z(new_n1152));
  NAND2_X1  g727(.A1(new_n997), .A2(new_n998), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT46), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT127), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1156), .A2(KEYINPUT47), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(KEYINPUT47), .ZN(new_n1158));
  INV_X1    g733(.A(new_n997), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n772), .A2(new_n779), .A3(new_n776), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1159), .A2(G1986), .A3(G290), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1005), .A2(new_n997), .B1(KEYINPUT48), .B2(new_n1163), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n1163), .A2(KEYINPUT48), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1162), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1157), .A2(new_n1158), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1149), .A2(new_n1167), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g743(.A1(new_n672), .A2(G319), .ZN(new_n1170));
  NOR3_X1   g744(.A1(G229), .A2(G227), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g745(.A1(new_n902), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g746(.A1(new_n980), .A2(new_n982), .ZN(new_n1173));
  NOR2_X1   g747(.A1(new_n1172), .A2(new_n1173), .ZN(G308));
  OR2_X1    g748(.A1(new_n1172), .A2(new_n1173), .ZN(G225));
endmodule


