

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U553 ( .A(n753), .B(KEYINPUT100), .ZN(n807) );
  AND2_X2 U554 ( .A1(n562), .A2(n561), .ZN(G164) );
  XOR2_X2 U555 ( .A(KEYINPUT67), .B(n572), .Z(n573) );
  INV_X2 U556 ( .A(G2105), .ZN(n555) );
  NOR2_X1 U557 ( .A1(G2104), .A2(G2105), .ZN(n553) );
  AND2_X1 U558 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U559 ( .A1(n730), .A2(n729), .ZN(n732) );
  NAND2_X1 U560 ( .A1(G160), .A2(n693), .ZN(n723) );
  AND2_X2 U561 ( .A1(G160), .A2(n693), .ZN(n691) );
  NOR2_X1 U562 ( .A1(G164), .A2(G1384), .ZN(n690) );
  XNOR2_X1 U563 ( .A(n567), .B(KEYINPUT65), .ZN(n569) );
  BUF_X1 U564 ( .A(n563), .Z(n564) );
  XOR2_X1 U565 ( .A(KEYINPUT17), .B(n553), .Z(n563) );
  AND2_X2 U566 ( .A1(G2104), .A2(G2105), .ZN(n865) );
  AND2_X2 U567 ( .A1(n766), .A2(G40), .ZN(n693) );
  NOR2_X1 U568 ( .A1(G543), .A2(G651), .ZN(n649) );
  XNOR2_X1 U569 ( .A(KEYINPUT66), .B(KEYINPUT23), .ZN(n568) );
  XOR2_X1 U570 ( .A(KEYINPUT29), .B(n719), .Z(n517) );
  NOR2_X1 U571 ( .A1(n757), .A2(n808), .ZN(n518) );
  AND2_X1 U572 ( .A1(n817), .A2(n786), .ZN(n519) );
  NOR2_X4 U573 ( .A1(n574), .A2(n573), .ZN(G160) );
  AND2_X1 U574 ( .A1(n811), .A2(n810), .ZN(n520) );
  OR2_X1 U575 ( .A1(n978), .A2(n705), .ZN(n521) );
  AND2_X1 U576 ( .A1(n700), .A2(n699), .ZN(n522) );
  INV_X1 U577 ( .A(KEYINPUT99), .ZN(n741) );
  XNOR2_X1 U578 ( .A(n742), .B(n741), .ZN(n743) );
  INV_X1 U579 ( .A(n989), .ZN(n761) );
  INV_X1 U580 ( .A(KEYINPUT13), .ZN(n583) );
  XOR2_X1 U581 ( .A(G543), .B(KEYINPUT0), .Z(n627) );
  NOR2_X1 U582 ( .A1(G651), .A2(n627), .ZN(n650) );
  NOR2_X2 U583 ( .A1(G2104), .A2(n555), .ZN(n864) );
  XOR2_X1 U584 ( .A(KEYINPUT68), .B(n524), .Z(n657) );
  NAND2_X1 U585 ( .A1(n649), .A2(G89), .ZN(n523) );
  XNOR2_X1 U586 ( .A(n523), .B(KEYINPUT4), .ZN(n526) );
  INV_X1 U587 ( .A(G651), .ZN(n528) );
  OR2_X1 U588 ( .A1(n528), .A2(n627), .ZN(n524) );
  NAND2_X1 U589 ( .A1(G76), .A2(n657), .ZN(n525) );
  NAND2_X1 U590 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n527), .B(KEYINPUT5), .ZN(n535) );
  NAND2_X1 U592 ( .A1(G51), .A2(n650), .ZN(n532) );
  NOR2_X1 U593 ( .A1(G543), .A2(n528), .ZN(n530) );
  XNOR2_X1 U594 ( .A(KEYINPUT69), .B(KEYINPUT1), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n530), .B(n529), .ZN(n653) );
  NAND2_X1 U596 ( .A1(G63), .A2(n653), .ZN(n531) );
  NAND2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U598 ( .A(KEYINPUT6), .B(n533), .Z(n534) );
  NAND2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n536), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U601 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U602 ( .A1(G53), .A2(n650), .ZN(n538) );
  NAND2_X1 U603 ( .A1(G65), .A2(n653), .ZN(n537) );
  NAND2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U605 ( .A(KEYINPUT73), .B(n539), .ZN(n543) );
  NAND2_X1 U606 ( .A1(n657), .A2(G78), .ZN(n541) );
  NAND2_X1 U607 ( .A1(G91), .A2(n649), .ZN(n540) );
  AND2_X1 U608 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U609 ( .A1(n543), .A2(n542), .ZN(G299) );
  NAND2_X1 U610 ( .A1(n653), .A2(G64), .ZN(n544) );
  XOR2_X1 U611 ( .A(KEYINPUT71), .B(n544), .Z(n546) );
  NAND2_X1 U612 ( .A1(n650), .A2(G52), .ZN(n545) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(KEYINPUT72), .B(n547), .ZN(n552) );
  NAND2_X1 U615 ( .A1(G90), .A2(n649), .ZN(n549) );
  NAND2_X1 U616 ( .A1(G77), .A2(n657), .ZN(n548) );
  NAND2_X1 U617 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U618 ( .A(KEYINPUT9), .B(n550), .Z(n551) );
  NOR2_X1 U619 ( .A1(n552), .A2(n551), .ZN(G171) );
  AND2_X1 U620 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U621 ( .A(G132), .ZN(G219) );
  INV_X1 U622 ( .A(G82), .ZN(G220) );
  NAND2_X1 U623 ( .A1(G138), .A2(n563), .ZN(n554) );
  XNOR2_X1 U624 ( .A(n554), .B(KEYINPUT90), .ZN(n562) );
  AND2_X4 U625 ( .A1(n555), .A2(G2104), .ZN(n861) );
  NAND2_X1 U626 ( .A1(G102), .A2(n861), .ZN(n557) );
  NAND2_X1 U627 ( .A1(G126), .A2(n864), .ZN(n556) );
  NAND2_X1 U628 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U629 ( .A1(G114), .A2(n865), .ZN(n558) );
  XNOR2_X1 U630 ( .A(KEYINPUT89), .B(n558), .ZN(n559) );
  NOR2_X1 U631 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U632 ( .A1(n564), .A2(G137), .ZN(n566) );
  NAND2_X1 U633 ( .A1(n865), .A2(G113), .ZN(n565) );
  NAND2_X1 U634 ( .A1(n566), .A2(n565), .ZN(n574) );
  NAND2_X1 U635 ( .A1(G101), .A2(n861), .ZN(n567) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n571) );
  NAND2_X1 U637 ( .A1(G125), .A2(n864), .ZN(n570) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U639 ( .A(KEYINPUT10), .B(KEYINPUT75), .Z(n576) );
  NAND2_X1 U640 ( .A1(G7), .A2(G661), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G223) );
  INV_X1 U642 ( .A(G223), .ZN(n834) );
  NAND2_X1 U643 ( .A1(n834), .A2(G567), .ZN(n577) );
  XOR2_X1 U644 ( .A(KEYINPUT11), .B(n577), .Z(G234) );
  XOR2_X1 U645 ( .A(KEYINPUT14), .B(KEYINPUT76), .Z(n579) );
  NAND2_X1 U646 ( .A1(G56), .A2(n653), .ZN(n578) );
  XNOR2_X1 U647 ( .A(n579), .B(n578), .ZN(n586) );
  NAND2_X1 U648 ( .A1(G68), .A2(n657), .ZN(n582) );
  NAND2_X1 U649 ( .A1(n649), .A2(G81), .ZN(n580) );
  XNOR2_X1 U650 ( .A(n580), .B(KEYINPUT12), .ZN(n581) );
  NAND2_X1 U651 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U652 ( .A(n584), .B(n583), .ZN(n585) );
  NOR2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U654 ( .A1(n650), .A2(G43), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n993) );
  INV_X1 U656 ( .A(G860), .ZN(n602) );
  OR2_X1 U657 ( .A1(n993), .A2(n602), .ZN(G153) );
  XNOR2_X1 U658 ( .A(G171), .B(KEYINPUT77), .ZN(G301) );
  NAND2_X1 U659 ( .A1(G868), .A2(G301), .ZN(n598) );
  NAND2_X1 U660 ( .A1(G54), .A2(n650), .ZN(n590) );
  NAND2_X1 U661 ( .A1(G79), .A2(n657), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n595) );
  NAND2_X1 U663 ( .A1(G92), .A2(n649), .ZN(n592) );
  NAND2_X1 U664 ( .A1(G66), .A2(n653), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U666 ( .A(KEYINPUT78), .B(n593), .ZN(n594) );
  NOR2_X1 U667 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U668 ( .A(n596), .B(KEYINPUT15), .ZN(n978) );
  INV_X1 U669 ( .A(G868), .ZN(n671) );
  NAND2_X1 U670 ( .A1(n978), .A2(n671), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n598), .A2(n597), .ZN(G284) );
  NOR2_X1 U672 ( .A1(G286), .A2(n671), .ZN(n599) );
  XOR2_X1 U673 ( .A(KEYINPUT79), .B(n599), .Z(n601) );
  NOR2_X1 U674 ( .A1(G868), .A2(G299), .ZN(n600) );
  NOR2_X1 U675 ( .A1(n601), .A2(n600), .ZN(G297) );
  NAND2_X1 U676 ( .A1(n602), .A2(G559), .ZN(n603) );
  INV_X1 U677 ( .A(n978), .ZN(n617) );
  NAND2_X1 U678 ( .A1(n603), .A2(n617), .ZN(n604) );
  XNOR2_X1 U679 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U680 ( .A1(G868), .A2(n993), .ZN(n607) );
  NAND2_X1 U681 ( .A1(G868), .A2(n617), .ZN(n605) );
  NOR2_X1 U682 ( .A1(G559), .A2(n605), .ZN(n606) );
  NOR2_X1 U683 ( .A1(n607), .A2(n606), .ZN(G282) );
  NAND2_X1 U684 ( .A1(n864), .A2(G123), .ZN(n608) );
  XNOR2_X1 U685 ( .A(n608), .B(KEYINPUT18), .ZN(n610) );
  NAND2_X1 U686 ( .A1(G111), .A2(n865), .ZN(n609) );
  NAND2_X1 U687 ( .A1(n610), .A2(n609), .ZN(n614) );
  NAND2_X1 U688 ( .A1(G99), .A2(n861), .ZN(n612) );
  NAND2_X1 U689 ( .A1(G135), .A2(n564), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n951) );
  XNOR2_X1 U692 ( .A(n951), .B(G2096), .ZN(n616) );
  INV_X1 U693 ( .A(G2100), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n616), .A2(n615), .ZN(G156) );
  NAND2_X1 U695 ( .A1(n617), .A2(G559), .ZN(n669) );
  XNOR2_X1 U696 ( .A(n993), .B(n669), .ZN(n618) );
  NOR2_X1 U697 ( .A1(n618), .A2(G860), .ZN(n626) );
  NAND2_X1 U698 ( .A1(G93), .A2(n649), .ZN(n620) );
  NAND2_X1 U699 ( .A1(G55), .A2(n650), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n625) );
  NAND2_X1 U701 ( .A1(G67), .A2(n653), .ZN(n621) );
  XNOR2_X1 U702 ( .A(n621), .B(KEYINPUT80), .ZN(n623) );
  NAND2_X1 U703 ( .A1(G80), .A2(n657), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n623), .A2(n622), .ZN(n624) );
  OR2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n672) );
  XOR2_X1 U706 ( .A(n626), .B(n672), .Z(G145) );
  NAND2_X1 U707 ( .A1(G87), .A2(n627), .ZN(n629) );
  NAND2_X1 U708 ( .A1(G74), .A2(G651), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U710 ( .A1(n653), .A2(n630), .ZN(n633) );
  NAND2_X1 U711 ( .A1(G49), .A2(n650), .ZN(n631) );
  XOR2_X1 U712 ( .A(KEYINPUT81), .B(n631), .Z(n632) );
  NAND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(G288) );
  NAND2_X1 U714 ( .A1(n657), .A2(G73), .ZN(n634) );
  XNOR2_X1 U715 ( .A(n634), .B(KEYINPUT2), .ZN(n641) );
  NAND2_X1 U716 ( .A1(G48), .A2(n650), .ZN(n636) );
  NAND2_X1 U717 ( .A1(G61), .A2(n653), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U719 ( .A1(n649), .A2(G86), .ZN(n637) );
  XOR2_X1 U720 ( .A(KEYINPUT82), .B(n637), .Z(n638) );
  NOR2_X1 U721 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U722 ( .A1(n641), .A2(n640), .ZN(G305) );
  NAND2_X1 U723 ( .A1(n653), .A2(G62), .ZN(n644) );
  NAND2_X1 U724 ( .A1(n657), .A2(G75), .ZN(n642) );
  XOR2_X1 U725 ( .A(KEYINPUT83), .B(n642), .Z(n643) );
  NAND2_X1 U726 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U727 ( .A1(G88), .A2(n649), .ZN(n646) );
  NAND2_X1 U728 ( .A1(G50), .A2(n650), .ZN(n645) );
  NAND2_X1 U729 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U730 ( .A1(n648), .A2(n647), .ZN(G166) );
  INV_X1 U731 ( .A(G166), .ZN(G303) );
  NAND2_X1 U732 ( .A1(G85), .A2(n649), .ZN(n652) );
  NAND2_X1 U733 ( .A1(G47), .A2(n650), .ZN(n651) );
  NAND2_X1 U734 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U735 ( .A1(n653), .A2(G60), .ZN(n654) );
  XOR2_X1 U736 ( .A(KEYINPUT70), .B(n654), .Z(n655) );
  NOR2_X1 U737 ( .A1(n656), .A2(n655), .ZN(n659) );
  NAND2_X1 U738 ( .A1(G72), .A2(n657), .ZN(n658) );
  NAND2_X1 U739 ( .A1(n659), .A2(n658), .ZN(G290) );
  XNOR2_X1 U740 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n661) );
  INV_X1 U741 ( .A(G299), .ZN(n994) );
  XNOR2_X1 U742 ( .A(G288), .B(n994), .ZN(n660) );
  XNOR2_X1 U743 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U744 ( .A(KEYINPUT86), .B(n662), .ZN(n664) );
  XNOR2_X1 U745 ( .A(n993), .B(KEYINPUT19), .ZN(n663) );
  XNOR2_X1 U746 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U747 ( .A(n665), .B(G305), .ZN(n666) );
  XNOR2_X1 U748 ( .A(n666), .B(G303), .ZN(n667) );
  XOR2_X1 U749 ( .A(n672), .B(n667), .Z(n668) );
  XNOR2_X1 U750 ( .A(n668), .B(G290), .ZN(n881) );
  XNOR2_X1 U751 ( .A(n669), .B(n881), .ZN(n670) );
  NAND2_X1 U752 ( .A1(n670), .A2(G868), .ZN(n674) );
  NAND2_X1 U753 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U754 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2078), .A2(G2084), .ZN(n675) );
  XNOR2_X1 U756 ( .A(n675), .B(KEYINPUT87), .ZN(n676) );
  XNOR2_X1 U757 ( .A(n676), .B(KEYINPUT20), .ZN(n677) );
  NAND2_X1 U758 ( .A1(n677), .A2(G2090), .ZN(n678) );
  XNOR2_X1 U759 ( .A(KEYINPUT21), .B(n678), .ZN(n679) );
  NAND2_X1 U760 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XOR2_X1 U761 ( .A(KEYINPUT74), .B(G57), .Z(G237) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U763 ( .A1(G108), .A2(G120), .ZN(n680) );
  NOR2_X1 U764 ( .A1(G237), .A2(n680), .ZN(n681) );
  NAND2_X1 U765 ( .A1(G69), .A2(n681), .ZN(n838) );
  NAND2_X1 U766 ( .A1(G567), .A2(n838), .ZN(n686) );
  NOR2_X1 U767 ( .A1(G220), .A2(G219), .ZN(n682) );
  XOR2_X1 U768 ( .A(KEYINPUT22), .B(n682), .Z(n683) );
  NOR2_X1 U769 ( .A1(G218), .A2(n683), .ZN(n684) );
  NAND2_X1 U770 ( .A1(G96), .A2(n684), .ZN(n839) );
  NAND2_X1 U771 ( .A1(G2106), .A2(n839), .ZN(n685) );
  NAND2_X1 U772 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U773 ( .A(KEYINPUT88), .B(n687), .Z(G319) );
  INV_X1 U774 ( .A(G319), .ZN(n922) );
  NAND2_X1 U775 ( .A1(G661), .A2(G483), .ZN(n688) );
  NOR2_X1 U776 ( .A1(n922), .A2(n688), .ZN(n837) );
  NAND2_X1 U777 ( .A1(n837), .A2(G36), .ZN(G176) );
  XNOR2_X1 U778 ( .A(n690), .B(KEYINPUT64), .ZN(n766) );
  NAND2_X1 U779 ( .A1(G1996), .A2(n691), .ZN(n692) );
  XNOR2_X1 U780 ( .A(n692), .B(KEYINPUT26), .ZN(n695) );
  INV_X1 U781 ( .A(G1341), .ZN(n1011) );
  NOR2_X1 U782 ( .A1(n691), .A2(n1011), .ZN(n694) );
  NAND2_X1 U783 ( .A1(KEYINPUT26), .A2(n694), .ZN(n698) );
  NAND2_X1 U784 ( .A1(n695), .A2(n698), .ZN(n697) );
  INV_X1 U785 ( .A(KEYINPUT97), .ZN(n696) );
  NAND2_X1 U786 ( .A1(n697), .A2(n696), .ZN(n700) );
  NAND2_X1 U787 ( .A1(n698), .A2(KEYINPUT97), .ZN(n699) );
  INV_X1 U788 ( .A(n993), .ZN(n701) );
  NAND2_X1 U789 ( .A1(n522), .A2(n701), .ZN(n704) );
  NAND2_X1 U790 ( .A1(G1348), .A2(n723), .ZN(n703) );
  NAND2_X1 U791 ( .A1(G2067), .A2(n691), .ZN(n702) );
  NAND2_X1 U792 ( .A1(n703), .A2(n702), .ZN(n705) );
  NAND2_X1 U793 ( .A1(n704), .A2(n521), .ZN(n707) );
  NAND2_X1 U794 ( .A1(n978), .A2(n705), .ZN(n706) );
  NAND2_X1 U795 ( .A1(n707), .A2(n706), .ZN(n713) );
  NAND2_X1 U796 ( .A1(n691), .A2(G2072), .ZN(n708) );
  XNOR2_X1 U797 ( .A(KEYINPUT27), .B(n708), .ZN(n711) );
  NAND2_X1 U798 ( .A1(G1956), .A2(n723), .ZN(n709) );
  XOR2_X1 U799 ( .A(KEYINPUT96), .B(n709), .Z(n710) );
  NOR2_X1 U800 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U801 ( .A1(n994), .A2(n714), .ZN(n712) );
  NAND2_X1 U802 ( .A1(n713), .A2(n712), .ZN(n718) );
  NOR2_X1 U803 ( .A1(n994), .A2(n714), .ZN(n716) );
  INV_X1 U804 ( .A(KEYINPUT28), .ZN(n715) );
  XNOR2_X1 U805 ( .A(n716), .B(n715), .ZN(n717) );
  NAND2_X1 U806 ( .A1(n718), .A2(n717), .ZN(n719) );
  INV_X1 U807 ( .A(n691), .ZN(n735) );
  XNOR2_X1 U808 ( .A(KEYINPUT25), .B(G2078), .ZN(n928) );
  NOR2_X1 U809 ( .A1(n735), .A2(n928), .ZN(n721) );
  AND2_X1 U810 ( .A1(n735), .A2(G1961), .ZN(n720) );
  NOR2_X1 U811 ( .A1(n721), .A2(n720), .ZN(n728) );
  NAND2_X1 U812 ( .A1(G171), .A2(n728), .ZN(n722) );
  NAND2_X1 U813 ( .A1(n517), .A2(n722), .ZN(n734) );
  NAND2_X2 U814 ( .A1(n723), .A2(G8), .ZN(n808) );
  NOR2_X1 U815 ( .A1(G1966), .A2(n808), .ZN(n748) );
  NOR2_X1 U816 ( .A1(G2084), .A2(n723), .ZN(n745) );
  NOR2_X1 U817 ( .A1(n748), .A2(n745), .ZN(n724) );
  NAND2_X1 U818 ( .A1(G8), .A2(n724), .ZN(n725) );
  XNOR2_X1 U819 ( .A(n725), .B(KEYINPUT30), .ZN(n726) );
  XNOR2_X1 U820 ( .A(n726), .B(KEYINPUT98), .ZN(n727) );
  NOR2_X1 U821 ( .A1(n727), .A2(G168), .ZN(n730) );
  NOR2_X1 U822 ( .A1(G171), .A2(n728), .ZN(n729) );
  INV_X1 U823 ( .A(KEYINPUT31), .ZN(n731) );
  XNOR2_X1 U824 ( .A(n732), .B(n731), .ZN(n733) );
  NAND2_X1 U825 ( .A1(n734), .A2(n733), .ZN(n749) );
  NAND2_X1 U826 ( .A1(n749), .A2(G286), .ZN(n740) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n808), .ZN(n737) );
  NOR2_X1 U828 ( .A1(G2090), .A2(n735), .ZN(n736) );
  NOR2_X1 U829 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U830 ( .A1(n738), .A2(G303), .ZN(n739) );
  NAND2_X1 U831 ( .A1(n740), .A2(n739), .ZN(n742) );
  NAND2_X1 U832 ( .A1(n743), .A2(G8), .ZN(n744) );
  XNOR2_X1 U833 ( .A(n744), .B(KEYINPUT32), .ZN(n752) );
  NAND2_X1 U834 ( .A1(G8), .A2(n745), .ZN(n746) );
  XNOR2_X1 U835 ( .A(KEYINPUT95), .B(n746), .ZN(n747) );
  NOR2_X1 U836 ( .A1(n748), .A2(n747), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U838 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n763) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n754) );
  NOR2_X1 U841 ( .A1(n763), .A2(n754), .ZN(n982) );
  INV_X1 U842 ( .A(KEYINPUT33), .ZN(n755) );
  AND2_X1 U843 ( .A1(n982), .A2(n755), .ZN(n756) );
  NAND2_X1 U844 ( .A1(n807), .A2(n756), .ZN(n759) );
  NAND2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n981) );
  INV_X1 U846 ( .A(n981), .ZN(n757) );
  OR2_X1 U847 ( .A1(KEYINPUT33), .A2(n518), .ZN(n758) );
  NAND2_X1 U848 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U849 ( .A(n760), .B(KEYINPUT101), .ZN(n762) );
  XNOR2_X1 U850 ( .A(G1981), .B(G305), .ZN(n989) );
  AND2_X1 U851 ( .A1(n762), .A2(n761), .ZN(n799) );
  INV_X1 U852 ( .A(n808), .ZN(n765) );
  AND2_X1 U853 ( .A1(n763), .A2(KEYINPUT33), .ZN(n764) );
  NAND2_X1 U854 ( .A1(n765), .A2(n764), .ZN(n787) );
  NAND2_X1 U855 ( .A1(G160), .A2(G40), .ZN(n767) );
  NOR2_X1 U856 ( .A1(n767), .A2(n766), .ZN(n829) );
  XOR2_X1 U857 ( .A(KEYINPUT92), .B(KEYINPUT38), .Z(n769) );
  NAND2_X1 U858 ( .A1(G105), .A2(n861), .ZN(n768) );
  XNOR2_X1 U859 ( .A(n769), .B(n768), .ZN(n773) );
  NAND2_X1 U860 ( .A1(G117), .A2(n865), .ZN(n771) );
  NAND2_X1 U861 ( .A1(G141), .A2(n564), .ZN(n770) );
  NAND2_X1 U862 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n775) );
  NAND2_X1 U864 ( .A1(n864), .A2(G129), .ZN(n774) );
  NAND2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n856) );
  NAND2_X1 U866 ( .A1(G1996), .A2(n856), .ZN(n784) );
  NAND2_X1 U867 ( .A1(G119), .A2(n864), .ZN(n777) );
  NAND2_X1 U868 ( .A1(G107), .A2(n865), .ZN(n776) );
  NAND2_X1 U869 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U870 ( .A(KEYINPUT91), .B(n778), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n861), .A2(G95), .ZN(n780) );
  NAND2_X1 U872 ( .A1(G131), .A2(n564), .ZN(n779) );
  AND2_X1 U873 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n875) );
  NAND2_X1 U875 ( .A1(G1991), .A2(n875), .ZN(n783) );
  NAND2_X1 U876 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U877 ( .A(KEYINPUT93), .B(n785), .Z(n952) );
  NAND2_X1 U878 ( .A1(n829), .A2(n952), .ZN(n817) );
  XNOR2_X1 U879 ( .A(G1986), .B(G290), .ZN(n998) );
  NAND2_X1 U880 ( .A1(n829), .A2(n998), .ZN(n786) );
  AND2_X1 U881 ( .A1(n787), .A2(n519), .ZN(n797) );
  NAND2_X1 U882 ( .A1(G104), .A2(n861), .ZN(n789) );
  NAND2_X1 U883 ( .A1(G140), .A2(n564), .ZN(n788) );
  NAND2_X1 U884 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U885 ( .A(KEYINPUT34), .B(n790), .ZN(n795) );
  NAND2_X1 U886 ( .A1(G128), .A2(n864), .ZN(n792) );
  NAND2_X1 U887 ( .A1(G116), .A2(n865), .ZN(n791) );
  NAND2_X1 U888 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U889 ( .A(KEYINPUT35), .B(n793), .Z(n794) );
  NOR2_X1 U890 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U891 ( .A(KEYINPUT36), .B(n796), .ZN(n871) );
  XNOR2_X1 U892 ( .A(G2067), .B(KEYINPUT37), .ZN(n826) );
  NOR2_X1 U893 ( .A1(n871), .A2(n826), .ZN(n970) );
  NAND2_X1 U894 ( .A1(n829), .A2(n970), .ZN(n824) );
  AND2_X1 U895 ( .A1(n797), .A2(n824), .ZN(n798) );
  NAND2_X1 U896 ( .A1(n799), .A2(n798), .ZN(n815) );
  INV_X1 U897 ( .A(n824), .ZN(n813) );
  NOR2_X1 U898 ( .A1(G2090), .A2(G303), .ZN(n800) );
  NAND2_X1 U899 ( .A1(G8), .A2(n800), .ZN(n805) );
  NOR2_X1 U900 ( .A1(G1981), .A2(G305), .ZN(n801) );
  XOR2_X1 U901 ( .A(n801), .B(KEYINPUT24), .Z(n802) );
  NOR2_X1 U902 ( .A1(n808), .A2(n802), .ZN(n803) );
  XNOR2_X1 U903 ( .A(n803), .B(KEYINPUT94), .ZN(n809) );
  INV_X1 U904 ( .A(n809), .ZN(n804) );
  AND2_X1 U905 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U906 ( .A1(n807), .A2(n806), .ZN(n811) );
  OR2_X1 U907 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U908 ( .A1(n519), .A2(n520), .ZN(n812) );
  OR2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U910 ( .A(n816), .B(KEYINPUT102), .ZN(n831) );
  NOR2_X1 U911 ( .A1(G1996), .A2(n856), .ZN(n961) );
  INV_X1 U912 ( .A(n817), .ZN(n821) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n818) );
  NOR2_X1 U914 ( .A1(G1991), .A2(n875), .ZN(n953) );
  NOR2_X1 U915 ( .A1(n818), .A2(n953), .ZN(n819) );
  XOR2_X1 U916 ( .A(KEYINPUT103), .B(n819), .Z(n820) );
  NOR2_X1 U917 ( .A1(n821), .A2(n820), .ZN(n822) );
  NOR2_X1 U918 ( .A1(n961), .A2(n822), .ZN(n823) );
  XNOR2_X1 U919 ( .A(n823), .B(KEYINPUT39), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n871), .A2(n826), .ZN(n967) );
  NAND2_X1 U922 ( .A1(n827), .A2(n967), .ZN(n828) );
  NAND2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n831), .A2(n830), .ZN(n833) );
  XNOR2_X1 U925 ( .A(KEYINPUT40), .B(KEYINPUT104), .ZN(n832) );
  XNOR2_X1 U926 ( .A(n833), .B(n832), .ZN(G329) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U929 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U931 ( .A1(n837), .A2(n836), .ZN(G188) );
  INV_X1 U933 ( .A(G120), .ZN(G236) );
  INV_X1 U934 ( .A(G108), .ZN(G238) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  NOR2_X1 U937 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  NAND2_X1 U939 ( .A1(n865), .A2(G112), .ZN(n840) );
  XNOR2_X1 U940 ( .A(n840), .B(KEYINPUT114), .ZN(n842) );
  NAND2_X1 U941 ( .A1(G100), .A2(n861), .ZN(n841) );
  NAND2_X1 U942 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n843), .B(KEYINPUT115), .ZN(n845) );
  NAND2_X1 U944 ( .A1(G136), .A2(n564), .ZN(n844) );
  NAND2_X1 U945 ( .A1(n845), .A2(n844), .ZN(n848) );
  NAND2_X1 U946 ( .A1(n864), .A2(G124), .ZN(n846) );
  XOR2_X1 U947 ( .A(KEYINPUT44), .B(n846), .Z(n847) );
  NOR2_X1 U948 ( .A1(n848), .A2(n847), .ZN(G162) );
  NAND2_X1 U949 ( .A1(G130), .A2(n864), .ZN(n850) );
  NAND2_X1 U950 ( .A1(G118), .A2(n865), .ZN(n849) );
  NAND2_X1 U951 ( .A1(n850), .A2(n849), .ZN(n855) );
  NAND2_X1 U952 ( .A1(G106), .A2(n861), .ZN(n852) );
  NAND2_X1 U953 ( .A1(G142), .A2(n564), .ZN(n851) );
  NAND2_X1 U954 ( .A1(n852), .A2(n851), .ZN(n853) );
  XOR2_X1 U955 ( .A(n853), .B(KEYINPUT45), .Z(n854) );
  NOR2_X1 U956 ( .A1(n855), .A2(n854), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U958 ( .A(n858), .B(KEYINPUT46), .Z(n860) );
  XNOR2_X1 U959 ( .A(KEYINPUT48), .B(KEYINPUT116), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n879) );
  NAND2_X1 U961 ( .A1(G103), .A2(n861), .ZN(n863) );
  NAND2_X1 U962 ( .A1(G139), .A2(n564), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n870) );
  NAND2_X1 U964 ( .A1(G127), .A2(n864), .ZN(n867) );
  NAND2_X1 U965 ( .A1(G115), .A2(n865), .ZN(n866) );
  NAND2_X1 U966 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U967 ( .A(KEYINPUT47), .B(n868), .Z(n869) );
  NOR2_X1 U968 ( .A1(n870), .A2(n869), .ZN(n956) );
  XNOR2_X1 U969 ( .A(n871), .B(n956), .ZN(n873) );
  XNOR2_X1 U970 ( .A(G160), .B(G164), .ZN(n872) );
  XNOR2_X1 U971 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U972 ( .A(n951), .B(n874), .ZN(n877) );
  XNOR2_X1 U973 ( .A(n875), .B(G162), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U975 ( .A(n879), .B(n878), .Z(n880) );
  NOR2_X1 U976 ( .A1(G37), .A2(n880), .ZN(G395) );
  XNOR2_X1 U977 ( .A(G286), .B(n978), .ZN(n882) );
  XNOR2_X1 U978 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U979 ( .A(n883), .B(G171), .ZN(n884) );
  NOR2_X1 U980 ( .A1(G37), .A2(n884), .ZN(G397) );
  XOR2_X1 U981 ( .A(G1966), .B(G1971), .Z(n886) );
  XNOR2_X1 U982 ( .A(G1986), .B(G1976), .ZN(n885) );
  XNOR2_X1 U983 ( .A(n886), .B(n885), .ZN(n898) );
  XOR2_X1 U984 ( .A(G1956), .B(G1961), .Z(n888) );
  XNOR2_X1 U985 ( .A(G1996), .B(G1981), .ZN(n887) );
  XNOR2_X1 U986 ( .A(n888), .B(n887), .ZN(n892) );
  XOR2_X1 U987 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n890) );
  XNOR2_X1 U988 ( .A(G1991), .B(KEYINPUT41), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n896) );
  XOR2_X1 U991 ( .A(KEYINPUT111), .B(G2474), .Z(n894) );
  XNOR2_X1 U992 ( .A(KEYINPUT110), .B(KEYINPUT109), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U995 ( .A(n898), .B(n897), .ZN(G229) );
  XOR2_X1 U996 ( .A(KEYINPUT43), .B(G2678), .Z(n900) );
  XNOR2_X1 U997 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U999 ( .A(KEYINPUT42), .B(G2090), .Z(n902) );
  XNOR2_X1 U1000 ( .A(G2067), .B(G2072), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1002 ( .A(n904), .B(n903), .Z(n906) );
  XNOR2_X1 U1003 ( .A(G2096), .B(G2100), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n908) );
  XOR2_X1 U1005 ( .A(G2078), .B(G2084), .Z(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(G227) );
  XOR2_X1 U1007 ( .A(G2454), .B(G2435), .Z(n910) );
  XNOR2_X1 U1008 ( .A(G2438), .B(G2427), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(n910), .B(n909), .ZN(n917) );
  XOR2_X1 U1010 ( .A(KEYINPUT105), .B(G2446), .Z(n912) );
  XNOR2_X1 U1011 ( .A(G2443), .B(G2430), .ZN(n911) );
  XNOR2_X1 U1012 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1013 ( .A(n913), .B(G2451), .Z(n915) );
  XNOR2_X1 U1014 ( .A(G1341), .B(G1348), .ZN(n914) );
  XNOR2_X1 U1015 ( .A(n915), .B(n914), .ZN(n916) );
  XNOR2_X1 U1016 ( .A(n917), .B(n916), .ZN(n918) );
  NAND2_X1 U1017 ( .A1(n918), .A2(G14), .ZN(n919) );
  XOR2_X1 U1018 ( .A(KEYINPUT106), .B(n919), .Z(G401) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n920) );
  XNOR2_X1 U1020 ( .A(KEYINPUT118), .B(n920), .ZN(n927) );
  NOR2_X1 U1021 ( .A1(G229), .A2(G227), .ZN(n921) );
  XNOR2_X1 U1022 ( .A(n921), .B(KEYINPUT49), .ZN(n925) );
  NOR2_X1 U1023 ( .A1(n922), .A2(G401), .ZN(n923) );
  XNOR2_X1 U1024 ( .A(KEYINPUT117), .B(n923), .ZN(n924) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(G225) );
  INV_X1 U1027 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1028 ( .A(G29), .B(KEYINPUT122), .Z(n948) );
  XNOR2_X1 U1029 ( .A(G27), .B(n928), .ZN(n938) );
  XOR2_X1 U1030 ( .A(G1991), .B(G25), .Z(n929) );
  NAND2_X1 U1031 ( .A1(G28), .A2(n929), .ZN(n930) );
  XNOR2_X1 U1032 ( .A(n930), .B(KEYINPUT121), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(G2067), .B(G26), .ZN(n932) );
  XNOR2_X1 U1034 ( .A(G2072), .B(G33), .ZN(n931) );
  NOR2_X1 U1035 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1036 ( .A1(n934), .A2(n933), .ZN(n936) );
  XNOR2_X1 U1037 ( .A(G32), .B(G1996), .ZN(n935) );
  NOR2_X1 U1038 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1040 ( .A(n939), .B(KEYINPUT53), .ZN(n942) );
  XOR2_X1 U1041 ( .A(G2084), .B(G34), .Z(n940) );
  XNOR2_X1 U1042 ( .A(KEYINPUT54), .B(n940), .ZN(n941) );
  NAND2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(KEYINPUT120), .B(G2090), .ZN(n943) );
  XNOR2_X1 U1045 ( .A(G35), .B(n943), .ZN(n944) );
  NOR2_X1 U1046 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1047 ( .A(n946), .B(KEYINPUT55), .ZN(n947) );
  NAND2_X1 U1048 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1049 ( .A1(G11), .A2(n949), .ZN(n977) );
  INV_X1 U1050 ( .A(G29), .ZN(n975) );
  XNOR2_X1 U1051 ( .A(KEYINPUT119), .B(KEYINPUT52), .ZN(n972) );
  XOR2_X1 U1052 ( .A(G2084), .B(G160), .Z(n950) );
  NOR2_X1 U1053 ( .A1(n951), .A2(n950), .ZN(n955) );
  NOR2_X1 U1054 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1055 ( .A1(n955), .A2(n954), .ZN(n966) );
  XOR2_X1 U1056 ( .A(G2072), .B(n956), .Z(n958) );
  XOR2_X1 U1057 ( .A(G164), .B(G2078), .Z(n957) );
  NOR2_X1 U1058 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1059 ( .A(KEYINPUT50), .B(n959), .ZN(n964) );
  XOR2_X1 U1060 ( .A(G2090), .B(G162), .Z(n960) );
  NOR2_X1 U1061 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1062 ( .A(KEYINPUT51), .B(n962), .Z(n963) );
  NAND2_X1 U1063 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1064 ( .A1(n966), .A2(n965), .ZN(n968) );
  NAND2_X1 U1065 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1067 ( .A(n972), .B(n971), .ZN(n973) );
  NOR2_X1 U1068 ( .A1(n973), .A2(KEYINPUT55), .ZN(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n1004) );
  XNOR2_X1 U1071 ( .A(KEYINPUT56), .B(G16), .ZN(n1002) );
  XOR2_X1 U1072 ( .A(G171), .B(G1961), .Z(n980) );
  XNOR2_X1 U1073 ( .A(n978), .B(G1348), .ZN(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n987) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n984) );
  AND2_X1 U1076 ( .A1(G303), .A2(G1971), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1078 ( .A(KEYINPUT123), .B(n985), .Z(n986) );
  NAND2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n992) );
  XOR2_X1 U1080 ( .A(G1966), .B(G168), .Z(n988) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1082 ( .A(n990), .B(KEYINPUT57), .ZN(n991) );
  NOR2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n1000) );
  XOR2_X1 U1084 ( .A(n993), .B(G1341), .Z(n996) );
  XNOR2_X1 U1085 ( .A(n994), .B(G1956), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1032) );
  XNOR2_X1 U1091 ( .A(G1986), .B(G24), .ZN(n1009) );
  XNOR2_X1 U1092 ( .A(G1976), .B(G23), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(G1971), .B(G22), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(KEYINPUT127), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(KEYINPUT58), .B(n1010), .ZN(n1026) );
  XOR2_X1 U1098 ( .A(G1981), .B(G6), .Z(n1013) );
  XNOR2_X1 U1099 ( .A(n1011), .B(G19), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XNOR2_X1 U1101 ( .A(G20), .B(G1956), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(KEYINPUT124), .B(n1016), .ZN(n1020) );
  XOR2_X1 U1104 ( .A(KEYINPUT125), .B(G4), .Z(n1018) );
  XNOR2_X1 U1105 ( .A(G1348), .B(KEYINPUT59), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(n1018), .B(n1017), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(n1021), .B(KEYINPUT60), .ZN(n1024) );
  XNOR2_X1 U1109 ( .A(KEYINPUT126), .B(G1966), .ZN(n1022) );
  XNOR2_X1 U1110 ( .A(G21), .B(n1022), .ZN(n1023) );
  NOR2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1028) );
  XNOR2_X1 U1113 ( .A(G5), .B(G1961), .ZN(n1027) );
  NOR2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1115 ( .A(KEYINPUT61), .B(n1029), .Z(n1030) );
  NOR2_X1 U1116 ( .A1(G16), .A2(n1030), .ZN(n1031) );
  NOR2_X1 U1117 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1118 ( .A(n1033), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

