//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n553, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n598, new_n601, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1177;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n461));
  INV_X1    g036(.A(G137), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g043(.A(new_n463), .B(KEYINPUT66), .C1(new_n465), .C2(new_n464), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n461), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n473), .ZN(new_n475));
  AOI211_X1 g050(.A(KEYINPUT67), .B(new_n475), .C1(new_n468), .C2(new_n469), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  AOI22_X1  g052(.A1(new_n477), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n478));
  INV_X1    g053(.A(G2105), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR3_X1   g055(.A1(new_n474), .A2(new_n476), .A3(new_n480), .ZN(G160));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n482));
  OR2_X1    g057(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n477), .A2(new_n482), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(new_n479), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n479), .A3(new_n484), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  OR2_X1    g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G112), .C2(new_n479), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n487), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n464), .B2(new_n465), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n477), .A2(new_n499), .A3(new_n496), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(G126), .B1(new_n464), .B2(new_n465), .ZN(new_n502));
  NAND2_X1  g077(.A1(G114), .A2(G2104), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G2105), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n472), .A2(G102), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n501), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  NAND2_X1  g083(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n512));
  NAND4_X1  g087(.A1(KEYINPUT70), .A2(KEYINPUT71), .A3(KEYINPUT5), .A4(G543), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT69), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n516), .B2(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(KEYINPUT69), .A3(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(KEYINPUT6), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n514), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n520), .A2(G543), .A3(new_n521), .ZN(new_n524));
  INV_X1    g099(.A(G50), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n522), .A2(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n516), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n526), .A2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  INV_X1    g105(.A(new_n522), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G89), .ZN(new_n532));
  INV_X1    g107(.A(new_n524), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G51), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n532), .A2(new_n534), .A3(new_n536), .A4(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n522), .A2(new_n540), .B1(new_n524), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n516), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(G171));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n522), .A2(new_n546), .B1(new_n524), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n516), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n553), .A2(new_n556), .ZN(G188));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n520), .A2(G53), .A3(G543), .A4(new_n521), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n560));
  OAI211_X1 g135(.A(KEYINPUT72), .B(new_n558), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT72), .B1(new_n559), .B2(new_n560), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT9), .B1(new_n559), .B2(KEYINPUT72), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n561), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT74), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n514), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n568), .A2(new_n516), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(G91), .B2(new_n531), .ZN(new_n570));
  OAI211_X1 g145(.A(new_n562), .B(KEYINPUT9), .C1(KEYINPUT72), .C2(new_n559), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n571), .A2(KEYINPUT74), .A3(new_n561), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n567), .A2(new_n570), .A3(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  NAND4_X1  g149(.A1(new_n514), .A2(new_n520), .A3(G87), .A4(new_n521), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n520), .A2(G49), .A3(G543), .A4(new_n521), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G288));
  NAND4_X1  g153(.A1(new_n514), .A2(new_n520), .A3(G86), .A4(new_n521), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n520), .A2(G48), .A3(G543), .A4(new_n521), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n514), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n516), .ZN(G305));
  AOI22_X1  g157(.A1(new_n531), .A2(G85), .B1(new_n533), .B2(G47), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n516), .B2(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n531), .A2(G92), .ZN(new_n587));
  XOR2_X1   g162(.A(new_n587), .B(KEYINPUT10), .Z(new_n588));
  XNOR2_X1  g163(.A(KEYINPUT75), .B(G66), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n514), .A2(new_n589), .B1(G79), .B2(G543), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT76), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(G54), .B2(new_n533), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n586), .B1(new_n594), .B2(G868), .ZN(G284));
  OAI21_X1  g170(.A(new_n586), .B1(new_n594), .B2(G868), .ZN(G321));
  NAND2_X1  g171(.A1(G286), .A2(G868), .ZN(new_n597));
  INV_X1    g172(.A(G299), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(G868), .ZN(G297));
  OAI21_X1  g174(.A(new_n597), .B1(new_n598), .B2(G868), .ZN(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n594), .B1(new_n601), .B2(G860), .ZN(G148));
  NAND2_X1  g177(.A1(new_n594), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G868), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g181(.A1(new_n486), .A2(G123), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n489), .A2(G135), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n479), .A2(G111), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(KEYINPUT79), .ZN(new_n610));
  OAI21_X1  g185(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n609), .A2(KEYINPUT79), .B1(new_n611), .B2(KEYINPUT80), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(KEYINPUT80), .B2(new_n611), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n607), .B(new_n608), .C1(new_n610), .C2(new_n613), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT81), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2096), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n477), .A2(new_n472), .ZN(new_n617));
  XOR2_X1   g192(.A(KEYINPUT77), .B(KEYINPUT12), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  AND2_X1   g195(.A1(KEYINPUT78), .A2(G2100), .ZN(new_n621));
  NOR2_X1   g196(.A1(KEYINPUT78), .A2(G2100), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n616), .B(new_n623), .C1(new_n621), .C2(new_n620), .ZN(G156));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2430), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2435), .ZN(new_n626));
  XOR2_X1   g201(.A(G2427), .B(G2438), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(KEYINPUT14), .ZN(new_n629));
  XOR2_X1   g204(.A(G2443), .B(G2446), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(KEYINPUT82), .B(KEYINPUT16), .Z(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n631), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n635), .B(new_n636), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G14), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(G401));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2067), .B(G2678), .Z(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(new_n644), .A3(KEYINPUT17), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT18), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2072), .B(G2078), .Z(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(new_n643), .B2(KEYINPUT18), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n647), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2096), .B(G2100), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(G227));
  INV_X1    g227(.A(KEYINPUT20), .ZN(new_n653));
  XOR2_X1   g228(.A(G1961), .B(G1966), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT83), .ZN(new_n655));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1971), .B(G1976), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n653), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n655), .A2(new_n656), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n662), .A2(new_n659), .A3(new_n657), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n657), .A2(new_n653), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n664), .A2(new_n661), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n660), .B(new_n663), .C1(new_n665), .C2(new_n659), .ZN(new_n666));
  XOR2_X1   g241(.A(G1991), .B(G1996), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G229));
  NAND2_X1  g247(.A1(new_n486), .A2(G129), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT93), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n472), .A2(G105), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT94), .ZN(new_n676));
  NAND3_X1  g251(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT26), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n489), .B2(G141), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n674), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  MUX2_X1   g255(.A(G32), .B(new_n680), .S(G29), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT95), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT27), .B(G1996), .Z(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n684), .ZN(new_n686));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  AND2_X1   g262(.A1(KEYINPUT30), .A2(G28), .ZN(new_n688));
  NOR2_X1   g263(.A1(KEYINPUT30), .A2(G28), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(new_n614), .B2(new_n687), .ZN(new_n691));
  INV_X1    g266(.A(G2072), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n687), .A2(G33), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n472), .A2(G103), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT25), .Z(new_n695));
  AOI22_X1  g270(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n696));
  INV_X1    g271(.A(G139), .ZN(new_n697));
  OAI221_X1 g272(.A(new_n695), .B1(new_n479), .B2(new_n696), .C1(new_n488), .C2(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n693), .B1(new_n698), .B2(G29), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n691), .B1(new_n692), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(G171), .A2(G16), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G5), .B2(G16), .ZN(new_n702));
  INV_X1    g277(.A(G1961), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n700), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NOR3_X1   g281(.A1(new_n685), .A2(new_n686), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n687), .A2(G26), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n486), .A2(G128), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n489), .A2(G140), .ZN(new_n711));
  NOR2_X1   g286(.A1(G104), .A2(G2105), .ZN(new_n712));
  OAI21_X1  g287(.A(G2104), .B1(new_n479), .B2(G116), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n710), .B(new_n711), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  AND3_X1   g289(.A1(new_n714), .A2(KEYINPUT91), .A3(G29), .ZN(new_n715));
  AOI21_X1  g290(.A(KEYINPUT91), .B1(new_n714), .B2(G29), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n709), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G2067), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT31), .B(G11), .ZN(new_n720));
  AND2_X1   g295(.A1(KEYINPUT24), .A2(G34), .ZN(new_n721));
  NOR2_X1   g296(.A1(KEYINPUT24), .A2(G34), .ZN(new_n722));
  NOR3_X1   g297(.A1(new_n721), .A2(new_n722), .A3(G29), .ZN(new_n723));
  INV_X1    g298(.A(G160), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(G29), .ZN(new_n725));
  INV_X1    g300(.A(G2084), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G16), .ZN(new_n728));
  NOR2_X1   g303(.A1(G168), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n728), .B2(G21), .ZN(new_n730));
  INV_X1    g305(.A(G1966), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n727), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT86), .B(G16), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G19), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n551), .B2(new_n734), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(G1341), .Z(new_n737));
  NOR2_X1   g312(.A1(G27), .A2(G29), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G164), .B2(G29), .ZN(new_n739));
  INV_X1    g314(.A(G2078), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n737), .B(new_n741), .C1(new_n692), .C2(new_n699), .ZN(new_n742));
  AOI211_X1 g317(.A(new_n732), .B(new_n742), .C1(new_n731), .C2(new_n730), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n707), .A2(new_n719), .A3(new_n720), .A4(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n734), .A2(KEYINPUT23), .A3(G20), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT23), .ZN(new_n746));
  INV_X1    g321(.A(G20), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n746), .B1(new_n733), .B2(new_n747), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n745), .B(new_n748), .C1(new_n598), .C2(new_n728), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G1956), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n687), .A2(G35), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G162), .B2(new_n687), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT29), .B(G2090), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n728), .A2(G4), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n594), .B2(new_n728), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT90), .B(G1348), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NOR4_X1   g333(.A1(new_n744), .A2(new_n750), .A3(new_n754), .A4(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n725), .A2(new_n726), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT92), .ZN(new_n761));
  MUX2_X1   g336(.A(G24), .B(G290), .S(new_n733), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1986), .ZN(new_n763));
  NAND2_X1  g338(.A1(G166), .A2(new_n733), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G22), .B2(new_n733), .ZN(new_n765));
  INV_X1    g340(.A(G1971), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT32), .B(G1981), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT88), .ZN(new_n769));
  MUX2_X1   g344(.A(G6), .B(G305), .S(G16), .Z(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n767), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n769), .B2(new_n771), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n765), .A2(new_n766), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n728), .A2(G23), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT89), .ZN(new_n776));
  NAND2_X1  g351(.A1(G288), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n575), .A2(new_n576), .A3(new_n577), .A4(KEYINPUT89), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n775), .B1(new_n779), .B2(new_n728), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT33), .B(G1976), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n773), .A2(new_n774), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT87), .B(KEYINPUT34), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n763), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n486), .A2(G119), .ZN(new_n787));
  NOR2_X1   g362(.A1(G95), .A2(G2105), .ZN(new_n788));
  OAI21_X1  g363(.A(G2104), .B1(new_n479), .B2(G107), .ZN(new_n789));
  AND3_X1   g364(.A1(new_n489), .A2(KEYINPUT84), .A3(G131), .ZN(new_n790));
  AOI21_X1  g365(.A(KEYINPUT84), .B1(new_n489), .B2(G131), .ZN(new_n791));
  OAI221_X1 g366(.A(new_n787), .B1(new_n788), .B2(new_n789), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  MUX2_X1   g367(.A(G25), .B(new_n792), .S(G29), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT85), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT35), .B(G1991), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n786), .B(new_n796), .C1(new_n785), .C2(new_n784), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT36), .ZN(new_n798));
  AND3_X1   g373(.A1(new_n759), .A2(new_n761), .A3(new_n798), .ZN(G311));
  NAND3_X1  g374(.A1(new_n759), .A2(new_n761), .A3(new_n798), .ZN(G150));
  AND2_X1   g375(.A1(new_n514), .A2(G67), .ZN(new_n801));
  AND2_X1   g376(.A1(G80), .A2(G543), .ZN(new_n802));
  OAI21_X1  g377(.A(G651), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(G93), .ZN(new_n804));
  INV_X1    g379(.A(G55), .ZN(new_n805));
  OAI22_X1  g380(.A1(new_n522), .A2(new_n804), .B1(new_n524), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n806), .A2(KEYINPUT96), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(KEYINPUT96), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n803), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(G860), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT37), .Z(new_n811));
  NAND2_X1  g386(.A1(new_n594), .A2(G559), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT38), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n809), .A2(new_n551), .ZN(new_n814));
  OAI221_X1 g389(.A(new_n803), .B1(new_n550), .B2(new_n548), .C1(new_n807), .C2(new_n808), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT39), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n813), .B(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n811), .B1(new_n818), .B2(G860), .ZN(G145));
  XNOR2_X1  g394(.A(new_n680), .B(G164), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n698), .A2(KEYINPUT99), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n714), .B(new_n821), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(G142), .ZN(new_n824));
  NOR2_X1   g399(.A1(G106), .A2(G2105), .ZN(new_n825));
  OAI21_X1  g400(.A(G2104), .B1(new_n479), .B2(G118), .ZN(new_n826));
  OAI22_X1  g401(.A1(new_n488), .A2(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(G130), .B2(new_n486), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n619), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n792), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT100), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n823), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n830), .A2(new_n831), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n823), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n724), .B(new_n614), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n493), .B(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n837), .B(new_n839), .Z(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n836), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(G37), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n833), .A2(new_n835), .A3(new_n840), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g421(.A(G868), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT106), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n779), .B(KEYINPUT104), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G290), .ZN(new_n850));
  XOR2_X1   g425(.A(G303), .B(G305), .Z(new_n851));
  INV_X1    g426(.A(KEYINPUT105), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT42), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n851), .A2(new_n852), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n850), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n855), .B1(new_n854), .B2(new_n857), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n848), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n603), .B(new_n816), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n598), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(G299), .A2(KEYINPUT101), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(new_n593), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n598), .A2(new_n594), .A3(new_n863), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n862), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT102), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(new_n868), .B2(KEYINPUT41), .ZN(new_n871));
  XNOR2_X1  g446(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT41), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n866), .A2(KEYINPUT102), .A3(new_n874), .A4(new_n867), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n871), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n869), .B1(new_n876), .B2(new_n862), .ZN(new_n877));
  INV_X1    g452(.A(new_n860), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(KEYINPUT106), .A3(new_n858), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n861), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n877), .A2(new_n861), .A3(new_n879), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n847), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n809), .A2(G868), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n883), .A2(KEYINPUT107), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT107), .ZN(new_n887));
  INV_X1    g462(.A(new_n882), .ZN(new_n888));
  OAI21_X1  g463(.A(G868), .B1(new_n888), .B2(new_n880), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n887), .B1(new_n889), .B2(new_n884), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n886), .A2(new_n890), .ZN(G295));
  NOR2_X1   g466(.A1(new_n883), .A2(new_n885), .ZN(G331));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n893));
  XNOR2_X1  g468(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n854), .A2(new_n857), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n816), .A2(G171), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n814), .A2(new_n815), .A3(G301), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(G286), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n897), .A2(G168), .A3(new_n898), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n876), .A2(new_n902), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n902), .A2(new_n868), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n896), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n902), .A2(new_n868), .ZN(new_n906));
  INV_X1    g481(.A(new_n896), .ZN(new_n907));
  AOI211_X1 g482(.A(new_n906), .B(new_n907), .C1(new_n876), .C2(new_n902), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n895), .B1(new_n909), .B2(new_n843), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n903), .A2(new_n896), .A3(new_n904), .ZN(new_n911));
  INV_X1    g486(.A(new_n872), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n902), .B1(new_n868), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT41), .B1(new_n866), .B2(new_n867), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n904), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n907), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n911), .A2(new_n843), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n917), .A2(new_n894), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n893), .B1(new_n910), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n893), .B1(new_n917), .B2(KEYINPUT43), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n921));
  INV_X1    g496(.A(new_n905), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n922), .A2(new_n843), .A3(new_n895), .A4(new_n911), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n921), .B1(new_n920), .B2(new_n923), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n919), .B1(new_n924), .B2(new_n925), .ZN(G397));
  INV_X1    g501(.A(G1384), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n507), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT45), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n469), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT66), .B1(new_n477), .B2(new_n463), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n473), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT67), .ZN(new_n934));
  INV_X1    g509(.A(new_n480), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n470), .A2(new_n461), .A3(new_n473), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n934), .A2(G40), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n930), .A2(new_n937), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n680), .A2(G1996), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n714), .B(new_n718), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n680), .A2(G1996), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n792), .B(new_n795), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n938), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AND2_X1   g519(.A1(G290), .A2(G1986), .ZN(new_n945));
  NOR2_X1   g520(.A1(G290), .A2(G1986), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n938), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT110), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n928), .A2(new_n951), .A3(KEYINPUT50), .ZN(new_n952));
  INV_X1    g527(.A(new_n506), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n953), .B1(new_n504), .B2(G2105), .ZN(new_n954));
  AOI21_X1  g529(.A(G1384), .B1(new_n954), .B2(new_n501), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT50), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT111), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n952), .A2(new_n957), .ZN(new_n958));
  AOI211_X1 g533(.A(KEYINPUT50), .B(G1384), .C1(new_n954), .C2(new_n501), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n937), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n958), .A2(new_n960), .A3(new_n726), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n955), .A2(KEYINPUT45), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT115), .ZN(new_n964));
  NAND4_X1  g539(.A1(G160), .A2(new_n930), .A3(new_n964), .A4(G40), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n955), .A2(KEYINPUT45), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT115), .B1(new_n937), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n963), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n961), .B1(new_n968), .B2(G1966), .ZN(new_n969));
  XOR2_X1   g544(.A(KEYINPUT113), .B(G8), .Z(new_n970));
  AND3_X1   g545(.A1(new_n969), .A2(G168), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT55), .ZN(new_n975));
  INV_X1    g550(.A(G8), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n975), .B1(G166), .B2(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(G303), .A2(KEYINPUT112), .A3(KEYINPUT55), .A4(G8), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n974), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND4_X1  g554(.A1(G160), .A2(new_n930), .A3(G40), .A4(new_n962), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n956), .B1(new_n507), .B2(new_n927), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n937), .A2(new_n981), .A3(new_n959), .ZN(new_n982));
  INV_X1    g557(.A(G2090), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n766), .A2(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n970), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n979), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n970), .B1(new_n937), .B2(new_n928), .ZN(new_n987));
  INV_X1    g562(.A(G1976), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n777), .B2(new_n778), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT52), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n581), .A2(new_n516), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n579), .A2(new_n580), .ZN(new_n992));
  INV_X1    g567(.A(G1981), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(G305), .A2(G1981), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT49), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n474), .A2(new_n476), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n999), .A2(G40), .A3(new_n935), .A4(new_n955), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n994), .A2(new_n995), .A3(KEYINPUT49), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n998), .A2(new_n1000), .A3(new_n970), .A4(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n989), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT52), .B1(G288), .B2(new_n988), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1000), .A2(new_n1003), .A3(new_n970), .A4(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n990), .A2(new_n1002), .A3(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n974), .A2(new_n977), .A3(new_n978), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n980), .A2(new_n766), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n958), .A2(new_n960), .A3(new_n983), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n976), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1006), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n971), .A2(KEYINPUT116), .A3(new_n986), .A4(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(G8), .A3(new_n1007), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n990), .A2(new_n1002), .A3(new_n1005), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n986), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n969), .A2(G168), .A3(new_n970), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1013), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT63), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1012), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n1010), .A2(new_n1007), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n971), .A2(KEYINPUT63), .A3(new_n1011), .A4(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1016), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1002), .A2(new_n988), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1026), .A2(G288), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n994), .B(KEYINPUT114), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n987), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1024), .A2(new_n1025), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n958), .A2(new_n960), .ZN(new_n1032));
  INV_X1    g607(.A(G1348), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1000), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n718), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT60), .ZN(new_n1038));
  OAI211_X1 g613(.A(KEYINPUT120), .B(new_n593), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1032), .A2(new_n1033), .B1(new_n1035), .B2(new_n718), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n593), .A2(KEYINPUT120), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n593), .A2(KEYINPUT120), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1041), .A2(new_n1042), .A3(KEYINPUT60), .A4(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1039), .A2(new_n1040), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT121), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1039), .A2(KEYINPUT121), .A3(new_n1040), .A4(new_n1044), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  XOR2_X1   g624(.A(KEYINPUT58), .B(G1341), .Z(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n937), .B2(new_n928), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1051), .B(KEYINPUT118), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(G1996), .B2(new_n980), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT119), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT59), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1053), .A2(new_n551), .A3(new_n1055), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1054), .A2(KEYINPUT59), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1056), .B(new_n1057), .ZN(new_n1058));
  OR3_X1    g633(.A1(new_n937), .A2(new_n981), .A3(new_n959), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n1060));
  INV_X1    g635(.A(G1956), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT117), .B1(new_n982), .B2(G1956), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n570), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(new_n565), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1067), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n963), .A2(new_n937), .A3(new_n966), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT56), .B(G2072), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1064), .A2(new_n1068), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1068), .B1(new_n1064), .B2(new_n1071), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT61), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1064), .A2(new_n1071), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1068), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT61), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(new_n1079), .A3(new_n1072), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1075), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1049), .A2(new_n1058), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1037), .A2(new_n594), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1073), .B1(new_n1078), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n969), .ZN(new_n1087));
  NAND2_X1  g662(.A1(G286), .A2(new_n970), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n969), .A2(new_n970), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT122), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n1095));
  AOI211_X1 g670(.A(new_n1095), .B(new_n1092), .C1(new_n969), .C2(new_n970), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n969), .A2(G8), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1091), .B1(new_n1098), .B2(new_n1088), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1089), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1069), .A2(new_n740), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT123), .B(G1961), .Z(new_n1104));
  AOI22_X1  g679(.A1(new_n1102), .A2(new_n1103), .B1(new_n1032), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1103), .A2(G2078), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n968), .A2(new_n1106), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1105), .A2(G301), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n999), .A2(KEYINPUT124), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n474), .B2(new_n476), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n930), .A2(G40), .A3(new_n935), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT125), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1114), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT125), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1115), .A2(new_n962), .A3(new_n1119), .A4(new_n1106), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1105), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(G171), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1109), .A2(new_n1122), .A3(KEYINPUT54), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1017), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(G171), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1120), .A2(G301), .A3(new_n1105), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT54), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1101), .A2(new_n1125), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1031), .B1(new_n1086), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT126), .B1(new_n1101), .B2(new_n1132), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n1127), .A2(new_n1017), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1134), .B1(new_n1101), .B2(new_n1132), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT126), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1099), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1136), .B(KEYINPUT62), .C1(new_n1137), .C2(new_n1089), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1133), .A2(new_n1135), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n950), .B1(new_n1131), .B2(new_n1139), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n942), .A2(new_n795), .A3(new_n792), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n714), .A2(G2067), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n938), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n938), .A2(new_n946), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT48), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n944), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n940), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n938), .B1(new_n1147), .B2(new_n680), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n930), .A2(new_n937), .A3(G1996), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n1149), .A2(KEYINPUT46), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(KEYINPUT46), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1148), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT47), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1143), .A2(new_n1146), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT127), .B1(new_n1140), .B2(new_n1154), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1133), .A2(new_n1135), .A3(new_n1138), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1029), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1047), .A2(new_n1048), .B1(new_n1075), .B2(new_n1080), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1084), .B1(new_n1158), .B2(new_n1058), .ZN(new_n1159));
  AOI21_X1  g734(.A(G301), .B1(new_n1120), .B2(new_n1105), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1160), .A2(new_n1108), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1017), .B1(new_n1161), .B2(KEYINPUT54), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1129), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1162), .B(new_n1163), .C1(new_n1137), .C2(new_n1089), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1025), .B(new_n1157), .C1(new_n1159), .C2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n949), .B1(new_n1156), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1154), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1155), .A2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g745(.A1(G229), .A2(new_n459), .ZN(new_n1172));
  OAI21_X1  g746(.A(new_n1172), .B1(new_n910), .B2(new_n918), .ZN(new_n1173));
  NOR2_X1   g747(.A1(G401), .A2(G227), .ZN(new_n1174));
  NAND2_X1  g748(.A1(new_n845), .A2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g749(.A1(new_n1173), .A2(new_n1175), .ZN(G308));
  INV_X1    g750(.A(new_n1175), .ZN(new_n1177));
  OAI211_X1 g751(.A(new_n1177), .B(new_n1172), .C1(new_n910), .C2(new_n918), .ZN(G225));
endmodule


