//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT85), .ZN(new_n203));
  XOR2_X1   g002(.A(G169gat), .B(G197gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n205), .B(new_n206), .Z(new_n207));
  XOR2_X1   g006(.A(new_n207), .B(KEYINPUT12), .Z(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT92), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT89), .ZN(new_n211));
  XNOR2_X1  g010(.A(G15gat), .B(G22gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT16), .ZN(new_n213));
  AOI21_X1  g012(.A(G1gat), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT88), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n214), .B(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT90), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n211), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(G8gat), .B1(new_n217), .B2(new_n211), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n211), .B(G8gat), .C1(new_n217), .C2(new_n218), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G29gat), .ZN(new_n224));
  INV_X1    g023(.A(G36gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT14), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT14), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(G29gat), .B2(G36gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(G29gat), .A2(G36gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G43gat), .B(G50gat), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n232), .A2(KEYINPUT15), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n231), .B1(new_n233), .B2(KEYINPUT87), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT15), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n235), .B1(new_n232), .B2(KEYINPUT86), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(KEYINPUT86), .B2(new_n232), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n233), .A2(KEYINPUT87), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n230), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n210), .B1(new_n223), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n241), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n243), .A2(new_n221), .A3(KEYINPUT92), .A4(new_n222), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n223), .A2(new_n241), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT93), .ZN(new_n247));
  NAND2_X1  g046(.A1(G229gat), .A2(G233gat), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n248), .B(KEYINPUT13), .Z(new_n249));
  NAND3_X1  g048(.A1(new_n246), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n247), .B1(new_n246), .B2(new_n249), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT17), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT91), .B1(new_n241), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT91), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n256), .B(KEYINPUT17), .C1(new_n238), .C2(new_n240), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n223), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n241), .A2(new_n254), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n261), .A2(new_n248), .A3(new_n245), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT18), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n261), .A2(KEYINPUT18), .A3(new_n248), .A4(new_n245), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n209), .B1(new_n253), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n246), .A2(new_n249), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT93), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n250), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n270), .A2(new_n208), .A3(new_n264), .A4(new_n265), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G22gat), .B(G50gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G228gat), .A2(G233gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT3), .ZN(new_n277));
  XNOR2_X1  g076(.A(G197gat), .B(G204gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT22), .ZN(new_n279));
  INV_X1    g078(.A(G211gat), .ZN(new_n280));
  INV_X1    g079(.A(G218gat), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G211gat), .B(G218gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n278), .A3(new_n282), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n286), .A2(KEYINPUT80), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT29), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n289), .B1(new_n286), .B2(KEYINPUT80), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n277), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n292));
  NAND2_X1  g091(.A1(G141gat), .A2(G148gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(G141gat), .A2(G148gat), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n292), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G141gat), .ZN(new_n297));
  INV_X1    g096(.A(G148gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n299), .A2(KEYINPUT75), .A3(new_n293), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT2), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n296), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(G155gat), .B(G162gat), .Z(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G155gat), .ZN(new_n305));
  INV_X1    g104(.A(G162gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n301), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(new_n305), .B2(new_n306), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n294), .A2(new_n295), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n276), .B1(new_n291), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n286), .A2(new_n287), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n313), .B(new_n314), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n302), .A2(new_n303), .B1(new_n309), .B2(new_n308), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT29), .B1(new_n316), .B2(new_n277), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n312), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT29), .B1(new_n286), .B2(new_n287), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n311), .B1(new_n319), .B2(KEYINPUT3), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(new_n315), .B2(new_n317), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n276), .ZN(new_n322));
  XNOR2_X1  g121(.A(G78gat), .B(G106gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(KEYINPUT31), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n318), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n325), .B1(new_n318), .B2(new_n322), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n274), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n318), .A2(new_n322), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n324), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(new_n273), .A3(new_n326), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G127gat), .B(G134gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT69), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G127gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n337), .A2(G134gat), .ZN(new_n338));
  INV_X1    g137(.A(G134gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n339), .A2(G127gat), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT69), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G113gat), .ZN(new_n342));
  INV_X1    g141(.A(G120gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G113gat), .A2(G120gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n336), .B(new_n341), .C1(KEYINPUT1), .C2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT70), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n334), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT70), .B1(new_n338), .B2(new_n340), .ZN(new_n350));
  INV_X1    g149(.A(new_n346), .ZN(new_n351));
  XOR2_X1   g150(.A(KEYINPUT71), .B(KEYINPUT1), .Z(new_n352));
  NAND4_X1  g151(.A1(new_n349), .A2(new_n350), .A3(new_n351), .A4(new_n352), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n347), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G183gat), .A2(G190gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  AND2_X1   g155(.A1(G169gat), .A2(G176gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT26), .ZN(new_n358));
  NOR2_X1   g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n359), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT26), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n356), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT28), .ZN(new_n365));
  INV_X1    g164(.A(G183gat), .ZN(new_n366));
  AOI21_X1  g165(.A(G190gat), .B1(new_n366), .B2(KEYINPUT27), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT27), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT66), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT66), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT27), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n366), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n367), .B1(new_n372), .B2(KEYINPUT67), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT67), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n374), .A2(new_n375), .A3(new_n366), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n365), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n368), .A2(G183gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n367), .A2(KEYINPUT28), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT68), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n367), .A2(KEYINPUT68), .A3(KEYINPUT28), .A4(new_n378), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n364), .B1(new_n377), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT25), .ZN(new_n385));
  OAI211_X1 g184(.A(KEYINPUT64), .B(KEYINPUT24), .C1(G183gat), .C2(G190gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n385), .B1(new_n386), .B2(new_n356), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT64), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT24), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n355), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n387), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT23), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n357), .B1(new_n361), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n359), .A2(KEYINPUT23), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(G190gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n366), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n389), .A2(KEYINPUT65), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n399), .A3(new_n355), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n356), .A2(KEYINPUT65), .A3(new_n389), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n393), .A2(new_n394), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT25), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n396), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n354), .B1(new_n384), .B2(new_n404), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n391), .A2(new_n395), .B1(new_n402), .B2(KEYINPUT25), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n347), .A2(new_n353), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n381), .A2(new_n382), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n372), .A2(KEYINPUT67), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n375), .B1(new_n374), .B2(new_n366), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n410), .A3(new_n367), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n408), .B1(new_n411), .B2(new_n365), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n406), .B(new_n407), .C1(new_n412), .C2(new_n364), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n405), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(G227gat), .ZN(new_n415));
  INV_X1    g214(.A(G233gat), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT34), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n414), .A2(KEYINPUT34), .A3(new_n418), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n405), .A2(new_n417), .A3(new_n413), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT32), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT33), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G15gat), .B(G43gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(G71gat), .B(G99gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n429), .B(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n426), .B1(new_n432), .B2(KEYINPUT33), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n425), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n424), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n333), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT72), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n433), .A2(new_n439), .A3(new_n435), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n425), .A2(new_n434), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n431), .B1(new_n425), .B2(new_n427), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT72), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT73), .B1(new_n444), .B2(new_n424), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT73), .ZN(new_n446));
  AOI211_X1 g245(.A(new_n446), .B(new_n423), .C1(new_n440), .C2(new_n443), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n438), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT4), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n354), .A2(new_n449), .A3(new_n316), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT4), .B1(new_n311), .B2(new_n407), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(G225gat), .A2(G233gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n311), .A2(KEYINPUT3), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n316), .A2(new_n277), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(new_n407), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n452), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(KEYINPUT76), .B(KEYINPUT5), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n460));
  XNOR2_X1  g259(.A(G1gat), .B(G29gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G57gat), .B(G85gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n462), .B(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n311), .B(new_n407), .ZN(new_n465));
  INV_X1    g264(.A(new_n453), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n458), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n452), .A2(new_n453), .A3(new_n456), .A4(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n459), .A2(new_n464), .A3(new_n467), .A4(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(KEYINPUT78), .B(KEYINPUT6), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n469), .A2(new_n467), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n464), .B1(new_n473), .B2(new_n459), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT79), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n464), .ZN(new_n476));
  INV_X1    g275(.A(new_n459), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n469), .A2(new_n467), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT79), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n479), .A2(new_n480), .A3(new_n470), .A4(new_n471), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n470), .A2(new_n471), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n475), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n315), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n406), .B1(new_n412), .B2(new_n364), .ZN(new_n485));
  INV_X1    g284(.A(G226gat), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n486), .A2(new_n416), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n487), .B1(new_n485), .B2(new_n289), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n484), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n384), .A2(new_n404), .ZN(new_n492));
  OAI22_X1  g291(.A1(new_n492), .A2(KEYINPUT29), .B1(new_n486), .B2(new_n416), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n493), .A2(new_n315), .A3(new_n488), .ZN(new_n494));
  XNOR2_X1  g293(.A(G8gat), .B(G36gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(G64gat), .ZN(new_n496));
  INV_X1    g295(.A(G92gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n491), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT30), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n498), .B1(new_n491), .B2(new_n494), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n491), .A2(new_n494), .A3(KEYINPUT30), .A4(new_n498), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n501), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n483), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT35), .B1(new_n448), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT83), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT83), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n509), .B(KEYINPUT35), .C1(new_n448), .C2(new_n506), .ZN(new_n510));
  INV_X1    g309(.A(new_n437), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n424), .A2(new_n436), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n513), .A2(KEYINPUT35), .A3(new_n333), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n502), .B1(new_n500), .B2(new_n499), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n515), .A2(KEYINPUT81), .A3(new_n504), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT81), .B1(new_n515), .B2(new_n504), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n482), .B1(new_n474), .B2(new_n472), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n514), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n508), .A2(new_n510), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n499), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n494), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n315), .B1(new_n493), .B2(new_n488), .ZN(new_n525));
  OR3_X1    g324(.A1(new_n524), .A2(KEYINPUT37), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n498), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT37), .B1(new_n524), .B2(new_n525), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT38), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT38), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n526), .A2(new_n531), .A3(new_n527), .A4(new_n528), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n523), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n333), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT40), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n452), .A2(new_n456), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(new_n466), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n476), .B1(new_n537), .B2(KEYINPUT39), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT39), .B1(new_n465), .B2(new_n466), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n539), .B1(new_n466), .B2(new_n536), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n535), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT82), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  OR3_X1    g342(.A1(new_n538), .A2(new_n540), .A3(new_n535), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n543), .A2(new_n470), .A3(new_n544), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n533), .B(new_n534), .C1(new_n518), .C2(new_n545), .ZN(new_n546));
  OAI211_X1 g345(.A(KEYINPUT36), .B(new_n511), .C1(new_n445), .C2(new_n447), .ZN(new_n547));
  INV_X1    g346(.A(new_n513), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n547), .B1(KEYINPUT36), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n506), .A2(new_n333), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n546), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n272), .B1(new_n521), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT95), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT97), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n553), .B(KEYINPUT95), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT97), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G71gat), .B(G78gat), .ZN(new_n560));
  INV_X1    g359(.A(G64gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n561), .A2(G57gat), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT96), .ZN(new_n563));
  INV_X1    g362(.A(G57gat), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n564), .A2(G64gat), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n562), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(new_n563), .B2(new_n565), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n556), .A2(new_n559), .A3(new_n560), .A4(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n557), .B1(new_n565), .B2(new_n562), .ZN(new_n569));
  NOR3_X1   g368(.A1(KEYINPUT94), .A2(G71gat), .A3(G78gat), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT94), .B1(G71gat), .B2(G78gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  AOI211_X1 g371(.A(new_n570), .B(new_n572), .C1(G71gat), .C2(G78gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n575), .A2(KEYINPUT98), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(KEYINPUT98), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT99), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n575), .A2(KEYINPUT98), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n575), .A2(KEYINPUT98), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT99), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(KEYINPUT21), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n583), .A2(new_n366), .A3(new_n259), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT21), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n578), .B1(new_n576), .B2(new_n577), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n580), .A2(KEYINPUT99), .A3(new_n581), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(G183gat), .B1(new_n588), .B2(new_n223), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n591));
  NAND2_X1  g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n591), .B(new_n592), .Z(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n584), .A2(new_n589), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT21), .B1(new_n580), .B2(new_n581), .ZN(new_n598));
  XNOR2_X1  g397(.A(G127gat), .B(G155gat), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n600), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n601), .A2(new_n280), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n280), .B1(new_n601), .B2(new_n602), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n597), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n594), .A2(new_n605), .A3(new_n596), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610));
  INV_X1    g409(.A(G85gat), .ZN(new_n611));
  OAI21_X1  g410(.A(KEYINPUT7), .B1(new_n611), .B2(new_n497), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT7), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n613), .A2(G85gat), .A3(G92gat), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n612), .A2(new_n614), .B1(new_n611), .B2(new_n497), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT8), .ZN(new_n616));
  NAND2_X1  g415(.A1(G99gat), .A2(G106gat), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT100), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n619), .B1(new_n618), .B2(new_n617), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G99gat), .B(G106gat), .Z(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT101), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n621), .A2(new_n622), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT102), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n258), .A2(new_n260), .A3(new_n628), .ZN(new_n629));
  AND2_X1   g428(.A1(G232gat), .A2(G233gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT41), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n631), .B1(new_n628), .B2(new_n243), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n610), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(KEYINPUT103), .ZN(new_n634));
  XOR2_X1   g433(.A(G134gat), .B(G162gat), .Z(new_n635));
  NOR2_X1   g434(.A1(new_n630), .A2(KEYINPUT41), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  OR3_X1    g437(.A1(new_n629), .A2(new_n610), .A3(new_n632), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n633), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n634), .A2(new_n639), .A3(new_n633), .A4(new_n637), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n609), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G176gat), .B(G204gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT105), .ZN(new_n647));
  XNOR2_X1  g446(.A(G120gat), .B(G148gat), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n647), .B(new_n648), .Z(new_n649));
  NAND2_X1  g448(.A1(G230gat), .A2(G233gat), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n624), .A2(KEYINPUT10), .A3(new_n627), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(new_n579), .B2(new_n582), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n628), .B1(new_n576), .B2(new_n577), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT10), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n625), .A2(KEYINPUT104), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n625), .B1(new_n623), .B2(KEYINPUT104), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n657), .A2(new_n658), .A3(new_n568), .A4(new_n574), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n655), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n651), .B1(new_n654), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n650), .B1(new_n655), .B2(new_n659), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n649), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n655), .A2(new_n656), .A3(new_n659), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n652), .B1(new_n586), .B2(new_n587), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n650), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n662), .ZN(new_n667));
  INV_X1    g466(.A(new_n649), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n663), .A2(new_n669), .A3(KEYINPUT106), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT106), .B1(new_n663), .B2(new_n669), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n645), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n552), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n483), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(G1gat), .ZN(G1324gat));
  INV_X1    g478(.A(new_n518), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT16), .B(G8gat), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n683), .A2(KEYINPUT42), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(KEYINPUT42), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n681), .A2(G8gat), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(G1325gat));
  OAI21_X1  g486(.A(G15gat), .B1(new_n675), .B2(new_n549), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n513), .A2(G15gat), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n688), .B1(new_n675), .B2(new_n689), .ZN(G1326gat));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n676), .A2(new_n691), .A3(new_n333), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT107), .B1(new_n675), .B2(new_n534), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT43), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(G22gat), .ZN(G1327gat));
  NOR3_X1   g495(.A1(new_n673), .A2(new_n609), .A3(new_n643), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n552), .A2(new_n224), .A3(new_n677), .A4(new_n697), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n521), .A2(new_n551), .ZN(new_n702));
  INV_X1    g501(.A(new_n643), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AOI211_X1 g503(.A(KEYINPUT44), .B(new_n643), .C1(new_n521), .C2(new_n551), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n672), .B(KEYINPUT109), .Z(new_n707));
  NAND2_X1  g506(.A1(new_n267), .A2(new_n271), .ZN(new_n708));
  INV_X1    g507(.A(new_n609), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n711), .A2(new_n677), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n700), .B1(new_n712), .B2(new_n224), .ZN(G1328gat));
  NAND4_X1  g512(.A1(new_n552), .A2(new_n225), .A3(new_n680), .A4(new_n697), .ZN(new_n714));
  AND2_X1   g513(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n715));
  NOR2_X1   g514(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n711), .A2(new_n680), .ZN(new_n718));
  OAI221_X1 g517(.A(new_n717), .B1(new_n715), .B2(new_n714), .C1(new_n718), .C2(new_n225), .ZN(G1329gat));
  INV_X1    g518(.A(G43gat), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n552), .A2(new_n720), .A3(new_n548), .A4(new_n697), .ZN(new_n721));
  INV_X1    g520(.A(new_n549), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n711), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n723), .B2(new_n720), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT47), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI211_X1 g525(.A(KEYINPUT47), .B(new_n721), .C1(new_n723), .C2(new_n720), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1330gat));
  NAND3_X1  g527(.A1(new_n706), .A2(new_n333), .A3(new_n710), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT111), .B1(new_n729), .B2(G50gat), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n534), .A2(G50gat), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n552), .A2(new_n697), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(new_n729), .B2(G50gat), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n732), .B(new_n735), .ZN(G1331gat));
  AOI21_X1  g535(.A(new_n708), .B1(new_n521), .B2(new_n551), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n707), .A2(new_n645), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(new_n483), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(new_n564), .ZN(G1332gat));
  INV_X1    g540(.A(KEYINPUT112), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n737), .A2(new_n738), .A3(KEYINPUT112), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n518), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT113), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT113), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n746), .A2(new_n750), .A3(new_n747), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  OR2_X1    g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1333gat));
  OAI21_X1  g553(.A(G71gat), .B1(new_n745), .B2(new_n549), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n513), .A2(G71gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n739), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g557(.A1(new_n746), .A2(new_n333), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g559(.A1(new_n609), .A2(new_n643), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n737), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT51), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(new_n672), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n764), .A2(new_n611), .A3(new_n677), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n609), .A2(new_n672), .A3(new_n708), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n704), .B2(new_n705), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(KEYINPUT114), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n769), .B(new_n766), .C1(new_n704), .C2(new_n705), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n768), .A2(new_n677), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G85gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n765), .A2(new_n772), .ZN(G1336gat));
  NOR4_X1   g572(.A1(new_n763), .A2(G92gat), .A3(new_n518), .A4(new_n707), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(KEYINPUT52), .ZN(new_n775));
  OAI21_X1  g574(.A(G92gat), .B1(new_n767), .B2(new_n518), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n768), .A2(new_n680), .A3(new_n770), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n778), .A2(KEYINPUT115), .A3(G92gat), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT115), .B1(new_n778), .B2(G92gat), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n779), .A2(new_n780), .A3(new_n774), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n777), .B1(new_n781), .B2(new_n782), .ZN(G1337gat));
  INV_X1    g582(.A(G99gat), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n764), .A2(new_n784), .A3(new_n548), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n768), .A2(new_n722), .A3(new_n770), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n786), .B2(new_n784), .ZN(G1338gat));
  OR4_X1    g586(.A1(G106gat), .A2(new_n763), .A3(new_n534), .A4(new_n707), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n789));
  OAI21_X1  g588(.A(G106gat), .B1(new_n767), .B2(new_n534), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n768), .A2(new_n333), .A3(new_n770), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G106gat), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n788), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n791), .B1(new_n794), .B2(new_n789), .ZN(G1339gat));
  INV_X1    g594(.A(new_n669), .ZN(new_n796));
  XOR2_X1   g595(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n797));
  AOI21_X1  g596(.A(new_n668), .B1(new_n661), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n654), .A2(new_n660), .A3(new_n651), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n666), .A2(KEYINPUT54), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n796), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n798), .A2(new_n800), .A3(KEYINPUT55), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n708), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n207), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n246), .A2(new_n249), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n248), .B1(new_n261), .B2(new_n245), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n271), .B(new_n809), .C1(new_n670), .C2(new_n671), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n703), .B1(new_n805), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n801), .A2(new_n802), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(new_n669), .A3(new_n804), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n271), .A2(new_n809), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n813), .A2(new_n643), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n709), .B1(new_n811), .B2(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n272), .A2(new_n609), .A3(new_n672), .A4(new_n643), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n644), .A2(KEYINPUT116), .A3(new_n272), .A4(new_n672), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n816), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n680), .A2(new_n483), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n448), .ZN(new_n824));
  AOI21_X1  g623(.A(G113gat), .B1(new_n824), .B2(new_n708), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n821), .A2(new_n534), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n513), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n821), .A2(KEYINPUT118), .A3(new_n534), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n822), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n272), .A2(new_n342), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n825), .B1(new_n832), .B2(new_n833), .ZN(G1340gat));
  NOR4_X1   g633(.A1(new_n830), .A2(new_n343), .A3(new_n707), .A4(new_n831), .ZN(new_n835));
  AOI21_X1  g634(.A(G120gat), .B1(new_n824), .B2(new_n673), .ZN(new_n836));
  OR3_X1    g635(.A1(new_n835), .A2(new_n836), .A3(KEYINPUT119), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT119), .B1(new_n835), .B2(new_n836), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1341gat));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n337), .A3(new_n609), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n830), .A2(new_n709), .A3(new_n831), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(new_n337), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g643(.A(KEYINPUT120), .B(new_n840), .C1(new_n841), .C2(new_n337), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(G1342gat));
  NAND3_X1  g645(.A1(new_n824), .A2(new_n339), .A3(new_n703), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n847), .A2(KEYINPUT56), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(KEYINPUT56), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n830), .A2(new_n643), .A3(new_n831), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n848), .B(new_n849), .C1(new_n850), .C2(new_n339), .ZN(G1343gat));
  OAI21_X1  g650(.A(new_n810), .B1(new_n272), .B2(new_n813), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n643), .ZN(new_n853));
  INV_X1    g652(.A(new_n815), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n609), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n820), .A2(new_n819), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n534), .A2(KEYINPUT57), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n549), .B(new_n822), .C1(new_n857), .C2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n861), .B1(new_n821), .B2(new_n333), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(G141gat), .B1(new_n863), .B2(new_n272), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT121), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n823), .A2(new_n534), .A3(new_n722), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n297), .A3(new_n708), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n865), .A2(new_n868), .A3(KEYINPUT58), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n864), .B(new_n867), .C1(KEYINPUT121), .C2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(G1344gat));
  NAND3_X1  g671(.A1(new_n866), .A2(new_n298), .A3(new_n673), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n821), .A2(KEYINPUT122), .A3(KEYINPUT57), .A4(new_n333), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n831), .A2(new_n722), .A3(new_n672), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n859), .B1(new_n816), .B2(new_n817), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n333), .B1(new_n855), .B2(new_n856), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(KEYINPUT57), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n875), .B(new_n876), .C1(new_n879), .C2(KEYINPUT122), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n874), .B1(new_n880), .B2(G148gat), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n874), .A2(G148gat), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n860), .A2(new_n862), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(new_n673), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n873), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g686(.A(KEYINPUT123), .B(new_n873), .C1(new_n881), .C2(new_n884), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1345gat));
  OAI21_X1  g688(.A(G155gat), .B1(new_n863), .B2(new_n709), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n866), .A2(new_n305), .A3(new_n609), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1346gat));
  OAI21_X1  g691(.A(G162gat), .B1(new_n863), .B2(new_n643), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n722), .A2(new_n534), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n643), .A2(G162gat), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n821), .A2(new_n822), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT124), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n893), .A2(KEYINPUT125), .A3(new_n897), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1347gat));
  NOR2_X1   g701(.A1(new_n518), .A2(new_n677), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  OR3_X1    g703(.A1(new_n857), .A2(new_n448), .A3(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(G169gat), .B1(new_n906), .B2(new_n708), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n830), .A2(new_n904), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n708), .A2(G169gat), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(G1348gat));
  INV_X1    g709(.A(G176gat), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n906), .A2(new_n911), .A3(new_n673), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n830), .A2(new_n707), .A3(new_n904), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n913), .B2(new_n911), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI211_X1 g715(.A(KEYINPUT126), .B(new_n912), .C1(new_n913), .C2(new_n911), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1349gat));
  NAND2_X1  g717(.A1(new_n366), .A2(KEYINPUT27), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n906), .A2(new_n919), .A3(new_n378), .A4(new_n609), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n830), .A2(new_n709), .A3(new_n904), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n366), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT60), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT60), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n924), .B(new_n920), .C1(new_n921), .C2(new_n366), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1350gat));
  NAND3_X1  g725(.A1(new_n906), .A2(new_n397), .A3(new_n703), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n828), .A2(new_n703), .A3(new_n829), .A4(new_n903), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n928), .A2(new_n929), .A3(G190gat), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n929), .B1(new_n928), .B2(G190gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(G1351gat));
  NOR3_X1   g731(.A1(new_n878), .A2(new_n722), .A3(new_n904), .ZN(new_n933));
  AOI21_X1  g732(.A(G197gat), .B1(new_n933), .B2(new_n708), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n935), .B1(new_n862), .B2(new_n877), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n936), .A2(new_n875), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n722), .A2(new_n904), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n708), .A2(G197gat), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n934), .B1(new_n940), .B2(new_n941), .ZN(G1352gat));
  INV_X1    g741(.A(new_n933), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n943), .A2(G204gat), .A3(new_n672), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT62), .ZN(new_n945));
  OAI21_X1  g744(.A(G204gat), .B1(new_n939), .B2(new_n707), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1353gat));
  NAND4_X1  g746(.A1(new_n936), .A2(new_n609), .A3(new_n875), .A4(new_n938), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT63), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n280), .B1(KEYINPUT127), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n951), .A2(new_n952), .A3(KEYINPUT63), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n948), .B(new_n950), .C1(KEYINPUT127), .C2(new_n949), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n933), .A2(new_n280), .A3(new_n609), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(G1354gat));
  AOI21_X1  g755(.A(G218gat), .B1(new_n933), .B2(new_n703), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n643), .A2(new_n281), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n940), .B2(new_n958), .ZN(G1355gat));
endmodule


