//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040;
  INV_X1    g000(.A(KEYINPUT28), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT0), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n188), .A2(new_n189), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n191), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT64), .B1(new_n192), .B2(G143), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(new_n194), .A3(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  AND4_X1   g016(.A1(KEYINPUT65), .A2(new_n202), .A3(new_n190), .A4(new_n193), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n194), .A2(G146), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n204), .B1(new_n199), .B2(new_n201), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT65), .B1(new_n205), .B2(new_n190), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n198), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT69), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT11), .ZN(new_n210));
  INV_X1    g024(.A(G134), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(G137), .ZN(new_n212));
  INV_X1    g026(.A(G137), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT11), .A3(G134), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(G137), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n212), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G131), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT66), .B(G131), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n218), .A2(new_n212), .A3(new_n214), .A4(new_n215), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  OAI211_X1 g034(.A(KEYINPUT69), .B(new_n198), .C1(new_n203), .C2(new_n206), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n209), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n205), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n225));
  OAI21_X1  g039(.A(G128), .B1(new_n204), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n196), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G131), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n213), .A2(G134), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n229), .B1(new_n230), .B2(new_n215), .ZN(new_n231));
  OR2_X1    g045(.A1(new_n231), .A2(KEYINPUT67), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(KEYINPUT67), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n228), .A2(new_n219), .A3(new_n232), .A4(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G119), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G116), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n237));
  INV_X1    g051(.A(G116), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n237), .B1(new_n238), .B2(G119), .ZN(new_n239));
  NOR3_X1   g053(.A1(new_n235), .A2(KEYINPUT68), .A3(G116), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n236), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  XOR2_X1   g055(.A(KEYINPUT2), .B(G113), .Z(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n242), .B(new_n236), .C1(new_n240), .C2(new_n239), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n234), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n222), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n220), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n234), .B1(new_n207), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n246), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n187), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  XOR2_X1   g069(.A(KEYINPUT26), .B(G101), .Z(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n257));
  XOR2_X1   g071(.A(new_n256), .B(new_n257), .Z(new_n258));
  OR2_X1    g072(.A1(KEYINPUT70), .A2(G237), .ZN(new_n259));
  NAND2_X1  g073(.A1(KEYINPUT70), .A2(G237), .ZN(new_n260));
  AOI21_X1  g074(.A(G953), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G210), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT72), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n262), .A2(KEYINPUT72), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n258), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OR2_X1    g080(.A1(new_n262), .A2(KEYINPUT72), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n256), .B(new_n257), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n263), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n270), .B(KEYINPUT74), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT75), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n222), .A2(new_n273), .A3(new_n234), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n273), .B1(new_n222), .B2(new_n234), .ZN(new_n275));
  NOR3_X1   g089(.A1(new_n274), .A2(new_n275), .A3(new_n246), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n255), .B(new_n272), .C1(new_n276), .C2(KEYINPUT28), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT30), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n252), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n222), .A2(new_n234), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n246), .B(new_n279), .C1(new_n280), .C2(new_n278), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n250), .ZN(new_n282));
  AOI21_X1  g096(.A(KEYINPUT29), .B1(new_n282), .B2(new_n270), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n250), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n247), .B1(new_n222), .B2(new_n234), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT28), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n270), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n288), .A2(KEYINPUT29), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n287), .B(new_n289), .C1(new_n276), .C2(KEYINPUT28), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT77), .ZN(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n246), .B1(new_n280), .B2(KEYINPUT75), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n222), .A2(new_n273), .A3(new_n234), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n187), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT77), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n296), .A2(new_n297), .A3(new_n287), .A4(new_n289), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n284), .A2(new_n291), .A3(new_n292), .A4(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G472), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT28), .B1(new_n293), .B2(new_n294), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n271), .B1(new_n301), .B2(new_n254), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n250), .A2(new_n288), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n250), .A2(KEYINPUT73), .A3(new_n288), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT31), .B1(new_n307), .B2(new_n281), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT73), .B1(new_n250), .B2(new_n288), .ZN(new_n309));
  AOI211_X1 g123(.A(new_n304), .B(new_n270), .C1(new_n222), .C2(new_n249), .ZN(new_n310));
  OAI211_X1 g124(.A(KEYINPUT31), .B(new_n281), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n302), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(G472), .A2(G902), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(KEYINPUT32), .A3(new_n314), .ZN(new_n315));
  XOR2_X1   g129(.A(KEYINPUT76), .B(KEYINPUT32), .Z(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n281), .B1(new_n309), .B2(new_n310), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT31), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n255), .B1(new_n276), .B2(KEYINPUT28), .ZN(new_n321));
  AOI22_X1  g135(.A1(new_n320), .A2(new_n311), .B1(new_n321), .B2(new_n271), .ZN(new_n322));
  INV_X1    g136(.A(new_n314), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n317), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n300), .A2(new_n315), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G469), .ZN(new_n326));
  INV_X1    g140(.A(G953), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G227), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(KEYINPUT84), .ZN(new_n329));
  XNOR2_X1  g143(.A(G110), .B(G140), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n329), .B(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G104), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT3), .B1(new_n333), .B2(G107), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n335));
  INV_X1    g149(.A(G107), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n336), .A3(G104), .ZN(new_n337));
  INV_X1    g151(.A(G101), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n333), .A2(G107), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n334), .A2(new_n337), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n333), .A2(G107), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n336), .A2(G104), .ZN(new_n342));
  OAI21_X1  g156(.A(G101), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n202), .A2(new_n193), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n226), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n344), .B1(new_n346), .B2(new_n224), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT10), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n205), .A2(new_n223), .B1(new_n226), .B2(new_n196), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n344), .A2(KEYINPUT87), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT87), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n340), .A2(new_n343), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n350), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n349), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n334), .A2(new_n337), .A3(new_n339), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT85), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT4), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n334), .A2(new_n337), .A3(KEYINPUT85), .A4(new_n339), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n358), .A2(new_n359), .A3(G101), .A4(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n209), .A2(new_n221), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n358), .A2(G101), .A3(new_n360), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT86), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n340), .A2(KEYINPUT4), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n364), .B1(new_n363), .B2(new_n365), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n355), .B1(new_n362), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n220), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n251), .B(new_n355), .C1(new_n362), .C2(new_n368), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n332), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n344), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n205), .A2(new_n223), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n189), .B1(new_n193), .B2(KEYINPUT1), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n205), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n373), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n350), .A2(new_n344), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(KEYINPUT12), .B1(new_n379), .B2(new_n220), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT12), .ZN(new_n381));
  AOI211_X1 g195(.A(new_n381), .B(new_n251), .C1(new_n377), .C2(new_n378), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT88), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n228), .A2(new_n373), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n220), .B1(new_n384), .B2(new_n347), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n381), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n379), .A2(KEYINPUT12), .A3(new_n220), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT88), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AND4_X1   g203(.A1(new_n371), .A2(new_n383), .A3(new_n332), .A4(new_n389), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n326), .B(new_n292), .C1(new_n372), .C2(new_n390), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n371), .A2(new_n332), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n386), .A2(new_n387), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n371), .A2(new_n393), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n392), .A2(new_n370), .B1(new_n394), .B2(new_n331), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G469), .ZN(new_n396));
  NAND2_X1  g210(.A1(G469), .A2(G902), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n391), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G110), .B(G122), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n246), .A2(new_n361), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n363), .A2(new_n365), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT86), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n401), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n351), .A2(new_n353), .ZN(new_n406));
  OAI211_X1 g220(.A(KEYINPUT5), .B(new_n236), .C1(new_n239), .C2(new_n240), .ZN(new_n407));
  INV_X1    g221(.A(G113), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n238), .A2(G119), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT5), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n245), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n406), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n400), .B1(new_n405), .B2(new_n414), .ZN(new_n415));
  OR2_X1    g229(.A1(new_n406), .A2(new_n413), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n246), .A2(new_n361), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n417), .B1(new_n366), .B2(new_n367), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n418), .A3(new_n399), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n415), .A2(KEYINPUT6), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G125), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n224), .A2(new_n421), .A3(new_n227), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(new_n207), .B2(G125), .ZN(new_n423));
  INV_X1    g237(.A(G224), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(G953), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n423), .B(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n428), .B(new_n400), .C1(new_n405), .C2(new_n414), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n420), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n350), .A2(new_n421), .ZN(new_n431));
  INV_X1    g245(.A(new_n198), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n202), .A2(new_n190), .A3(new_n193), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT65), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n205), .A2(KEYINPUT65), .A3(new_n190), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n432), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n426), .B(new_n431), .C1(new_n437), .C2(new_n421), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT7), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT91), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n426), .B1(new_n440), .B2(KEYINPUT7), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n441), .B1(new_n440), .B2(KEYINPUT7), .ZN(new_n442));
  OAI22_X1  g256(.A1(new_n438), .A2(new_n439), .B1(new_n423), .B2(new_n442), .ZN(new_n443));
  XOR2_X1   g257(.A(new_n399), .B(KEYINPUT8), .Z(new_n444));
  NAND2_X1  g258(.A1(new_n411), .A2(KEYINPUT89), .ZN(new_n445));
  OAI21_X1  g259(.A(G113), .B1(new_n236), .B2(KEYINPUT5), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n445), .A2(new_n407), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(new_n245), .A3(new_n373), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT90), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n450), .A2(new_n451), .B1(new_n413), .B2(new_n344), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n449), .A2(new_n373), .A3(KEYINPUT90), .A4(new_n245), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n444), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n443), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(G902), .B1(new_n455), .B2(new_n419), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n430), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(G210), .B1(G237), .B2(G902), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n430), .A2(new_n456), .A3(new_n458), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(G214), .B1(G237), .B2(G902), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT9), .B(G234), .ZN(new_n464));
  OAI21_X1  g278(.A(G221), .B1(new_n464), .B2(G902), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n398), .A2(new_n462), .A3(new_n463), .A4(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G475), .ZN(new_n467));
  XNOR2_X1  g281(.A(G113), .B(G122), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(new_n333), .ZN(new_n469));
  XNOR2_X1  g283(.A(G125), .B(G140), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n192), .ZN(new_n471));
  NAND2_X1  g285(.A1(KEYINPUT79), .A2(G125), .ZN(new_n472));
  INV_X1    g286(.A(G140), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(KEYINPUT79), .A2(G125), .A3(G140), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(G146), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  AND2_X1   g291(.A1(KEYINPUT70), .A2(G237), .ZN(new_n478));
  NOR2_X1   g292(.A1(KEYINPUT70), .A2(G237), .ZN(new_n479));
  OAI211_X1 g293(.A(G214), .B(new_n327), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT92), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n481), .A2(new_n194), .ZN(new_n482));
  NOR2_X1   g296(.A1(KEYINPUT92), .A2(G143), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n483), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n261), .A2(G214), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(KEYINPUT18), .A2(G131), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n488), .B1(new_n484), .B2(new_n486), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n477), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n484), .A2(new_n486), .A3(new_n218), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n218), .B1(new_n484), .B2(new_n486), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT17), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(KEYINPUT17), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n474), .A2(KEYINPUT16), .A3(new_n475), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT16), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(new_n421), .B2(G140), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n498), .A2(new_n192), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n192), .B1(new_n498), .B2(new_n500), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n469), .B(new_n492), .C1(new_n496), .C2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n484), .A2(new_n486), .ZN(new_n507));
  INV_X1    g321(.A(new_n218), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n510), .A3(new_n493), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n503), .A3(new_n497), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n469), .B1(new_n512), .B2(new_n492), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n292), .B1(new_n506), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n467), .B1(new_n514), .B2(KEYINPUT93), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n492), .B1(new_n496), .B2(new_n504), .ZN(new_n516));
  INV_X1    g330(.A(new_n469), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(G902), .B1(new_n518), .B2(new_n505), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT93), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n502), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT19), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n470), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n474), .A2(KEYINPUT19), .A3(new_n475), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n523), .B1(new_n527), .B2(G146), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(new_n509), .B2(new_n493), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n507), .A2(new_n487), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n530), .A2(new_n489), .B1(new_n471), .B2(new_n476), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n517), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n505), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(G475), .A2(G902), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT20), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n505), .A2(new_n532), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT20), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n538), .A3(new_n534), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n189), .A2(G143), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n194), .A2(G128), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n541), .A2(new_n542), .A3(G134), .ZN(new_n543));
  XOR2_X1   g357(.A(G116), .B(G122), .Z(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(G107), .ZN(new_n545));
  XNOR2_X1  g359(.A(G116), .B(G122), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n336), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n543), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT94), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n194), .A2(G128), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT13), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n549), .B(new_n550), .C1(new_n542), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n189), .A2(G143), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n541), .B1(KEYINPUT13), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT94), .B1(new_n550), .B2(new_n551), .ZN(new_n555));
  OAI211_X1 g369(.A(G134), .B(new_n552), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n548), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n238), .A2(KEYINPUT14), .A3(G122), .ZN(new_n558));
  OAI211_X1 g372(.A(G107), .B(new_n558), .C1(new_n544), .C2(KEYINPUT14), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n211), .B1(new_n550), .B2(new_n553), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n559), .B(new_n547), .C1(new_n543), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(G217), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n464), .A2(new_n563), .A3(G953), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT95), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT95), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n557), .A2(new_n561), .A3(new_n567), .A4(new_n564), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n562), .A2(new_n565), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n292), .ZN(new_n571));
  INV_X1    g385(.A(G478), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(KEYINPUT15), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(G952), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(G953), .ZN(new_n576));
  INV_X1    g390(.A(G234), .ZN(new_n577));
  INV_X1    g391(.A(G237), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT21), .B(G898), .ZN(new_n580));
  XOR2_X1   g394(.A(new_n580), .B(KEYINPUT96), .Z(new_n581));
  AOI211_X1 g395(.A(new_n292), .B(new_n327), .C1(G234), .C2(G237), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n579), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n573), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n570), .A2(new_n292), .A3(new_n585), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n574), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n522), .A2(new_n540), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n466), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT78), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n590), .B1(new_n189), .B2(G119), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n235), .A2(KEYINPUT78), .A3(G128), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n189), .A2(G119), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT24), .B(G110), .ZN(new_n595));
  OR2_X1    g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT23), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n235), .A2(G128), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n189), .A2(KEYINPUT23), .A3(G119), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(G110), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n596), .B(new_n602), .C1(new_n501), .C2(new_n502), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n594), .A2(new_n595), .ZN(new_n604));
  INV_X1    g418(.A(G110), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n598), .A2(new_n600), .A3(new_n605), .A4(new_n599), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n604), .A2(KEYINPUT80), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(new_n523), .A3(new_n471), .ZN(new_n608));
  AOI21_X1  g422(.A(KEYINPUT80), .B1(new_n604), .B2(new_n606), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n603), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT22), .B(G137), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n327), .A2(G221), .A3(G234), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n603), .B(new_n613), .C1(new_n608), .C2(new_n609), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n292), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT81), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT25), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n617), .A2(KEYINPUT81), .A3(KEYINPUT25), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n563), .B1(G234), .B2(new_n292), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT82), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n620), .A2(KEYINPUT82), .A3(new_n621), .A4(new_n622), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n622), .A2(G902), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT83), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n615), .A2(new_n616), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n625), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n325), .A2(new_n589), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G101), .ZN(G3));
  NOR2_X1   g447(.A1(new_n322), .A2(new_n323), .ZN(new_n634));
  OAI21_X1  g448(.A(G472), .B1(new_n322), .B2(G902), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n634), .B1(new_n635), .B2(KEYINPUT97), .ZN(new_n636));
  INV_X1    g450(.A(G472), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n313), .B2(new_n292), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT97), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n398), .A2(new_n465), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n641), .A2(new_n630), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n462), .A2(new_n463), .A3(new_n584), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT33), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n557), .A2(new_n561), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n565), .A2(KEYINPUT98), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT99), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n647), .B1(new_n557), .B2(new_n561), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n648), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n647), .ZN(new_n653));
  OAI21_X1  g467(.A(KEYINPUT33), .B1(new_n562), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(KEYINPUT99), .B1(new_n654), .B2(new_n650), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n652), .A2(new_n655), .B1(new_n570), .B2(new_n645), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n572), .A2(G902), .ZN(new_n657));
  AOI22_X1  g471(.A1(new_n656), .A2(new_n657), .B1(new_n572), .B2(new_n571), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n658), .B1(new_n522), .B2(new_n540), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n644), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n643), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G104), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  NAND2_X1  g479(.A1(new_n574), .A2(new_n586), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n536), .A2(KEYINPUT101), .A3(new_n539), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n538), .B1(new_n537), .B2(new_n534), .ZN(new_n669));
  AOI211_X1 g483(.A(KEYINPUT20), .B(new_n535), .C1(new_n505), .C2(new_n532), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n522), .A2(new_n666), .A3(new_n667), .A4(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n644), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n643), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT35), .B(G107), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  NOR2_X1   g490(.A1(new_n614), .A2(KEYINPUT36), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n610), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n628), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n625), .A2(new_n626), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(KEYINPUT103), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n625), .A2(new_n684), .A3(new_n681), .A4(new_n626), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n466), .ZN(new_n687));
  INV_X1    g501(.A(new_n588), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n687), .A2(new_n636), .A3(new_n688), .A4(new_n640), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT37), .B(G110), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G12));
  AND2_X1   g507(.A1(new_n687), .A2(new_n325), .ZN(new_n694));
  INV_X1    g508(.A(G900), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n582), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n579), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n672), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G128), .ZN(G30));
  INV_X1    g515(.A(new_n465), .ZN(new_n702));
  OAI21_X1  g516(.A(G469), .B1(new_n395), .B2(G902), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n702), .B1(new_n703), .B2(new_n391), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n697), .B(KEYINPUT39), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n706), .B(KEYINPUT40), .Z(new_n707));
  INV_X1    g521(.A(new_n318), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n285), .A2(new_n286), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n272), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n292), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G472), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n324), .A2(new_n315), .A3(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT38), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n462), .B(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n463), .ZN(new_n716));
  OAI21_X1  g530(.A(G475), .B1(new_n519), .B2(new_n520), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n514), .A2(KEYINPUT93), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n540), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n666), .ZN(new_n720));
  NOR4_X1   g534(.A1(new_n715), .A2(new_n716), .A3(new_n682), .A4(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n707), .A2(new_n713), .A3(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(new_n722), .B(KEYINPUT106), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G143), .ZN(G45));
  AOI211_X1 g538(.A(new_n698), .B(new_n658), .C1(new_n522), .C2(new_n540), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n694), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G146), .ZN(G48));
  OAI21_X1  g541(.A(new_n292), .B1(new_n372), .B2(new_n390), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(G469), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(KEYINPUT107), .A3(new_n391), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n728), .A2(new_n731), .A3(G469), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n702), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n325), .A2(new_n631), .A3(new_n661), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT41), .B(G113), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G15));
  NAND4_X1  g550(.A1(new_n325), .A2(new_n631), .A3(new_n673), .A4(new_n733), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G116), .ZN(G18));
  AND3_X1   g552(.A1(new_n430), .A2(new_n456), .A3(new_n458), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n458), .B1(new_n430), .B2(new_n456), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n463), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI211_X1 g555(.A(new_n702), .B(new_n741), .C1(new_n730), .C2(new_n732), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n683), .A2(new_n688), .A3(new_n685), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n325), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G119), .ZN(G21));
  NAND2_X1  g559(.A1(new_n296), .A2(new_n287), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n271), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n320), .A2(new_n311), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n323), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n638), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n644), .A2(new_n720), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n750), .A2(new_n751), .A3(new_n733), .A4(new_n631), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G122), .ZN(G24));
  INV_X1    g567(.A(new_n658), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n719), .A2(new_n754), .A3(new_n697), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n625), .A2(new_n626), .A3(new_n681), .ZN(new_n756));
  NOR4_X1   g570(.A1(new_n638), .A2(new_n749), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n742), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G125), .ZN(G27));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT42), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT32), .ZN(new_n762));
  AOI211_X1 g576(.A(new_n762), .B(new_n323), .C1(new_n748), .C2(new_n302), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT32), .B1(new_n313), .B2(new_n314), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n630), .B1(new_n765), .B2(new_n300), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n739), .A2(new_n740), .A3(new_n716), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n725), .A2(new_n704), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n761), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n325), .A2(new_n768), .A3(new_n761), .A4(new_n631), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n760), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n762), .B1(new_n322), .B2(new_n323), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n315), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n299), .A2(G472), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n768), .B(new_n631), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT42), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(KEYINPUT108), .A3(new_n770), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n772), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(new_n229), .ZN(G33));
  NAND2_X1  g594(.A1(new_n704), .A2(new_n767), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n325), .A2(new_n631), .A3(new_n699), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  INV_X1    g598(.A(new_n391), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n395), .A2(KEYINPUT45), .ZN(new_n786));
  XOR2_X1   g600(.A(new_n786), .B(KEYINPUT110), .Z(new_n787));
  INV_X1    g601(.A(new_n395), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n326), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n790), .A2(KEYINPUT109), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(KEYINPUT109), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n787), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n397), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT46), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n785), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n796), .B1(new_n795), .B2(new_n794), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n465), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n799), .A2(new_n705), .ZN(new_n800));
  INV_X1    g614(.A(new_n719), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(KEYINPUT43), .A3(new_n754), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n802), .A2(KEYINPUT112), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(KEYINPUT112), .ZN(new_n804));
  XOR2_X1   g618(.A(new_n658), .B(KEYINPUT111), .Z(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n719), .ZN(new_n806));
  OAI22_X1  g620(.A1(new_n803), .A2(new_n804), .B1(KEYINPUT43), .B2(new_n806), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n641), .A2(KEYINPUT113), .A3(new_n682), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT113), .B1(new_n641), .B2(new_n682), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT44), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n800), .A2(new_n767), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G137), .ZN(G39));
  INV_X1    g629(.A(new_n767), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n325), .A2(new_n631), .A3(new_n755), .A4(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n797), .A2(KEYINPUT47), .A3(new_n465), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT47), .B1(new_n797), .B2(new_n465), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G140), .ZN(G42));
  INV_X1    g635(.A(new_n579), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n807), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n750), .A2(new_n631), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(new_n816), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT118), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n818), .A2(new_n819), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n730), .A2(new_n732), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n702), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n828), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n733), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(new_n816), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n823), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n750), .A2(new_n682), .ZN(new_n836));
  INV_X1    g650(.A(new_n713), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n834), .A2(new_n631), .A3(new_n822), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n801), .A2(new_n658), .ZN(new_n839));
  OAI22_X1  g653(.A1(new_n835), .A2(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT50), .ZN(new_n841));
  INV_X1    g655(.A(new_n715), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n842), .A2(new_n833), .A3(new_n463), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n841), .B1(new_n826), .B2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n823), .A2(KEYINPUT50), .A3(new_n825), .A4(new_n843), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n840), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT51), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n832), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n823), .A2(new_n766), .A3(new_n834), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n850), .B(KEYINPUT48), .Z(new_n851));
  INV_X1    g665(.A(new_n742), .ZN(new_n852));
  OAI221_X1 g666(.A(new_n576), .B1(new_n660), .B2(new_n838), .C1(new_n826), .C2(new_n852), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n849), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  AND4_X1   g668(.A1(new_n734), .A2(new_n737), .A3(new_n744), .A4(new_n752), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n540), .B(new_n666), .C1(new_n718), .C2(new_n717), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n857), .A2(new_n659), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n644), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n642), .A2(new_n630), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n636), .A2(new_n859), .A3(new_n860), .A4(new_n640), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n689), .A2(new_n861), .A3(new_n632), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n667), .A2(new_n671), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n570), .A2(new_n292), .A3(new_n585), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n585), .B1(new_n570), .B2(new_n292), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n864), .A2(new_n865), .A3(new_n698), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n866), .B1(new_n717), .B2(new_n718), .ZN(new_n867));
  OAI21_X1  g681(.A(KEYINPUT114), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n574), .A2(new_n586), .A3(new_n697), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n515), .B2(new_n521), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT114), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n870), .A2(new_n871), .A3(new_n667), .A4(new_n671), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n683), .A2(new_n868), .A3(new_n872), .A4(new_n685), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n699), .A2(new_n631), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n325), .ZN(new_n876));
  INV_X1    g690(.A(new_n757), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n782), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n855), .A2(new_n862), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT115), .B1(new_n779), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n734), .A2(new_n737), .A3(new_n744), .A4(new_n752), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n781), .B1(new_n876), .B2(new_n877), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n689), .A2(new_n861), .A3(new_n632), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT115), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n885), .A2(new_n886), .A3(new_n772), .A4(new_n778), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n687), .B(new_n325), .C1(new_n699), .C2(new_n725), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n720), .A2(new_n741), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n698), .A2(KEYINPUT116), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n698), .A2(KEYINPUT116), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n682), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n713), .A2(new_n704), .A3(new_n889), .A4(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n888), .A2(new_n893), .A3(new_n758), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT52), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT52), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n888), .A2(new_n758), .A3(new_n896), .A4(new_n893), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n881), .A2(new_n887), .A3(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT53), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n899), .B(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT54), .ZN(new_n902));
  INV_X1    g716(.A(new_n818), .ZN(new_n903));
  INV_X1    g717(.A(new_n819), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n903), .A2(KEYINPUT119), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT119), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(new_n818), .B2(new_n819), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n905), .A2(new_n907), .A3(new_n831), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n847), .B1(new_n908), .B2(new_n828), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT51), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n899), .A2(new_n900), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT54), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n883), .A2(new_n884), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n777), .A2(KEYINPUT53), .A3(new_n770), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n914), .A2(new_n915), .A3(new_n855), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n895), .A2(new_n897), .ZN(new_n917));
  OAI21_X1  g731(.A(KEYINPUT117), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT117), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n898), .A2(new_n919), .A3(new_n885), .A4(new_n915), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n912), .A2(new_n913), .A3(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n854), .A2(new_n902), .A3(new_n911), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n575), .A2(new_n327), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n801), .A2(new_n463), .A3(new_n465), .A4(new_n754), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n842), .A2(new_n630), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n830), .B(KEYINPUT49), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n927), .A2(new_n837), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n925), .A2(new_n929), .ZN(G75));
  NAND2_X1  g744(.A1(new_n420), .A2(new_n429), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(new_n427), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT55), .Z(new_n933));
  AOI22_X1  g747(.A1(new_n899), .A2(new_n900), .B1(new_n918), .B2(new_n920), .ZN(new_n934));
  INV_X1    g748(.A(G210), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n934), .A2(new_n935), .A3(new_n292), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n933), .B1(new_n936), .B2(KEYINPUT56), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n327), .A2(G952), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT120), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n934), .B2(new_n292), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n914), .A2(new_n772), .A3(new_n778), .A4(new_n855), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n917), .B1(new_n943), .B2(KEYINPUT115), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT53), .B1(new_n944), .B2(new_n887), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n918), .A2(new_n920), .ZN(new_n946));
  OAI211_X1 g760(.A(KEYINPUT120), .B(G902), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n942), .A2(new_n459), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n933), .A2(KEYINPUT56), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n940), .B1(new_n948), .B2(new_n949), .ZN(G51));
  INV_X1    g764(.A(new_n793), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n942), .A2(new_n951), .A3(new_n947), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT121), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n372), .A2(new_n390), .ZN(new_n954));
  OAI21_X1  g768(.A(KEYINPUT54), .B1(new_n945), .B2(new_n946), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n922), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n397), .B(KEYINPUT57), .Z(new_n957));
  AOI21_X1  g771(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n952), .B1(new_n953), .B2(new_n958), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n956), .A2(new_n957), .ZN(new_n960));
  OAI21_X1  g774(.A(KEYINPUT121), .B1(new_n960), .B2(new_n954), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n938), .B1(new_n959), .B2(new_n961), .ZN(G54));
  NAND2_X1  g776(.A1(KEYINPUT58), .A2(G475), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT122), .Z(new_n964));
  NAND3_X1  g778(.A1(new_n942), .A2(new_n947), .A3(new_n964), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n965), .A2(new_n533), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n533), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n966), .A2(new_n967), .A3(new_n938), .ZN(G60));
  NAND2_X1  g782(.A1(new_n902), .A2(new_n922), .ZN(new_n969));
  NAND2_X1  g783(.A1(G478), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT59), .Z(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n656), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n956), .A2(new_n656), .A3(new_n972), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n973), .A2(new_n938), .A3(new_n974), .ZN(G63));
  INV_X1    g789(.A(KEYINPUT61), .ZN(new_n976));
  NAND2_X1  g790(.A1(G217), .A2(G902), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT60), .ZN(new_n978));
  OAI21_X1  g792(.A(KEYINPUT123), .B1(new_n934), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n615), .A2(new_n616), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT123), .ZN(new_n981));
  INV_X1    g795(.A(new_n978), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n981), .B(new_n982), .C1(new_n945), .C2(new_n946), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n979), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n939), .ZN(new_n985));
  INV_X1    g799(.A(new_n678), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n986), .B1(new_n979), .B2(new_n983), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n976), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n987), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n989), .A2(KEYINPUT61), .A3(new_n939), .A4(new_n984), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n988), .A2(new_n990), .ZN(G66));
  INV_X1    g805(.A(new_n581), .ZN(new_n992));
  OAI21_X1  g806(.A(G953), .B1(new_n992), .B2(new_n424), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n882), .A2(new_n884), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n993), .B1(new_n994), .B2(G953), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n931), .B1(G898), .B2(new_n327), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n995), .B(new_n996), .ZN(G69));
  INV_X1    g811(.A(G227), .ZN(new_n998));
  OAI21_X1  g812(.A(G953), .B1(new_n998), .B2(new_n695), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT126), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n279), .B1(new_n280), .B2(new_n278), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT124), .Z(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(new_n527), .Z(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(new_n779), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n799), .A2(new_n705), .A3(new_n766), .A4(new_n889), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n888), .A2(new_n758), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n1007), .A2(new_n783), .ZN(new_n1008));
  AND4_X1   g822(.A1(new_n1005), .A2(new_n820), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(G953), .B1(new_n1009), .B2(new_n814), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n327), .A2(G900), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1004), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT125), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n723), .A2(new_n1007), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1014), .B1(new_n1015), .B2(KEYINPUT62), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT62), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n723), .A2(KEYINPUT125), .A3(new_n1017), .A4(new_n1007), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n325), .A2(new_n631), .ZN(new_n1020));
  NOR4_X1   g834(.A1(new_n1020), .A2(new_n706), .A3(new_n816), .A4(new_n858), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1021), .B1(new_n1015), .B2(KEYINPUT62), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1019), .A2(new_n814), .A3(new_n820), .A4(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1004), .B1(new_n1023), .B2(new_n327), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1000), .B1(new_n1013), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1000), .ZN(new_n1026));
  AND2_X1   g840(.A1(new_n1023), .A2(new_n327), .ZN(new_n1027));
  OAI211_X1 g841(.A(new_n1012), .B(new_n1026), .C1(new_n1027), .C2(new_n1004), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1025), .A2(new_n1028), .ZN(G72));
  NAND2_X1  g843(.A1(G472), .A2(G902), .ZN(new_n1030));
  XOR2_X1   g844(.A(new_n1030), .B(KEYINPUT63), .Z(new_n1031));
  INV_X1    g845(.A(new_n994), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1031), .B1(new_n1023), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1033), .A2(new_n288), .A3(new_n282), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1009), .A2(new_n814), .A3(new_n994), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1035), .A2(new_n1031), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n282), .A2(new_n288), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n938), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n288), .B1(new_n281), .B2(new_n250), .ZN(new_n1039));
  OAI211_X1 g853(.A(new_n901), .B(new_n1031), .C1(new_n708), .C2(new_n1039), .ZN(new_n1040));
  AND3_X1   g854(.A1(new_n1034), .A2(new_n1038), .A3(new_n1040), .ZN(G57));
endmodule


