//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 1 1 1 1 1 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  XNOR2_X1  g000(.A(KEYINPUT2), .B(G113), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G116), .B(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n189), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(new_n187), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT67), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G134), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT67), .A3(G137), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(KEYINPUT66), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT66), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G137), .ZN(new_n202));
  AND2_X1   g016(.A1(KEYINPUT11), .A2(G134), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT11), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n205), .B1(new_n197), .B2(G137), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n199), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G131), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n199), .A2(new_n204), .A3(new_n209), .A4(new_n206), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT64), .A2(G146), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(G143), .A3(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n213), .A2(G143), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(KEYINPUT0), .A2(G128), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT65), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n216), .A2(new_n222), .A3(new_n218), .A4(new_n219), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  OR2_X1    g039(.A1(new_n219), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G143), .ZN(new_n227));
  AND2_X1   g041(.A1(KEYINPUT64), .A2(G146), .ZN(new_n228));
  NOR2_X1   g042(.A1(KEYINPUT64), .A2(G146), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n213), .A2(G143), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n226), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n211), .A2(new_n224), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G128), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(KEYINPUT1), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n216), .A2(new_n218), .A3(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n230), .A2(new_n231), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n235), .B1(new_n216), .B2(KEYINPUT1), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(G134), .B1(new_n200), .B2(new_n202), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n197), .A2(G137), .ZN(new_n242));
  OAI21_X1  g056(.A(G131), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(new_n210), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT30), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n234), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(new_n210), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT68), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n243), .A2(new_n210), .A3(KEYINPUT68), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n240), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n245), .B1(new_n252), .B2(new_n234), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n193), .B1(new_n247), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n193), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n252), .A2(new_n255), .A3(new_n234), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT69), .B(G953), .ZN(new_n257));
  INV_X1    g071(.A(G237), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(G210), .A3(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n259), .B(KEYINPUT71), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G101), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n260), .B(new_n263), .Z(new_n264));
  NAND3_X1  g078(.A1(new_n254), .A2(new_n256), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT31), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n256), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n230), .A2(new_n231), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT1), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n228), .A2(new_n229), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n270), .B1(new_n271), .B2(G143), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n269), .B1(new_n272), .B2(new_n235), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n249), .A2(new_n248), .B1(new_n273), .B2(new_n237), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n232), .B1(new_n221), .B2(new_n223), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n274), .A2(new_n251), .B1(new_n275), .B2(new_n211), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n246), .B1(new_n276), .B2(new_n245), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n268), .B1(new_n277), .B2(new_n193), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(KEYINPUT31), .A3(new_n264), .ZN(new_n279));
  INV_X1    g093(.A(new_n264), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT28), .B1(new_n276), .B2(new_n255), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n234), .A2(new_n244), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n193), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n252), .A2(KEYINPUT28), .A3(new_n255), .A4(new_n234), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n280), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT28), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n256), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(new_n284), .A3(new_n283), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(KEYINPUT72), .A3(new_n280), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n267), .A2(new_n279), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(G472), .A2(G902), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(KEYINPUT32), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT31), .B1(new_n278), .B2(new_n264), .ZN(new_n297));
  AND4_X1   g111(.A1(KEYINPUT31), .A2(new_n254), .A3(new_n256), .A4(new_n264), .ZN(new_n298));
  INV_X1    g112(.A(new_n292), .ZN(new_n299));
  AOI21_X1  g113(.A(KEYINPUT72), .B1(new_n291), .B2(new_n280), .ZN(new_n300));
  OAI22_X1  g114(.A1(new_n297), .A2(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT32), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n302), .A3(new_n294), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n296), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n278), .A2(new_n280), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n291), .A2(new_n264), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT29), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  XOR2_X1   g121(.A(KEYINPUT74), .B(G902), .Z(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n281), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n255), .B1(new_n252), .B2(new_n234), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT28), .B1(new_n268), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n290), .A2(KEYINPUT73), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n264), .A2(KEYINPUT29), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n309), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(G472), .B1(new_n307), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n304), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n321));
  INV_X1    g135(.A(G140), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n321), .B1(G125), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT76), .B(G125), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(new_n322), .ZN(new_n325));
  AND2_X1   g139(.A1(KEYINPUT76), .A2(G125), .ZN(new_n326));
  NOR2_X1   g140(.A1(KEYINPUT76), .A2(G125), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(new_n321), .A3(G140), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n320), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n328), .A2(KEYINPUT16), .A3(G140), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n213), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G125), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT77), .B1(new_n333), .B2(G140), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n334), .B1(new_n328), .B2(G140), .ZN(new_n335));
  NOR4_X1   g149(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT77), .A4(new_n322), .ZN(new_n336));
  OAI21_X1  g150(.A(KEYINPUT16), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n331), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(G146), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT23), .ZN(new_n341));
  INV_X1    g155(.A(G119), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n341), .B1(new_n342), .B2(G128), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n235), .A2(KEYINPUT23), .A3(G119), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(G128), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT75), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT75), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n343), .A2(new_n344), .A3(new_n348), .A4(new_n345), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(G110), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n235), .A2(G119), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n345), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT24), .B(G110), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n350), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n340), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(G125), .B(G140), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n271), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n352), .A2(new_n353), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n359), .B1(G110), .B2(new_n346), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n339), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n257), .A2(G221), .A3(G234), .ZN(new_n362));
  XOR2_X1   g176(.A(KEYINPUT22), .B(G137), .Z(new_n363));
  OR2_X1    g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n363), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n356), .A2(new_n361), .A3(new_n366), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n364), .A2(KEYINPUT78), .A3(new_n365), .ZN(new_n368));
  AOI21_X1  g182(.A(KEYINPUT78), .B1(new_n364), .B2(new_n365), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n354), .B1(new_n332), .B2(new_n339), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n360), .A2(new_n358), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n330), .A2(new_n331), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n372), .B1(new_n373), .B2(G146), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n370), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n367), .A2(new_n375), .A3(new_n309), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT79), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT25), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G217), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(new_n309), .B2(G234), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n376), .A2(new_n378), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n367), .A2(new_n375), .A3(KEYINPUT25), .A4(new_n309), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(KEYINPUT79), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n381), .A2(G902), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n367), .A2(new_n375), .A3(new_n387), .ZN(new_n388));
  XOR2_X1   g202(.A(new_n388), .B(KEYINPUT80), .Z(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n319), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT94), .B(G475), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n325), .A2(new_n329), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n358), .B1(new_n395), .B2(new_n213), .ZN(new_n396));
  INV_X1    g210(.A(G953), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT69), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT69), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G953), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n398), .A2(new_n400), .A3(G214), .A4(new_n258), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n227), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n257), .A2(G143), .A3(G214), .A4(new_n258), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(KEYINPUT18), .A3(G131), .ZN(new_n405));
  NAND2_X1  g219(.A1(KEYINPUT18), .A2(G131), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n402), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n396), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT17), .ZN(new_n409));
  AOI211_X1 g223(.A(new_n409), .B(new_n209), .C1(new_n402), .C2(new_n403), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n404), .A2(G131), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n402), .A2(new_n403), .A3(new_n209), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n410), .B1(new_n413), .B2(KEYINPUT93), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n404), .A2(KEYINPUT93), .A3(KEYINPUT17), .A4(G131), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n332), .A2(new_n339), .A3(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n408), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT95), .ZN(new_n418));
  XNOR2_X1  g232(.A(G113), .B(G122), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(G104), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT95), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n421), .B(new_n408), .C1(new_n414), .C2(new_n416), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n418), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT96), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n420), .B(KEYINPUT92), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n408), .B(new_n426), .C1(new_n414), .C2(new_n416), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n418), .A2(KEYINPUT96), .A3(new_n420), .A4(new_n422), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n425), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G902), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n394), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(G116), .B(G122), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(KEYINPUT97), .ZN(new_n433));
  INV_X1    g247(.A(G107), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(G128), .B(G143), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(new_n197), .ZN(new_n438));
  INV_X1    g252(.A(G116), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(KEYINPUT14), .A3(G122), .ZN(new_n440));
  INV_X1    g254(.A(new_n432), .ZN(new_n441));
  OAI211_X1 g255(.A(G107), .B(new_n440), .C1(new_n441), .C2(KEYINPUT14), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT98), .B1(new_n436), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n437), .A2(KEYINPUT13), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n235), .A2(KEYINPUT13), .A3(G143), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(new_n197), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n445), .A2(new_n447), .B1(new_n197), .B2(new_n437), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n433), .A2(new_n434), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n448), .B1(new_n436), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT98), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n435), .A2(new_n451), .A3(new_n438), .A4(new_n442), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n444), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT9), .B(G234), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(KEYINPUT81), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(G217), .A3(new_n397), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n456), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n444), .A2(new_n450), .A3(new_n452), .A4(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n308), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G478), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(KEYINPUT15), .ZN(new_n462));
  XOR2_X1   g276(.A(new_n460), .B(new_n462), .Z(new_n463));
  INV_X1    g277(.A(KEYINPUT19), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n357), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n465), .B1(new_n395), .B2(new_n464), .ZN(new_n466));
  INV_X1    g280(.A(new_n271), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n339), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n411), .A2(new_n412), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n408), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n420), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n427), .ZN(new_n472));
  INV_X1    g286(.A(G475), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n473), .A3(new_n430), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT20), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n431), .A2(new_n463), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(G214), .B1(G237), .B2(G902), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n273), .A2(new_n328), .A3(new_n237), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n275), .A2(new_n328), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT88), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n397), .A2(G224), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n485), .B(KEYINPUT89), .Z(new_n486));
  OAI21_X1  g300(.A(KEYINPUT88), .B1(new_n275), .B2(new_n328), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n484), .A2(KEYINPUT7), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n217), .B1(new_n271), .B2(G143), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n222), .B1(new_n489), .B2(new_n219), .ZN(new_n490));
  INV_X1    g304(.A(new_n223), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n233), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n483), .A3(new_n324), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(new_n487), .A3(new_n480), .ZN(new_n494));
  INV_X1    g308(.A(new_n486), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT7), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G104), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT3), .B1(new_n499), .B2(G107), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT3), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n434), .A3(G104), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n499), .A2(G107), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT4), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n505), .A3(G101), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT83), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT83), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n504), .A2(new_n508), .A3(new_n505), .A4(G101), .ZN(new_n509));
  INV_X1    g323(.A(G101), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n500), .A2(new_n502), .A3(new_n510), .A4(new_n503), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n511), .A2(KEYINPUT4), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n504), .A2(G101), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n507), .A2(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n499), .A2(G107), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n434), .A2(G104), .ZN(new_n516));
  OAI21_X1  g330(.A(G101), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(G113), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT87), .B(KEYINPUT5), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n439), .A2(G119), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT5), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT87), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT87), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT5), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n189), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n523), .A2(new_n529), .B1(new_n189), .B2(new_n188), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n514), .A2(new_n193), .B1(new_n519), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(G110), .B(G122), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n523), .A2(new_n529), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n190), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT91), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n535), .A3(new_n518), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT91), .B1(new_n530), .B2(new_n519), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n523), .B1(new_n524), .B2(new_n191), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(new_n519), .A3(new_n190), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n532), .B(KEYINPUT8), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n531), .A2(new_n532), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n488), .A2(new_n496), .A3(new_n498), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n430), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT90), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n507), .A2(new_n509), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n512), .A2(new_n513), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n193), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n530), .A2(new_n519), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n550), .A3(new_n532), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT6), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n532), .B1(new_n549), .B2(new_n550), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n531), .A2(KEYINPUT6), .A3(new_n532), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n493), .A2(new_n487), .A3(new_n486), .A4(new_n480), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n496), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n546), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n552), .A2(new_n553), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n549), .A2(new_n550), .ZN(new_n561));
  INV_X1    g375(.A(new_n532), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(KEYINPUT6), .A3(new_n551), .ZN(new_n564));
  AND4_X1   g378(.A1(new_n546), .A2(new_n558), .A3(new_n560), .A4(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n545), .B1(new_n559), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G210), .B1(G237), .B2(G902), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n564), .A2(new_n560), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n486), .B1(new_n484), .B2(new_n487), .ZN(new_n571));
  INV_X1    g385(.A(new_n557), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT90), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n558), .A2(new_n546), .A3(new_n560), .A4(new_n564), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(new_n567), .A3(new_n545), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n479), .B1(new_n569), .B2(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n397), .A2(G952), .ZN(new_n579));
  INV_X1    g393(.A(G234), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n579), .B1(new_n580), .B2(new_n258), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n257), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n583), .B(new_n308), .C1(new_n580), .C2(new_n258), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(KEYINPUT99), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT21), .B(G898), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n582), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n455), .A2(new_n430), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n589), .A2(G221), .ZN(new_n590));
  INV_X1    g404(.A(G469), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(new_n430), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n257), .A2(G227), .ZN(new_n593));
  XOR2_X1   g407(.A(G110), .B(G140), .Z(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n275), .A2(new_n547), .A3(new_n548), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT84), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n514), .A2(KEYINPUT84), .A3(new_n275), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n211), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n216), .A2(new_n218), .A3(new_n236), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT1), .B1(new_n227), .B2(G146), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n216), .A2(new_n218), .B1(G128), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT85), .B1(new_n605), .B2(new_n518), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n235), .B1(new_n231), .B2(KEYINPUT1), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n237), .B1(new_n489), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT85), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n610), .A3(new_n519), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n606), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n240), .ZN(new_n613));
  OAI21_X1  g427(.A(KEYINPUT10), .B1(new_n613), .B2(new_n518), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n600), .A2(new_n601), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n601), .B1(new_n600), .B2(new_n615), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n595), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g432(.A1(new_n598), .A2(new_n599), .B1(new_n612), .B2(new_n614), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n595), .B1(new_n619), .B2(new_n601), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT12), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n606), .A2(new_n611), .B1(new_n613), .B2(new_n518), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n621), .B1(new_n622), .B2(new_n601), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n609), .A2(new_n610), .A3(new_n519), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n610), .B1(new_n609), .B2(new_n519), .ZN(new_n625));
  OAI22_X1  g439(.A1(new_n624), .A2(new_n625), .B1(new_n240), .B2(new_n519), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n626), .A2(KEYINPUT12), .A3(new_n211), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n620), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n308), .B1(new_n618), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n592), .B1(new_n630), .B2(new_n591), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n595), .B(KEYINPUT82), .ZN(new_n632));
  INV_X1    g446(.A(new_n628), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n632), .B1(new_n633), .B2(new_n616), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n600), .A2(new_n615), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n211), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n600), .A2(new_n601), .A3(new_n615), .ZN(new_n637));
  INV_X1    g451(.A(new_n595), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n636), .B1(new_n639), .B2(KEYINPUT86), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT86), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n620), .A2(new_n641), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n634), .B(G469), .C1(new_n640), .C2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n590), .B1(new_n631), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n477), .A2(new_n578), .A3(new_n588), .A4(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n392), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(new_n510), .ZN(G3));
  NOR2_X1   g461(.A1(new_n293), .A2(new_n295), .ZN(new_n648));
  OAI21_X1  g462(.A(G472), .B1(new_n293), .B2(new_n308), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT100), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI211_X1 g465(.A(KEYINPUT100), .B(G472), .C1(new_n293), .C2(new_n308), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n651), .A2(new_n644), .A3(new_n391), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT102), .B(G478), .ZN(new_n654));
  OR3_X1    g468(.A1(new_n460), .A2(KEYINPUT103), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT103), .B1(new_n460), .B2(new_n654), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT101), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT33), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n457), .B2(new_n459), .ZN(new_n660));
  NOR2_X1   g474(.A1(KEYINPUT101), .A2(KEYINPUT33), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n457), .A2(new_n657), .A3(new_n658), .A4(new_n459), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n308), .A2(new_n461), .ZN(new_n666));
  AOI22_X1  g480(.A1(new_n655), .A2(new_n656), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n429), .A2(new_n430), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n393), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n474), .B(KEYINPUT20), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n667), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n588), .A3(new_n578), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n653), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT34), .B(G104), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n674), .B(KEYINPUT104), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n673), .B(new_n675), .ZN(G6));
  NOR2_X1   g490(.A1(new_n431), .A2(new_n476), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n578), .A2(new_n588), .A3(new_n463), .A4(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n653), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT35), .B(G107), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G9));
  NAND2_X1  g495(.A1(new_n649), .A2(new_n650), .ZN(new_n682));
  INV_X1    g496(.A(new_n648), .ZN(new_n683));
  INV_X1    g497(.A(new_n370), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT36), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n684), .A2(new_n356), .A3(new_n685), .A4(new_n361), .ZN(new_n686));
  OAI22_X1  g500(.A1(new_n371), .A2(new_n374), .B1(new_n370), .B2(KEYINPUT36), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n686), .A2(new_n387), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n382), .B2(new_n385), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n682), .A2(new_n683), .A3(new_n652), .A4(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n645), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT37), .B(G110), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G12));
  AOI21_X1  g508(.A(new_n689), .B1(new_n304), .B2(new_n318), .ZN(new_n695));
  AOI211_X1 g509(.A(new_n568), .B(new_n544), .C1(new_n574), .C2(new_n575), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n567), .B1(new_n576), .B2(new_n545), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n478), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n638), .B1(new_n636), .B2(new_n637), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n628), .A2(new_n637), .A3(new_n638), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n591), .B(new_n309), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n592), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n643), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n590), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n698), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n695), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n427), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n423), .B2(new_n424), .ZN(new_n709));
  AOI21_X1  g523(.A(G902), .B1(new_n709), .B2(new_n428), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n463), .B(new_n670), .C1(new_n710), .C2(new_n394), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT105), .B(G900), .Z(new_n712));
  NAND2_X1  g526(.A1(new_n585), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n581), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n707), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n235), .ZN(G30));
  XNOR2_X1  g533(.A(new_n714), .B(KEYINPUT39), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n644), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT106), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT40), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n463), .B1(new_n431), .B2(new_n476), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n725), .A2(new_n479), .A3(new_n690), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n569), .A2(new_n577), .ZN(new_n727));
  XOR2_X1   g541(.A(new_n727), .B(KEYINPUT38), .Z(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n278), .A2(new_n280), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n268), .A2(new_n312), .ZN(new_n731));
  AOI21_X1  g545(.A(G902), .B1(new_n731), .B2(new_n280), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(G472), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n304), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n724), .A2(new_n726), .A3(new_n729), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G143), .ZN(G45));
  NAND2_X1  g551(.A1(new_n655), .A2(new_n656), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n665), .A2(new_n666), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n740), .B(new_n714), .C1(new_n431), .C2(new_n476), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n707), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n213), .ZN(G48));
  AOI21_X1  g557(.A(new_n390), .B1(new_n304), .B2(new_n318), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n588), .B(new_n478), .C1(new_n696), .C2(new_n697), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n699), .A2(new_n700), .ZN(new_n747));
  OAI21_X1  g561(.A(G469), .B1(new_n747), .B2(new_n308), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(KEYINPUT107), .A3(new_n701), .ZN(new_n749));
  OR3_X1    g563(.A1(new_n630), .A2(KEYINPUT107), .A3(new_n591), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n590), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n744), .A2(new_n746), .A3(new_n751), .A4(new_n671), .ZN(new_n752));
  XNOR2_X1  g566(.A(KEYINPUT41), .B(G113), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(G15));
  NOR2_X1   g568(.A1(new_n745), .A2(new_n711), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n744), .A3(new_n751), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G116), .ZN(G18));
  NOR4_X1   g571(.A1(new_n431), .A2(new_n476), .A3(new_n463), .A4(new_n587), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n695), .A2(new_n751), .A3(new_n758), .A4(new_n578), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G119), .ZN(G21));
  NOR2_X1   g574(.A1(new_n698), .A2(new_n725), .ZN(new_n761));
  INV_X1    g575(.A(G472), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n762), .B1(new_n301), .B2(new_n309), .ZN(new_n763));
  XOR2_X1   g577(.A(new_n294), .B(KEYINPUT108), .Z(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n315), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n311), .A2(new_n313), .A3(KEYINPUT109), .A4(new_n314), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n280), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n279), .A2(new_n267), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n765), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n763), .A2(new_n771), .A3(new_n390), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n761), .A2(new_n751), .A3(new_n588), .A4(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G122), .ZN(G24));
  INV_X1    g588(.A(new_n741), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n763), .A2(new_n771), .A3(new_n689), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n751), .A2(new_n775), .A3(new_n776), .A4(new_n578), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G125), .ZN(G27));
  INV_X1    g592(.A(KEYINPUT42), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n569), .A2(new_n478), .A3(new_n577), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n705), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n744), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n779), .B1(new_n782), .B2(new_n741), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n744), .A2(new_n781), .A3(KEYINPUT42), .A4(new_n775), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XOR2_X1   g599(.A(KEYINPUT110), .B(G131), .Z(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(G33));
  NOR2_X1   g601(.A1(new_n782), .A2(new_n717), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(new_n197), .ZN(G36));
  INV_X1    g603(.A(new_n701), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n634), .B1(new_n640), .B2(new_n642), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n591), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n794));
  OAI22_X1  g608(.A1(new_n793), .A2(new_n794), .B1(new_n792), .B2(new_n791), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n702), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT46), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n790), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(KEYINPUT46), .B(new_n702), .C1(new_n795), .C2(new_n796), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n590), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n677), .A2(new_n740), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT43), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n651), .A2(new_n652), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT43), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n677), .A2(new_n805), .A3(new_n740), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n803), .A2(new_n804), .A3(new_n690), .A4(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT44), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n780), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n803), .A2(new_n806), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(KEYINPUT44), .A3(new_n804), .A4(new_n690), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n801), .A2(new_n809), .A3(new_n811), .A4(new_n720), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G137), .ZN(G39));
  INV_X1    g627(.A(new_n780), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n390), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n815), .A2(new_n319), .A3(new_n741), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n799), .A2(new_n800), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n704), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT47), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n801), .A2(KEYINPUT47), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n817), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(new_n322), .ZN(G42));
  NAND4_X1  g638(.A1(new_n728), .A2(new_n478), .A3(new_n704), .A4(new_n391), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n749), .A2(new_n750), .ZN(new_n826));
  XOR2_X1   g640(.A(new_n826), .B(KEYINPUT49), .Z(new_n827));
  OR4_X1    g641(.A1(new_n735), .A2(new_n825), .A3(new_n802), .A4(new_n827), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n735), .A2(new_n581), .A3(new_n390), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n751), .A3(new_n814), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n677), .A2(new_n667), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n751), .A2(new_n814), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n810), .A2(new_n582), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n810), .A2(KEYINPUT116), .A3(new_n582), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n833), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n832), .B1(new_n838), .B2(new_n776), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n772), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n841), .B1(new_n836), .B2(new_n837), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n728), .A2(new_n479), .A3(new_n751), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT50), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n844), .A2(KEYINPUT117), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n842), .B(new_n843), .C1(new_n847), .C2(KEYINPUT50), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n840), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n826), .A2(new_n590), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n821), .A2(new_n822), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(new_n814), .A3(new_n842), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n849), .A2(KEYINPUT51), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n842), .A2(new_n578), .A3(new_n751), .ZN(new_n854));
  INV_X1    g668(.A(new_n671), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n854), .B(new_n579), .C1(new_n855), .C2(new_n830), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n838), .A2(new_n744), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n857), .A2(KEYINPUT48), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(KEYINPUT48), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n853), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n788), .B1(new_n783), .B2(new_n784), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n752), .A2(new_n759), .A3(new_n773), .A4(new_n756), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n645), .A2(new_n392), .B1(new_n653), .B2(new_n672), .ZN(new_n864));
  OAI22_X1  g678(.A1(new_n653), .A2(new_n678), .B1(new_n645), .B2(new_n691), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT112), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n775), .A2(new_n776), .A3(new_n867), .ZN(new_n868));
  NOR4_X1   g682(.A1(new_n431), .A2(new_n476), .A3(new_n463), .A4(new_n715), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n319), .A2(new_n690), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n781), .A2(new_n775), .A3(new_n776), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n871), .A2(new_n781), .B1(KEYINPUT112), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n862), .A2(new_n863), .A3(new_n866), .A4(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n695), .B(new_n706), .C1(new_n716), .C2(new_n775), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n714), .B(KEYINPUT113), .ZN(new_n876));
  AOI211_X1 g690(.A(new_n688), .B(new_n876), .C1(new_n382), .C2(new_n385), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n703), .A2(new_n877), .A3(new_n704), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT114), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT114), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n703), .A2(new_n877), .A3(new_n880), .A4(new_n704), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n761), .A2(new_n879), .A3(new_n735), .A4(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n875), .A2(new_n882), .A3(new_n777), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT115), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n875), .A2(new_n882), .A3(KEYINPUT115), .A4(new_n777), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT52), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n874), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n885), .A2(KEYINPUT52), .A3(new_n886), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n888), .A2(KEYINPUT53), .A3(new_n889), .ZN(new_n890));
  AND4_X1   g704(.A1(new_n862), .A2(new_n863), .A3(new_n866), .A4(new_n873), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n885), .A2(new_n886), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT52), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n883), .A2(KEYINPUT52), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n891), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n890), .B1(new_n896), .B2(KEYINPUT53), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT54), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n891), .A2(new_n894), .A3(new_n889), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT53), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT54), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n888), .A2(KEYINPUT53), .A3(new_n895), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n898), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT51), .B1(new_n849), .B2(new_n852), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n861), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(G952), .A2(G953), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n828), .B1(new_n907), .B2(new_n908), .ZN(G75));
  NOR2_X1   g723(.A1(new_n257), .A2(G952), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n570), .B(new_n558), .ZN(new_n911));
  XNOR2_X1  g725(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n901), .A2(new_n903), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n914), .A2(new_n308), .A3(new_n568), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT56), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT53), .B1(new_n888), .B2(new_n889), .ZN(new_n918));
  AND4_X1   g732(.A1(KEYINPUT53), .A2(new_n891), .A3(new_n895), .A4(new_n894), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n308), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(KEYINPUT119), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT119), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n914), .A2(new_n922), .A3(new_n308), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n921), .A2(new_n568), .A3(new_n923), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n913), .A2(new_n916), .ZN(new_n925));
  AOI211_X1 g739(.A(new_n910), .B(new_n917), .C1(new_n924), .C2(new_n925), .ZN(G51));
  XNOR2_X1  g740(.A(new_n592), .B(KEYINPUT57), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n902), .B1(new_n901), .B2(new_n903), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n904), .B1(new_n928), .B2(KEYINPUT120), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT120), .ZN(new_n930));
  AOI211_X1 g744(.A(new_n930), .B(new_n902), .C1(new_n901), .C2(new_n903), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n927), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n747), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n795), .A2(new_n796), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n921), .A2(new_n935), .A3(new_n923), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n910), .B1(new_n934), .B2(new_n936), .ZN(G54));
  AND2_X1   g751(.A1(KEYINPUT58), .A2(G475), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n921), .A2(new_n923), .A3(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n472), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n910), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n921), .A2(new_n472), .A3(new_n923), .A4(new_n938), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(G60));
  NAND2_X1  g758(.A1(G478), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT59), .Z(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n898), .B2(new_n904), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n942), .B1(new_n947), .B2(new_n665), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n929), .A2(new_n931), .ZN(new_n949));
  INV_X1    g763(.A(new_n665), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n950), .A2(new_n946), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n948), .B1(new_n949), .B2(new_n951), .ZN(G63));
  XNOR2_X1  g766(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n380), .A2(new_n430), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n914), .A2(new_n686), .A3(new_n687), .A4(new_n955), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n914), .A2(new_n955), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n367), .A2(new_n375), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n942), .B(new_n956), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT61), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(G66));
  NAND2_X1  g775(.A1(new_n863), .A2(new_n866), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n257), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT122), .Z(new_n964));
  INV_X1    g778(.A(G224), .ZN(new_n965));
  OAI21_X1  g779(.A(G953), .B1(new_n586), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n570), .B1(G898), .B2(new_n257), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(G69));
  AOI21_X1  g783(.A(new_n257), .B1(G227), .B2(G900), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT126), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n761), .A2(new_n744), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n801), .A2(new_n720), .A3(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n875), .A2(new_n777), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n812), .A2(new_n973), .A3(new_n974), .A4(new_n862), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n823), .A2(new_n975), .A3(new_n583), .ZN(new_n976));
  INV_X1    g790(.A(G900), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n257), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n971), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n978), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n812), .A2(new_n974), .A3(new_n862), .ZN(new_n981));
  INV_X1    g795(.A(new_n822), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n801), .A2(KEYINPUT47), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n816), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n981), .A2(new_n984), .A3(new_n973), .ZN(new_n985));
  OAI211_X1 g799(.A(KEYINPUT126), .B(new_n980), .C1(new_n985), .C2(new_n583), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n277), .B(KEYINPUT123), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(new_n466), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n979), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n812), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n722), .A2(new_n392), .A3(new_n780), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n855), .A2(new_n711), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT124), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n990), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n736), .A2(KEYINPUT62), .A3(new_n974), .ZN(new_n995));
  AOI21_X1  g809(.A(KEYINPUT62), .B1(new_n736), .B2(new_n974), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n984), .B(new_n994), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n988), .A2(new_n583), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n989), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n970), .B1(new_n1000), .B2(KEYINPUT125), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT125), .ZN(new_n1002));
  INV_X1    g816(.A(new_n970), .ZN(new_n1003));
  AOI211_X1 g817(.A(new_n1002), .B(new_n1003), .C1(new_n989), .C2(new_n999), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1001), .A2(new_n1004), .ZN(G72));
  INV_X1    g819(.A(new_n730), .ZN(new_n1006));
  NAND2_X1  g820(.A1(G472), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT63), .Z(new_n1008));
  NAND4_X1  g822(.A1(new_n897), .A2(new_n305), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1009), .B(KEYINPUT127), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1008), .B1(new_n997), .B2(new_n962), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n730), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1008), .B1(new_n985), .B2(new_n962), .ZN(new_n1013));
  INV_X1    g827(.A(new_n305), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n910), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n1010), .A2(new_n1016), .ZN(G57));
endmodule


