//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1206, new_n1207;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT65), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G137), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  OR2_X1    g043(.A1(new_n460), .A2(new_n461), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(G160));
  NOR2_X1   g048(.A1(new_n462), .A2(new_n465), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n478), .B1(G136), .B2(new_n463), .ZN(G162));
  INV_X1    g054(.A(G138), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(KEYINPUT67), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n481), .B(new_n483), .C1(new_n460), .C2(new_n461), .ZN(new_n484));
  OR2_X1    g059(.A1(G102), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n469), .A2(new_n481), .ZN(new_n488));
  XNOR2_X1  g063(.A(KEYINPUT67), .B(KEYINPUT4), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n460), .C2(new_n461), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n491), .B(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  XNOR2_X1  g070(.A(KEYINPUT5), .B(G543), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n496), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n497));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n496), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n499), .A2(new_n504), .ZN(G166));
  AND2_X1   g080(.A1(G63), .A2(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n496), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n496), .A2(new_n508), .A3(G89), .ZN(new_n509));
  NAND3_X1  g084(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n510));
  XNOR2_X1  g085(.A(new_n510), .B(KEYINPUT7), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n509), .A2(new_n511), .A3(KEYINPUT70), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g088(.A(KEYINPUT70), .B1(new_n509), .B2(new_n511), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n507), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G51), .ZN(new_n516));
  OAI21_X1  g091(.A(KEYINPUT68), .B1(new_n501), .B2(new_n502), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(new_n498), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT68), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n517), .A2(new_n522), .A3(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT69), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n517), .A2(new_n522), .A3(new_n525), .A4(G543), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n516), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n515), .A2(new_n527), .ZN(G168));
  NAND2_X1  g103(.A1(G77), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(new_n496), .ZN(new_n530));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n530), .A2(new_n503), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n532), .A2(G651), .B1(new_n533), .B2(G90), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n536), .B1(new_n524), .B2(new_n526), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n535), .A2(new_n537), .ZN(G171));
  AOI22_X1  g113(.A1(new_n496), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n498), .ZN(new_n540));
  INV_X1    g115(.A(G543), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n541), .B1(new_n508), .B2(KEYINPUT68), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n525), .B1(new_n542), .B2(new_n522), .ZN(new_n543));
  INV_X1    g118(.A(new_n526), .ZN(new_n544));
  OAI21_X1  g119(.A(G43), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n533), .A2(G81), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n545), .A2(KEYINPUT71), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT71), .ZN(new_n548));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n549), .B1(new_n524), .B2(new_n526), .ZN(new_n550));
  INV_X1    g125(.A(new_n546), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n540), .B1(new_n547), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n530), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n533), .A2(G91), .ZN(new_n563));
  AND2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n542), .A2(G53), .A3(new_n522), .ZN(new_n565));
  AND2_X1   g140(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  XNOR2_X1  g143(.A(KEYINPUT72), .B(KEYINPUT9), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(KEYINPUT73), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n570), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT73), .ZN(new_n573));
  NOR3_X1   g148(.A1(new_n572), .A2(new_n567), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n564), .B1(new_n571), .B2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G171), .ZN(G301));
  INV_X1    g151(.A(G168), .ZN(G286));
  INV_X1    g152(.A(G166), .ZN(G303));
  NAND2_X1  g153(.A1(new_n533), .A2(G87), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n542), .A2(G49), .A3(new_n522), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n496), .B2(G74), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G288));
  AOI22_X1  g157(.A1(new_n496), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n503), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n496), .A2(G61), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n498), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT74), .ZN(new_n589));
  AND2_X1   g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n588), .A2(new_n589), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n585), .B1(new_n590), .B2(new_n591), .ZN(G305));
  OAI21_X1  g167(.A(G47), .B1(new_n543), .B2(new_n544), .ZN(new_n593));
  NAND2_X1  g168(.A1(G72), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G60), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n530), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g171(.A(KEYINPUT75), .B(G85), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n596), .A2(G651), .B1(new_n533), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n593), .A2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  AND3_X1   g175(.A1(new_n496), .A2(new_n508), .A3(G92), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT76), .ZN(new_n602));
  XOR2_X1   g177(.A(new_n602), .B(KEYINPUT10), .Z(new_n603));
  INV_X1    g178(.A(G54), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n604), .B1(new_n524), .B2(new_n526), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT77), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n496), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(new_n498), .ZN(new_n608));
  OR3_X1    g183(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n606), .B1(new_n605), .B2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n603), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n600), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n600), .B1(new_n613), .B2(G868), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  INV_X1    g191(.A(new_n564), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n573), .B1(new_n572), .B2(new_n567), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n568), .A2(KEYINPUT73), .A3(new_n570), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n616), .B1(new_n620), .B2(G868), .ZN(G297));
  XOR2_X1   g196(.A(G297), .B(KEYINPUT78), .Z(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n613), .B1(new_n623), .B2(G860), .ZN(G148));
  NOR2_X1   g199(.A1(new_n553), .A2(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n613), .A2(new_n623), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT79), .Z(G323));
  XOR2_X1   g203(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n629));
  XNOR2_X1  g204(.A(G323), .B(new_n629), .ZN(G282));
  NAND2_X1  g205(.A1(new_n469), .A2(new_n466), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  INV_X1    g208(.A(G2100), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n463), .A2(G135), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n474), .A2(G123), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n465), .A2(G111), .ZN(new_n639));
  OAI21_X1  g214(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n637), .B(new_n638), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(G2096), .Z(new_n642));
  NAND3_X1  g217(.A1(new_n635), .A2(new_n636), .A3(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(KEYINPUT14), .A3(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT81), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n651), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT82), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n651), .A2(new_n653), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n651), .A2(new_n653), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(new_n655), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n657), .A2(new_n660), .A3(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT84), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g241(.A1(new_n657), .A2(KEYINPUT84), .A3(new_n660), .A4(new_n663), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT83), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n657), .A2(new_n663), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n669), .B1(new_n670), .B2(new_n659), .ZN(new_n671));
  AOI211_X1 g246(.A(KEYINPUT83), .B(new_n660), .C1(new_n657), .C2(new_n663), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n668), .B(G14), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT85), .ZN(G401));
  XNOR2_X1  g249(.A(G2084), .B(G2090), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2072), .B(G2078), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(KEYINPUT17), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n678), .B1(new_n679), .B2(new_n676), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT87), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n676), .A2(new_n677), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n682), .A2(new_n675), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n679), .A2(new_n676), .A3(new_n675), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n681), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G2096), .B(G2100), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G227));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT89), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n693), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(G1956), .B(G2474), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT90), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1961), .B(G1966), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT91), .B(KEYINPUT20), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NAND4_X1  g278(.A1(new_n697), .A2(new_n699), .A3(new_n701), .A4(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n699), .A2(new_n701), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n702), .B1(new_n696), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n699), .A2(new_n701), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n696), .A2(new_n708), .A3(new_n705), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n697), .A2(new_n707), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n704), .A2(new_n706), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT92), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(G1991), .B(G1996), .Z(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n711), .A2(KEYINPUT92), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n711), .A2(KEYINPUT92), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n718), .A2(new_n719), .A3(new_n713), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n715), .A2(new_n717), .A3(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n717), .B1(new_n715), .B2(new_n720), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n691), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n720), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n713), .B1(new_n718), .B2(new_n719), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n716), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n727), .A2(new_n690), .A3(new_n721), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(G229));
  MUX2_X1   g305(.A(G6), .B(G305), .S(G16), .Z(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT32), .B(G1981), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G16), .ZN(new_n734));
  NOR2_X1   g309(.A1(G166), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n734), .B2(G22), .ZN(new_n736));
  INV_X1    g311(.A(G1971), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G288), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(new_n734), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n734), .B2(G23), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT33), .B(G1976), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT95), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n736), .A2(new_n737), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n738), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n741), .A2(new_n743), .ZN(new_n747));
  NOR3_X1   g322(.A1(new_n733), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(KEYINPUT34), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(KEYINPUT34), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n463), .A2(G131), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n474), .A2(G119), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n465), .A2(G107), .ZN(new_n754));
  OAI21_X1  g329(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n752), .B(new_n753), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT94), .Z(new_n757));
  XOR2_X1   g332(.A(KEYINPUT93), .B(G29), .Z(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G25), .B2(new_n759), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT35), .B(G1991), .Z(new_n762));
  AND2_X1   g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  MUX2_X1   g339(.A(G24), .B(G290), .S(G16), .Z(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1986), .ZN(new_n766));
  NOR4_X1   g341(.A1(new_n763), .A2(new_n764), .A3(new_n766), .A4(KEYINPUT96), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n750), .A2(new_n751), .A3(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(KEYINPUT36), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n734), .A2(G20), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT23), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n620), .B2(new_n734), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT107), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G1956), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n769), .A2(KEYINPUT36), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n770), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(G32), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n778), .A2(G29), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n466), .A2(G105), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n463), .A2(G141), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n474), .A2(G129), .ZN(new_n782));
  NAND3_X1  g357(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT26), .Z(new_n784));
  AND4_X1   g359(.A1(new_n780), .A2(new_n781), .A3(new_n782), .A4(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n779), .B1(new_n786), .B2(G29), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT27), .B(G1996), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT101), .B(KEYINPUT24), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n789), .A2(G34), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n789), .A2(G34), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n790), .A2(new_n759), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G160), .B2(G29), .ZN(new_n793));
  OAI22_X1  g368(.A1(new_n787), .A2(new_n788), .B1(G2084), .B2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(G1961), .ZN(new_n795));
  NOR2_X1   g370(.A1(G5), .A2(G16), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT103), .Z(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G301), .B2(new_n734), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n794), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT105), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n734), .A2(G19), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n553), .B2(new_n734), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(G1341), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n734), .A2(G4), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n613), .B2(new_n734), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n800), .B(new_n803), .C1(G1348), .C2(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n798), .A2(new_n795), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT31), .B(G11), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT102), .ZN(new_n809));
  INV_X1    g384(.A(G28), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(KEYINPUT30), .ZN(new_n811));
  AOI21_X1  g386(.A(G29), .B1(new_n810), .B2(KEYINPUT30), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n809), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(G168), .A2(new_n734), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n734), .B2(G21), .ZN(new_n815));
  INV_X1    g390(.A(G1966), .ZN(new_n816));
  OAI221_X1 g391(.A(new_n813), .B1(new_n641), .B2(new_n758), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  AOI211_X1 g392(.A(new_n807), .B(new_n817), .C1(new_n816), .C2(new_n815), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT104), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n818), .A2(new_n819), .B1(G1348), .B2(new_n805), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n759), .A2(G35), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G162), .B2(new_n759), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT29), .Z(new_n823));
  INV_X1    g398(.A(G2090), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT106), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT25), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n463), .A2(G139), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n465), .B2(new_n832), .ZN(new_n833));
  MUX2_X1   g408(.A(G33), .B(new_n833), .S(G29), .Z(new_n834));
  AOI22_X1  g409(.A1(new_n787), .A2(new_n788), .B1(new_n834), .B2(G2072), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n793), .A2(G2084), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n835), .B(new_n836), .C1(G2072), .C2(new_n834), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n758), .A2(G26), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT99), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT28), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n463), .A2(G140), .ZN(new_n841));
  NOR2_X1   g416(.A1(G104), .A2(G2105), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT98), .Z(new_n843));
  OAI21_X1  g418(.A(G2104), .B1(new_n465), .B2(G116), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n474), .A2(KEYINPUT97), .A3(G128), .ZN(new_n845));
  AOI21_X1  g420(.A(KEYINPUT97), .B1(new_n474), .B2(G128), .ZN(new_n846));
  OAI221_X1 g421(.A(new_n841), .B1(new_n843), .B2(new_n844), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n840), .B1(G29), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT100), .B(G2067), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n759), .A2(G27), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(G164), .B2(new_n759), .ZN(new_n852));
  INV_X1    g427(.A(G2078), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n823), .B2(new_n824), .ZN(new_n855));
  NOR4_X1   g430(.A1(new_n826), .A2(new_n837), .A3(new_n850), .A4(new_n855), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n820), .B(new_n856), .C1(new_n819), .C2(new_n818), .ZN(new_n857));
  NOR3_X1   g432(.A1(new_n777), .A2(new_n806), .A3(new_n857), .ZN(G311));
  INV_X1    g433(.A(G311), .ZN(G150));
  NOR2_X1   g434(.A1(new_n612), .A2(new_n623), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT38), .ZN(new_n861));
  INV_X1    g436(.A(new_n540), .ZN(new_n862));
  AOI21_X1  g437(.A(KEYINPUT71), .B1(new_n545), .B2(new_n546), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n550), .A2(new_n548), .A3(new_n551), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(G55), .B1(new_n543), .B2(new_n544), .ZN(new_n866));
  NAND2_X1  g441(.A1(G80), .A2(G543), .ZN(new_n867));
  INV_X1    g442(.A(G67), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n867), .B1(new_n530), .B2(new_n868), .ZN(new_n869));
  AOI22_X1  g444(.A1(new_n869), .A2(G651), .B1(new_n533), .B2(G93), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n865), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n871), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n553), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n861), .B(new_n875), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n876), .A2(KEYINPUT39), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(KEYINPUT39), .ZN(new_n878));
  NOR3_X1   g453(.A1(new_n877), .A2(new_n878), .A3(G860), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n871), .A2(G860), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT37), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n879), .A2(new_n881), .ZN(G145));
  INV_X1    g457(.A(G37), .ZN(new_n883));
  XOR2_X1   g458(.A(G160), .B(new_n641), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(G162), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n847), .A2(new_n494), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n847), .A2(new_n494), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n785), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n786), .A3(new_n888), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n833), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n632), .B(new_n756), .Z(new_n894));
  NAND2_X1  g469(.A1(new_n474), .A2(G130), .ZN(new_n895));
  XOR2_X1   g470(.A(new_n895), .B(KEYINPUT108), .Z(new_n896));
  NAND2_X1  g471(.A1(new_n463), .A2(G142), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n465), .A2(G118), .ZN(new_n898));
  OAI21_X1  g473(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n896), .B(new_n897), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n894), .B(new_n900), .Z(new_n901));
  INV_X1    g476(.A(new_n833), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n890), .A2(new_n902), .A3(new_n891), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n893), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n901), .B1(new_n893), .B2(new_n903), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n886), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(KEYINPUT109), .ZN(new_n908));
  INV_X1    g483(.A(new_n906), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(new_n909), .A3(new_n885), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n904), .A2(KEYINPUT109), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n883), .B(new_n907), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT40), .ZN(G395));
  AOI211_X1 g488(.A(new_n540), .B(new_n871), .C1(new_n552), .C2(new_n547), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n547), .A2(new_n552), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n873), .B1(new_n915), .B2(new_n862), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n626), .B(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n603), .A2(new_n620), .A3(new_n611), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n620), .B1(new_n603), .B2(new_n611), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n612), .A2(G299), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n603), .A2(new_n620), .A3(new_n611), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(KEYINPUT41), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n918), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n920), .A2(new_n921), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n927), .B1(new_n928), .B2(new_n918), .ZN(new_n929));
  XNOR2_X1  g504(.A(G288), .B(KEYINPUT110), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(G305), .ZN(new_n931));
  XNOR2_X1  g506(.A(G290), .B(G166), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n931), .B(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(KEYINPUT42), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n929), .B(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(G868), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(G868), .B2(new_n873), .ZN(G295));
  OAI21_X1  g512(.A(new_n936), .B1(G868), .B2(new_n873), .ZN(G331));
  INV_X1    g513(.A(new_n514), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n939), .A2(new_n512), .B1(new_n496), .B2(new_n506), .ZN(new_n940));
  INV_X1    g515(.A(new_n527), .ZN(new_n941));
  INV_X1    g516(.A(new_n537), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n940), .A2(new_n941), .A3(new_n942), .A4(new_n534), .ZN(new_n943));
  OAI22_X1  g518(.A1(new_n515), .A2(new_n527), .B1(new_n535), .B2(new_n537), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n872), .A2(new_n874), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT113), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n872), .A2(new_n874), .A3(new_n945), .A4(KEYINPUT113), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n943), .A2(new_n944), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(new_n914), .B2(new_n916), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n875), .A2(KEYINPUT112), .A3(new_n951), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n950), .A2(new_n928), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n952), .A2(new_n946), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n922), .A2(new_n957), .A3(new_n925), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n933), .A3(new_n958), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n957), .A2(new_n921), .A3(new_n920), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT113), .B1(new_n917), .B2(new_n945), .ZN(new_n961));
  INV_X1    g536(.A(new_n949), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n954), .B(new_n955), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n926), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n960), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n959), .B(new_n883), .C1(new_n965), .C2(new_n933), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n956), .A2(new_n958), .ZN(new_n968));
  OAI211_X1 g543(.A(KEYINPUT114), .B(new_n883), .C1(new_n968), .C2(new_n933), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT114), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n933), .B1(new_n956), .B2(new_n958), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n970), .B1(new_n971), .B2(G37), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n972), .A3(new_n959), .ZN(new_n973));
  OAI211_X1 g548(.A(KEYINPUT44), .B(new_n967), .C1(new_n973), .C2(KEYINPUT43), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT115), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n975), .B1(new_n966), .B2(KEYINPUT43), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n959), .A2(new_n883), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n978));
  INV_X1    g553(.A(new_n933), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n954), .A2(new_n955), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n926), .B1(new_n980), .B2(new_n950), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n979), .B1(new_n981), .B2(new_n960), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n977), .A2(KEYINPUT115), .A3(new_n978), .A4(new_n982), .ZN(new_n983));
  AOI22_X1  g558(.A1(KEYINPUT43), .A2(new_n973), .B1(new_n976), .B2(new_n983), .ZN(new_n984));
  XOR2_X1   g559(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n985));
  OAI21_X1  g560(.A(new_n974), .B1(new_n984), .B2(new_n985), .ZN(G397));
  INV_X1    g561(.A(G40), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n468), .A2(new_n472), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G1384), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n488), .A2(new_n489), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n484), .A2(new_n486), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n491), .B(KEYINPUT66), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n989), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n988), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  XOR2_X1   g571(.A(new_n847), .B(G2067), .Z(new_n997));
  XNOR2_X1  g572(.A(new_n997), .B(KEYINPUT116), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n785), .ZN(new_n999));
  INV_X1    g574(.A(new_n996), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1996), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1001), .B1(new_n1002), .B2(new_n998), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n996), .A2(G1996), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1003), .B1(new_n785), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(new_n762), .A3(new_n757), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n847), .A2(G2067), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n996), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1004), .A2(KEYINPUT46), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT125), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1001), .B(new_n1010), .C1(KEYINPUT46), .C2(new_n1004), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT47), .ZN(new_n1012));
  XOR2_X1   g587(.A(new_n756), .B(new_n762), .Z(new_n1013));
  NAND2_X1  g588(.A1(new_n1000), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1005), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(G290), .A2(G1986), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1000), .A2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g592(.A(new_n1017), .B(KEYINPUT48), .Z(new_n1018));
  OAI21_X1  g593(.A(new_n1012), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1008), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT124), .ZN(new_n1021));
  AND2_X1   g596(.A1(G290), .A2(G1986), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1000), .B1(new_n1022), .B2(new_n1016), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1005), .A2(new_n1023), .A3(new_n1014), .ZN(new_n1024));
  INV_X1    g599(.A(G8), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1384), .B1(new_n490), .B2(new_n493), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n994), .A2(KEYINPUT50), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1028), .A2(new_n1029), .A3(new_n988), .ZN(new_n1030));
  INV_X1    g605(.A(G2084), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n463), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n470), .A2(new_n471), .ZN(new_n1033));
  OAI211_X1 g608(.A(G40), .B(new_n1032), .C1(new_n1033), .C2(new_n465), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1034), .B1(new_n994), .B2(new_n995), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1026), .A2(KEYINPUT45), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1030), .A2(new_n1031), .B1(new_n1037), .B2(new_n816), .ZN(new_n1038));
  AOI211_X1 g613(.A(KEYINPUT51), .B(new_n1025), .C1(new_n1038), .C2(G168), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1025), .B1(new_n1038), .B2(G168), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1037), .A2(new_n816), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1034), .B1(new_n994), .B2(KEYINPUT50), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n1028), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1041), .B1(G2084), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G286), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1040), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1039), .B1(new_n1046), .B2(KEYINPUT51), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT122), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(G2078), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  OAI221_X1 g626(.A(new_n1048), .B1(new_n1037), .B2(new_n1051), .C1(new_n1030), .C2(G1961), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1037), .A2(new_n1051), .ZN(new_n1053));
  AOI21_X1  g628(.A(G1961), .B1(new_n1042), .B2(new_n1028), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT122), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1037), .A2(KEYINPUT117), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1035), .A2(new_n1058), .A3(new_n1036), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT53), .B1(new_n1060), .B2(new_n853), .ZN(new_n1061));
  OAI21_X1  g636(.A(G171), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1035), .A2(new_n1058), .A3(new_n1036), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1058), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n853), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n1049), .ZN(new_n1066));
  OAI22_X1  g641(.A1(new_n1030), .A2(G1961), .B1(new_n1037), .B2(new_n1051), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1066), .A2(G301), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1062), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1047), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n994), .B2(new_n1034), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1026), .A2(new_n988), .A3(KEYINPUT121), .ZN(new_n1075));
  XOR2_X1   g650(.A(KEYINPUT58), .B(G1341), .Z(new_n1076));
  NAND3_X1  g651(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1077), .B1(new_n1037), .B2(G1996), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1078), .A2(KEYINPUT59), .A3(new_n553), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT59), .B1(new_n1078), .B2(new_n553), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT60), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n603), .A2(new_n1081), .A3(new_n611), .ZN(new_n1082));
  AOI21_X1  g657(.A(G2067), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1083));
  AOI21_X1  g658(.A(G1348), .B1(new_n1042), .B2(new_n1028), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  NOR3_X1   g660(.A1(new_n1079), .A2(new_n1080), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT61), .ZN(new_n1087));
  NAND2_X1  g662(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1088));
  INV_X1    g663(.A(G1956), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1043), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1091), .B(new_n564), .C1(new_n572), .C2(new_n567), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT56), .B(G2072), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1035), .A2(new_n1036), .A3(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1088), .A2(new_n1090), .A3(new_n1092), .A4(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1088), .A2(new_n1092), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1087), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n613), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1083), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1084), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n612), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT60), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1106), .A2(KEYINPUT61), .A3(new_n1095), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1086), .A2(new_n1098), .A3(new_n1103), .A4(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1097), .B1(new_n1102), .B2(new_n1095), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1056), .A2(new_n1061), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1071), .B1(new_n1111), .B2(G301), .ZN(new_n1112));
  AOI211_X1 g687(.A(KEYINPUT123), .B(new_n1067), .C1(new_n1065), .C2(new_n1049), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT123), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1115));
  OAI21_X1  g690(.A(G171), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT55), .ZN(new_n1119));
  XOR2_X1   g694(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n1120));
  NOR2_X1   g695(.A1(G166), .A2(new_n1025), .ZN(new_n1121));
  MUX2_X1   g696(.A(new_n1119), .B(new_n1120), .S(new_n1121), .Z(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1124), .A2(new_n737), .B1(new_n824), .B2(new_n1030), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1123), .B1(new_n1125), .B2(new_n1025), .ZN(new_n1126));
  INV_X1    g701(.A(G1981), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1127), .B(new_n585), .C1(new_n590), .C2(new_n591), .ZN(new_n1128));
  OAI21_X1  g703(.A(G1981), .B1(new_n584), .B2(new_n588), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT49), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1026), .A2(new_n988), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(G8), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1136), .A2(KEYINPUT119), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1136), .A2(KEYINPUT119), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1135), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT52), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n739), .B2(G1976), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n739), .A2(G1976), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1133), .A2(G8), .A3(new_n1142), .ZN(new_n1143));
  MUX2_X1   g718(.A(new_n1141), .B(new_n1140), .S(new_n1143), .Z(new_n1144));
  NAND2_X1  g719(.A1(new_n1139), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1057), .A2(new_n737), .A3(new_n1059), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1030), .A2(new_n824), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1025), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n1122), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1126), .A2(new_n1146), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1072), .A2(new_n1110), .A3(new_n1117), .A4(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(G8), .B1(new_n1044), .B2(G286), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1038), .A2(G168), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT51), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1039), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1157), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1151), .A2(new_n1062), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(G288), .A2(G1976), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1139), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1128), .ZN(new_n1166));
  OAI211_X1 g741(.A(G8), .B(new_n1133), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1146), .A2(new_n1149), .A3(new_n1122), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1038), .A2(new_n1025), .A3(G286), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1126), .A2(new_n1146), .A3(new_n1150), .A4(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT63), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1145), .B1(new_n1149), .B2(new_n1122), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1174), .A2(new_n1126), .A3(KEYINPUT63), .A4(new_n1170), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1169), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1153), .B(new_n1163), .C1(new_n1176), .C2(KEYINPUT120), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1169), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT120), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1021), .B(new_n1024), .C1(new_n1177), .C2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1176), .A2(KEYINPUT120), .ZN(new_n1186));
  AOI22_X1  g761(.A1(new_n1108), .A2(new_n1109), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1187));
  AOI21_X1  g762(.A(KEYINPUT54), .B1(new_n1062), .B2(new_n1069), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n1188), .A2(new_n1151), .A3(new_n1047), .ZN(new_n1189));
  AOI22_X1  g764(.A1(new_n1187), .A2(new_n1189), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1185), .A2(new_n1186), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1021), .B1(new_n1191), .B2(new_n1024), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1020), .B1(new_n1184), .B2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n1195));
  NAND2_X1  g769(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n1196));
  NAND2_X1  g770(.A1(new_n976), .A2(new_n983), .ZN(new_n1197));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g772(.A1(G227), .A2(new_n458), .ZN(new_n1199));
  XOR2_X1   g773(.A(new_n1199), .B(KEYINPUT126), .Z(new_n1200));
  NAND4_X1  g774(.A1(new_n729), .A2(new_n912), .A3(new_n673), .A4(new_n1200), .ZN(new_n1201));
  INV_X1    g775(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g776(.A(new_n1195), .B1(new_n1198), .B2(new_n1202), .ZN(new_n1203));
  AOI211_X1 g777(.A(KEYINPUT127), .B(new_n1201), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1204));
  NOR2_X1   g778(.A1(new_n1203), .A2(new_n1204), .ZN(G308));
  OAI21_X1  g779(.A(KEYINPUT127), .B1(new_n984), .B2(new_n1201), .ZN(new_n1206));
  NAND3_X1  g780(.A1(new_n1198), .A2(new_n1195), .A3(new_n1202), .ZN(new_n1207));
  NAND2_X1  g781(.A1(new_n1206), .A2(new_n1207), .ZN(G225));
endmodule


