//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G140), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  AND2_X1   g004(.A1(new_n190), .A2(G227), .ZN(new_n191));
  XOR2_X1   g005(.A(new_n189), .B(new_n191), .Z(new_n192));
  INV_X1    g006(.A(KEYINPUT67), .ZN(new_n193));
  XNOR2_X1  g007(.A(G143), .B(G146), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n193), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G143), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  AND4_X1   g015(.A1(new_n193), .A2(new_n196), .A3(new_n199), .A4(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n195), .B1(new_n199), .B2(KEYINPUT1), .ZN(new_n203));
  OAI22_X1  g017(.A1(new_n197), .A2(new_n202), .B1(new_n194), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT76), .ZN(new_n205));
  INV_X1    g019(.A(G101), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G104), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  AOI21_X1  g024(.A(KEYINPUT3), .B1(new_n210), .B2(G107), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(G107), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n206), .B(new_n209), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n208), .A2(G104), .ZN(new_n214));
  OAI21_X1  g028(.A(G101), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n204), .A2(new_n205), .A3(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT1), .B1(new_n200), .B2(G146), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n219), .A2(G128), .B1(new_n199), .B2(new_n201), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n196), .A2(new_n199), .A3(new_n201), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT67), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n194), .A2(new_n193), .A3(new_n196), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n220), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT76), .B1(new_n224), .B2(new_n216), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n218), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT10), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n200), .A2(KEYINPUT64), .A3(G146), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT64), .B1(new_n200), .B2(G146), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n199), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AND2_X1   g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n230), .A2(new_n233), .B1(new_n194), .B2(new_n231), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G101), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT4), .A3(new_n213), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT4), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n238), .A3(G101), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n226), .A2(new_n227), .B1(new_n234), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n219), .A2(G128), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n230), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n200), .A2(G146), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT64), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n246), .B1(new_n198), .B2(G143), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n200), .A2(KEYINPUT64), .A3(G146), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n245), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT68), .B1(new_n249), .B2(new_n203), .ZN(new_n250));
  AOI221_X4 g064(.A(KEYINPUT70), .B1(new_n223), .B2(new_n222), .C1(new_n244), .C2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n244), .A2(new_n250), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n222), .A2(new_n223), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI211_X1 g069(.A(KEYINPUT10), .B(new_n217), .C1(new_n251), .C2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT11), .ZN(new_n257));
  INV_X1    g071(.A(G134), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n257), .B1(new_n258), .B2(G137), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(G137), .ZN(new_n260));
  INV_X1    g074(.A(G137), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(KEYINPUT11), .A3(G134), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G131), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT65), .B(G131), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n265), .A2(new_n260), .A3(new_n259), .A4(new_n262), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n241), .A2(new_n256), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT77), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n205), .B1(new_n204), .B2(new_n217), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n224), .A2(KEYINPUT76), .A3(new_n216), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n227), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n240), .A2(new_n234), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n217), .A2(KEYINPUT10), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n242), .B1(new_n230), .B2(new_n243), .ZN(new_n278));
  NOR3_X1   g092(.A1(new_n249), .A2(KEYINPUT68), .A3(new_n203), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n254), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT70), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n244), .A2(new_n250), .B1(new_n223), .B2(new_n222), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n252), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n277), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n271), .B1(new_n276), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n241), .A2(new_n256), .A3(KEYINPUT77), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n267), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT78), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n270), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n285), .A2(KEYINPUT78), .A3(new_n267), .A4(new_n286), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n192), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OAI22_X1  g105(.A1(new_n272), .A2(new_n273), .B1(new_n280), .B2(new_n217), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n267), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT12), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT12), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n292), .A2(new_n295), .A3(new_n267), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n269), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n192), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n187), .B(new_n188), .C1(new_n291), .C2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(G469), .A2(G902), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n289), .A2(new_n192), .A3(new_n290), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n297), .A2(new_n298), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(G469), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n300), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G221), .ZN(new_n306));
  XOR2_X1   g120(.A(KEYINPUT9), .B(G234), .Z(new_n307));
  AOI21_X1  g121(.A(new_n306), .B1(new_n307), .B2(new_n188), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT22), .B(G137), .ZN(new_n311));
  INV_X1    g125(.A(G234), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n306), .A2(new_n312), .A3(G953), .ZN(new_n313));
  XOR2_X1   g127(.A(new_n311), .B(new_n313), .Z(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G119), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n316), .A2(G128), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(G128), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT24), .B(G110), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT16), .ZN(new_n323));
  INV_X1    g137(.A(G140), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n324), .A3(G125), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(G125), .ZN(new_n326));
  INV_X1    g140(.A(G125), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n325), .B1(new_n329), .B2(new_n323), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n198), .ZN(new_n331));
  OAI211_X1 g145(.A(G146), .B(new_n325), .C1(new_n329), .C2(new_n323), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n322), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT23), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT72), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n317), .B(new_n335), .C1(KEYINPUT71), .C2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT23), .B1(new_n195), .B2(G119), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT71), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT71), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n319), .A2(new_n341), .A3(KEYINPUT23), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n336), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n338), .B1(new_n343), .B2(new_n318), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n344), .A2(KEYINPUT73), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G110), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n347), .B1(new_n344), .B2(KEYINPUT73), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n334), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(G125), .B(G140), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT74), .B1(new_n350), .B2(new_n198), .ZN(new_n351));
  AND4_X1   g165(.A1(KEYINPUT74), .A2(new_n326), .A3(new_n328), .A4(new_n198), .ZN(new_n352));
  OR2_X1    g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n332), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n343), .A2(new_n318), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n337), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n347), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n320), .A2(new_n321), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n354), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n315), .B1(new_n349), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT73), .ZN(new_n361));
  OAI21_X1  g175(.A(G110), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n333), .B1(new_n362), .B2(new_n345), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n344), .A2(G110), .ZN(new_n364));
  INV_X1    g178(.A(new_n358), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n332), .B(new_n353), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n363), .A2(new_n366), .A3(new_n314), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n360), .A2(new_n367), .A3(new_n188), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT25), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n360), .A2(new_n367), .A3(KEYINPUT25), .A4(new_n188), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(KEYINPUT75), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G217), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n373), .B1(G234), .B2(new_n188), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT75), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n368), .A2(new_n375), .A3(new_n369), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n372), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n374), .A2(G902), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n360), .A2(new_n367), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n266), .ZN(new_n381));
  INV_X1    g195(.A(G131), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n261), .A2(G134), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n382), .B1(new_n260), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(new_n251), .B2(new_n255), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n234), .A2(new_n267), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n387), .B(KEYINPUT69), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(KEYINPUT30), .A3(new_n388), .ZN(new_n389));
  XOR2_X1   g203(.A(G116), .B(G119), .Z(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT2), .B(G113), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n390), .B(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT30), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n387), .A2(KEYINPUT66), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT66), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n234), .A2(new_n267), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n385), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n282), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n393), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n389), .A2(new_n392), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n392), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n386), .A2(new_n402), .A3(new_n388), .ZN(new_n403));
  NOR2_X1   g217(.A1(G237), .A2(G953), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G210), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(new_n206), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n407));
  XOR2_X1   g221(.A(new_n406), .B(new_n407), .Z(new_n408));
  NAND3_X1  g222(.A1(new_n401), .A2(new_n403), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT31), .ZN(new_n410));
  INV_X1    g224(.A(new_n408), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT28), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n392), .B1(new_n397), .B2(new_n399), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n412), .B1(new_n403), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n392), .B1(new_n267), .B2(new_n234), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT28), .B1(new_n386), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n411), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT31), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n401), .A2(new_n418), .A3(new_n403), .A4(new_n408), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n410), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(G472), .A2(G902), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n420), .A2(KEYINPUT32), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT32), .B1(new_n420), .B2(new_n421), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n398), .B1(new_n281), .B2(new_n283), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT69), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n387), .B(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n392), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n403), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n416), .B1(new_n429), .B2(KEYINPUT28), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n408), .A2(KEYINPUT29), .ZN(new_n431));
  AOI21_X1  g245(.A(G902), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n414), .A2(new_n416), .A3(new_n411), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n408), .B1(new_n401), .B2(new_n403), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT29), .ZN(new_n436));
  OAI21_X1  g250(.A(G472), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n380), .B1(new_n424), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G214), .B1(G237), .B2(G902), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n190), .A2(G224), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n234), .A2(new_n327), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n254), .B(new_n327), .C1(new_n278), .C2(new_n279), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n442), .B1(new_n443), .B2(KEYINPUT82), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(KEYINPUT82), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n441), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT82), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n448), .B1(new_n282), .B2(new_n327), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n445), .B(new_n440), .C1(new_n449), .C2(new_n442), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT81), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n237), .A2(new_n392), .A3(new_n239), .ZN(new_n454));
  OR2_X1    g268(.A1(new_n390), .A2(new_n391), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n456));
  INV_X1    g270(.A(G116), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(G119), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n459), .B(G113), .C1(new_n390), .C2(new_n456), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n217), .A2(new_n455), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n454), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(G110), .B(G122), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n453), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n454), .A2(new_n461), .A3(KEYINPUT81), .A4(new_n463), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT80), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n462), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n454), .A2(KEYINPUT80), .A3(new_n461), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n464), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT6), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n452), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT84), .ZN(new_n477));
  OR2_X1    g291(.A1(new_n477), .A2(KEYINPUT7), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(KEYINPUT7), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n440), .A3(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n480), .B1(new_n444), .B2(new_n446), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT85), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n444), .A2(new_n446), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(KEYINPUT7), .A3(new_n440), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n463), .B(KEYINPUT8), .Z(new_n486));
  INV_X1    g300(.A(KEYINPUT5), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n459), .B(G113), .C1(new_n487), .C2(new_n390), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n455), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n486), .B1(new_n489), .B2(new_n217), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT83), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n460), .A2(new_n455), .A3(new_n216), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n491), .B1(new_n490), .B2(new_n492), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT85), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n496), .B(new_n480), .C1(new_n444), .C2(new_n446), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n495), .A2(new_n467), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n188), .B1(new_n485), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G210), .B1(G237), .B2(G902), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(KEYINPUT86), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n476), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n501), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n495), .A2(new_n467), .A3(new_n497), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n444), .A2(new_n446), .A3(new_n441), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n505), .A2(KEYINPUT7), .B1(new_n481), .B2(KEYINPUT85), .ZN(new_n506));
  AOI21_X1  g320(.A(G902), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n475), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n474), .B1(new_n467), .B2(new_n471), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n451), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n503), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n439), .B1(new_n502), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(G475), .A2(G902), .ZN(new_n513));
  XNOR2_X1  g327(.A(G113), .B(G122), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(new_n210), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n404), .A2(G214), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n200), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n404), .A2(G143), .A3(G214), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n265), .A3(new_n518), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n519), .A2(KEYINPUT88), .ZN(new_n520));
  INV_X1    g334(.A(new_n265), .ZN(new_n521));
  INV_X1    g335(.A(new_n518), .ZN(new_n522));
  AOI21_X1  g336(.A(G143), .B1(new_n404), .B2(G214), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT88), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n517), .A2(new_n525), .A3(new_n265), .A4(new_n518), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT89), .B1(new_n520), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n519), .A2(KEYINPUT88), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT89), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n529), .A2(new_n530), .A3(new_n524), .A4(new_n526), .ZN(new_n531));
  INV_X1    g345(.A(new_n332), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n350), .B(KEYINPUT19), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n532), .B1(new_n198), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n528), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  OAI22_X1  g349(.A1(new_n351), .A2(new_n352), .B1(new_n198), .B2(new_n350), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT87), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT87), .ZN(new_n538));
  OAI221_X1 g352(.A(new_n538), .B1(new_n198), .B2(new_n350), .C1(new_n351), .C2(new_n352), .ZN(new_n539));
  NAND2_X1  g353(.A1(KEYINPUT18), .A2(G131), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n517), .A2(new_n518), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n540), .B1(new_n517), .B2(new_n518), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n537), .A2(new_n539), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n515), .B1(new_n535), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n521), .B(KEYINPUT17), .C1(new_n522), .C2(new_n523), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n331), .A2(new_n546), .A3(new_n332), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n529), .A2(new_n548), .A3(new_n524), .A4(new_n526), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n550), .A2(new_n544), .A3(new_n515), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n513), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT20), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT20), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n554), .B(new_n513), .C1(new_n545), .C2(new_n551), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n515), .B1(new_n550), .B2(new_n544), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n188), .B1(new_n551), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT90), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT90), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n560), .B(new_n188), .C1(new_n551), .C2(new_n557), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(G475), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  OR2_X1    g378(.A1(KEYINPUT93), .A2(G952), .ZN(new_n565));
  NAND2_X1  g379(.A1(KEYINPUT93), .A2(G952), .ZN(new_n566));
  AOI21_X1  g380(.A(G953), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G237), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n567), .B1(new_n312), .B2(new_n568), .ZN(new_n569));
  OAI211_X1 g383(.A(G902), .B(G953), .C1(new_n312), .C2(new_n568), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(KEYINPUT94), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT21), .B(G898), .Z(new_n572));
  OAI21_X1  g386(.A(new_n569), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G478), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n574), .A2(KEYINPUT15), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n200), .A2(G128), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n195), .A2(G143), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT91), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n578), .B1(new_n576), .B2(new_n577), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n258), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT13), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n582), .B1(new_n195), .B2(G143), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n577), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n576), .A2(new_n582), .ZN(new_n585));
  OAI21_X1  g399(.A(G134), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G122), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(G116), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n457), .A2(G122), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(G107), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n588), .A2(new_n589), .A3(new_n208), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n581), .A2(new_n586), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT92), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n581), .A2(new_n586), .A3(new_n593), .A4(KEYINPUT92), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n588), .A2(KEYINPUT14), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n590), .A2(new_n599), .A3(G107), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n588), .B(new_n589), .C1(KEYINPUT14), .C2(new_n208), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n580), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(G134), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n602), .B1(new_n605), .B2(new_n581), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n598), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n307), .A2(G217), .A3(new_n190), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n609), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n598), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n575), .B1(new_n613), .B2(new_n188), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n611), .B1(new_n598), .B2(new_n607), .ZN(new_n615));
  AOI211_X1 g429(.A(new_n609), .B(new_n606), .C1(new_n596), .C2(new_n597), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n188), .B(new_n575), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n564), .A2(new_n573), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT95), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n564), .A2(KEYINPUT95), .A3(new_n573), .A4(new_n619), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n512), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n310), .A2(new_n438), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(new_n206), .ZN(G3));
  INV_X1    g440(.A(KEYINPUT96), .ZN(new_n627));
  INV_X1    g441(.A(G472), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n420), .A2(new_n188), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n630), .B1(new_n420), .B2(new_n188), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n631), .A2(new_n632), .A3(new_n380), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n310), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n501), .B1(new_n476), .B2(new_n499), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n507), .A2(new_n503), .A3(new_n510), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n636), .A2(KEYINPUT97), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT97), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n507), .A2(new_n510), .A3(new_n639), .A4(new_n503), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n638), .A2(new_n439), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n610), .A2(KEYINPUT33), .A3(new_n612), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT99), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n615), .A2(new_n616), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n646), .A2(KEYINPUT99), .A3(KEYINPUT33), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT33), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n649), .B1(new_n615), .B2(new_n616), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT98), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT98), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n652), .B(new_n649), .C1(new_n615), .C2(new_n616), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n574), .A2(G902), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n648), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT100), .B(G478), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n658), .B1(new_n646), .B2(G902), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n661), .A2(KEYINPUT101), .A3(new_n564), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT101), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n663), .B1(new_n660), .B2(new_n563), .ZN(new_n664));
  INV_X1    g478(.A(new_n573), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n662), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n635), .A2(new_n642), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT34), .B(G104), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G6));
  NOR3_X1   g483(.A1(new_n563), .A2(new_n665), .A3(new_n619), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n635), .A2(new_n642), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(new_n208), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT102), .B(KEYINPUT35), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G9));
  NAND2_X1  g488(.A1(new_n363), .A2(new_n366), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n315), .A2(KEYINPUT36), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n378), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n370), .A2(KEYINPUT75), .A3(new_n371), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n376), .A2(new_n374), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n682), .A2(new_n631), .A3(new_n632), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n310), .A2(new_n624), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT103), .B(KEYINPUT37), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(new_n347), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n684), .B(new_n686), .ZN(G12));
  AOI21_X1  g501(.A(new_n641), .B1(new_n424), .B2(new_n437), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n563), .A2(new_n619), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n569), .B1(new_n571), .B2(G900), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n310), .A2(new_n681), .A3(new_n688), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G128), .ZN(G30));
  XOR2_X1   g507(.A(new_n690), .B(KEYINPUT39), .Z(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n310), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT40), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n628), .A2(new_n188), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n628), .B1(new_n429), .B2(new_n411), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n698), .B1(new_n699), .B2(new_n409), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n700), .B(KEYINPUT104), .Z(new_n701));
  NAND2_X1  g515(.A1(new_n424), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT105), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n502), .A2(new_n511), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT38), .ZN(new_n705));
  INV_X1    g519(.A(new_n439), .ZN(new_n706));
  INV_X1    g520(.A(new_n619), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n563), .A2(new_n707), .ZN(new_n708));
  NOR4_X1   g522(.A1(new_n705), .A2(new_n706), .A3(new_n681), .A4(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n697), .A2(new_n703), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n696), .A2(KEYINPUT40), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(new_n200), .ZN(G45));
  NAND3_X1  g527(.A1(new_n660), .A2(new_n563), .A3(new_n690), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n310), .A2(new_n681), .A3(new_n688), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G146), .ZN(G48));
  NAND2_X1  g531(.A1(new_n420), .A2(new_n421), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT32), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n420), .A2(KEYINPUT32), .A3(new_n421), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n437), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n666), .A2(new_n722), .A3(new_n642), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n287), .A2(new_n288), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n290), .A3(new_n269), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n299), .B1(new_n725), .B2(new_n298), .ZN(new_n726));
  OAI21_X1  g540(.A(G469), .B1(new_n726), .B2(G902), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n309), .A3(new_n300), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n380), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n723), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g546(.A(KEYINPUT41), .B(G113), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G15));
  NAND2_X1  g548(.A1(new_n688), .A2(new_n670), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n731), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n457), .ZN(G18));
  INV_X1    g551(.A(new_n722), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n738), .A2(new_n641), .A3(new_n682), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n622), .A2(new_n623), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n729), .A3(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n739), .A2(new_n729), .A3(KEYINPUT106), .A4(new_n740), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G119), .ZN(G21));
  OAI211_X1 g560(.A(new_n410), .B(new_n419), .C1(new_n408), .C2(new_n430), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n421), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n628), .B1(new_n420), .B2(new_n188), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n748), .B1(new_n749), .B2(KEYINPUT107), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n751));
  AOI211_X1 g565(.A(new_n751), .B(new_n628), .C1(new_n420), .C2(new_n188), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n750), .A2(new_n380), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n641), .A2(new_n708), .ZN(new_n754));
  AND4_X1   g568(.A1(new_n573), .A2(new_n753), .A3(new_n729), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n587), .ZN(G24));
  NOR4_X1   g570(.A1(new_n750), .A2(new_n752), .A3(new_n682), .A4(new_n714), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n728), .A2(new_n641), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XOR2_X1   g573(.A(KEYINPUT108), .B(G125), .Z(new_n760));
  XNOR2_X1  g574(.A(new_n759), .B(new_n760), .ZN(G27));
  INV_X1    g575(.A(new_n437), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n762), .B1(new_n763), .B2(new_n720), .ZN(new_n764));
  OAI21_X1  g578(.A(KEYINPUT110), .B1(new_n422), .B2(new_n423), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n380), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n297), .A2(new_n767), .A3(new_n298), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n767), .B1(new_n297), .B2(new_n298), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n302), .A3(G469), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n300), .A2(new_n301), .A3(new_n771), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n636), .A2(new_n439), .A3(new_n637), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n772), .A2(new_n309), .A3(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n766), .A2(KEYINPUT42), .A3(new_n715), .A4(new_n774), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n774), .A2(new_n438), .A3(new_n715), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n775), .B1(KEYINPUT42), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G131), .ZN(G33));
  NAND3_X1  g592(.A1(new_n774), .A2(new_n438), .A3(new_n691), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G134), .ZN(G36));
  NAND3_X1  g594(.A1(new_n770), .A2(new_n302), .A3(KEYINPUT45), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(G469), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT45), .B1(new_n302), .B2(new_n303), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n301), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n300), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT46), .B1(new_n784), .B2(new_n301), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n309), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n788), .A2(new_n694), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n636), .A2(new_n439), .A3(new_n637), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n661), .A2(new_n563), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT43), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT43), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n793), .B1(new_n661), .B2(new_n563), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n631), .A2(new_n632), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n792), .A2(KEYINPUT111), .A3(new_n794), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n797), .A2(new_n799), .A3(new_n681), .A4(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT44), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n790), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(new_n802), .B2(new_n801), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n789), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(new_n261), .ZN(G39));
  XNOR2_X1  g620(.A(new_n788), .B(KEYINPUT47), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n738), .A2(new_n715), .A3(new_n380), .A4(new_n773), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT112), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(new_n324), .ZN(G42));
  NOR2_X1   g625(.A1(new_n308), .A2(new_n706), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n705), .A2(new_n730), .A3(new_n791), .A4(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n727), .A2(new_n300), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n813), .B1(KEYINPUT49), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n703), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n816), .B(new_n817), .C1(KEYINPUT49), .C2(new_n815), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n662), .A2(new_n664), .ZN(new_n819));
  NOR4_X1   g633(.A1(new_n728), .A2(new_n380), .A3(new_n569), .A4(new_n790), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n821), .A2(new_n567), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n569), .B1(new_n792), .B2(new_n794), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n823), .A2(new_n753), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n642), .A3(new_n729), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n822), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n822), .A2(KEYINPUT117), .A3(new_n827), .A4(new_n828), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n728), .A2(new_n790), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n766), .A2(new_n823), .A3(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT48), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n831), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT118), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n824), .A2(new_n773), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n814), .A2(new_n308), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n839), .B1(new_n807), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n824), .A2(new_n706), .A3(new_n705), .A4(new_n729), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n842), .A2(KEYINPUT50), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n750), .A2(new_n752), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n833), .A2(new_n823), .A3(new_n681), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n842), .A2(KEYINPUT50), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n817), .A2(new_n564), .A3(new_n661), .A4(new_n820), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n843), .A2(new_n845), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n838), .B1(new_n841), .B2(new_n848), .ZN(new_n849));
  OR3_X1    g663(.A1(new_n841), .A2(new_n838), .A3(new_n848), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n837), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n757), .A2(new_n774), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n619), .A2(new_n556), .A3(new_n562), .A4(new_n690), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n377), .B2(new_n678), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n773), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n424), .B2(new_n437), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT114), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n310), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n854), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n681), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n790), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n305), .A2(new_n862), .A3(new_n722), .A4(new_n309), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT114), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n779), .A2(new_n853), .A3(new_n859), .A4(new_n864), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n310), .B(new_n624), .C1(new_n438), .C2(new_n683), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n706), .B1(new_n636), .B2(new_n637), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n310), .A2(new_n633), .A3(new_n867), .A4(new_n670), .ZN(new_n868));
  AOI221_X4 g682(.A(new_n665), .B1(new_n556), .B2(new_n562), .C1(new_n656), .C2(new_n659), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT113), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n869), .A2(new_n870), .A3(new_n867), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n870), .B1(new_n869), .B2(new_n867), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(new_n310), .A3(new_n633), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n866), .A2(new_n868), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n865), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n739), .B(new_n310), .C1(new_n691), .C2(new_n715), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT52), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n772), .A2(new_n309), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n682), .A2(new_n690), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n880), .A2(new_n641), .A3(new_n708), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n879), .A2(new_n881), .A3(new_n702), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n877), .A2(new_n878), .A3(new_n759), .A4(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n692), .A2(new_n716), .A3(new_n759), .A4(new_n882), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT52), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n876), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n731), .B1(new_n723), .B2(new_n735), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(new_n755), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n745), .A2(new_n888), .A3(new_n777), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n886), .A2(KEYINPUT53), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT53), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n876), .A2(new_n885), .A3(new_n883), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n745), .A2(new_n888), .A3(new_n777), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n852), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT115), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n886), .B(new_n889), .C1(new_n896), .C2(new_n891), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n876), .A2(new_n885), .A3(new_n883), .A4(new_n896), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n898), .B(KEYINPUT53), .C1(new_n892), .C2(new_n893), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT54), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n836), .A2(KEYINPUT118), .ZN(new_n901));
  NOR4_X1   g715(.A1(new_n851), .A2(new_n895), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(G952), .A2(G953), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT119), .Z(new_n904));
  OAI21_X1  g718(.A(new_n818), .B1(new_n902), .B2(new_n904), .ZN(G75));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n190), .A2(G952), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n897), .A2(G902), .A3(new_n899), .A4(new_n501), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT56), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n508), .A2(new_n509), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(new_n451), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT55), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT120), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n915), .B1(new_n909), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n908), .B1(new_n911), .B2(new_n917), .ZN(new_n918));
  AND4_X1   g732(.A1(KEYINPUT120), .A2(new_n909), .A3(new_n910), .A4(new_n914), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n906), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n909), .A2(new_n910), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n909), .A2(new_n916), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n921), .B1(new_n922), .B2(new_n915), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n911), .A2(new_n917), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n923), .A2(KEYINPUT121), .A3(new_n924), .A4(new_n908), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n920), .A2(new_n925), .ZN(G51));
  NAND2_X1  g740(.A1(new_n897), .A2(new_n899), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n927), .A2(new_n188), .A3(new_n784), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT122), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n301), .B(KEYINPUT57), .Z(new_n931));
  NOR2_X1   g745(.A1(new_n927), .A2(new_n852), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n931), .B1(new_n932), .B2(new_n900), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(new_n291), .B2(new_n299), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n907), .B1(new_n930), .B2(new_n934), .ZN(G54));
  INV_X1    g749(.A(new_n927), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n936), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n545), .A2(new_n551), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(new_n907), .ZN(G60));
  NAND2_X1  g755(.A1(new_n648), .A2(new_n654), .ZN(new_n942));
  NAND2_X1  g756(.A1(G478), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT59), .Z(new_n944));
  NOR2_X1   g758(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n932), .B2(new_n900), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n908), .ZN(new_n947));
  INV_X1    g761(.A(new_n944), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n948), .B1(new_n900), .B2(new_n895), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n942), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n949), .A2(KEYINPUT123), .A3(new_n942), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n947), .B1(new_n952), .B2(new_n953), .ZN(G63));
  NAND2_X1  g768(.A1(G217), .A2(G902), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT60), .Z(new_n956));
  NAND2_X1  g770(.A1(new_n936), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n360), .A2(new_n367), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n936), .A2(new_n677), .A3(new_n956), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n959), .A2(new_n908), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT61), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n959), .A2(KEYINPUT61), .A3(new_n908), .A4(new_n960), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(G66));
  AOI21_X1  g779(.A(new_n190), .B1(new_n572), .B2(G224), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n745), .A2(new_n888), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n967), .A2(new_n875), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n966), .B1(new_n969), .B2(new_n190), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n912), .B1(G898), .B2(new_n190), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n970), .B(new_n971), .Z(G69));
  AOI21_X1  g786(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n389), .A2(new_n400), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n533), .B(KEYINPUT124), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT125), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n877), .A2(new_n759), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n712), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT62), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n980), .A2(new_n810), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n661), .A2(new_n564), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n438), .B(new_n773), .C1(new_n982), .C2(new_n689), .ZN(new_n983));
  OAI22_X1  g797(.A1(new_n789), .A2(new_n804), .B1(new_n696), .B2(new_n983), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT126), .Z(new_n985));
  NAND2_X1  g799(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n977), .B1(new_n986), .B2(new_n190), .ZN(new_n987));
  INV_X1    g801(.A(new_n976), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n988), .B1(G900), .B2(G953), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n777), .B(new_n779), .C1(new_n807), .C2(new_n809), .ZN(new_n991));
  INV_X1    g805(.A(new_n789), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n992), .A2(new_n754), .A3(new_n766), .ZN(new_n993));
  NOR4_X1   g807(.A1(new_n991), .A2(new_n993), .A3(new_n805), .A4(new_n978), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n990), .B1(new_n994), .B2(new_n190), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n973), .B1(new_n987), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n190), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n989), .ZN(new_n998));
  INV_X1    g812(.A(new_n973), .ZN(new_n999));
  AOI21_X1  g813(.A(G953), .B1(new_n981), .B2(new_n985), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n998), .B(new_n999), .C1(new_n1000), .C2(new_n977), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n996), .A2(new_n1001), .ZN(G72));
  XNOR2_X1  g816(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(new_n698), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1005), .B1(new_n994), .B2(new_n968), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n401), .A2(new_n403), .A3(new_n411), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n908), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n401), .A2(new_n403), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n408), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n981), .A2(new_n985), .A3(new_n968), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1010), .B1(new_n1011), .B2(new_n1004), .ZN(new_n1012));
  INV_X1    g826(.A(new_n409), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1004), .B1(new_n1013), .B2(new_n435), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1014), .B1(new_n890), .B2(new_n894), .ZN(new_n1015));
  NOR3_X1   g829(.A1(new_n1008), .A2(new_n1012), .A3(new_n1015), .ZN(G57));
endmodule


