//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  AND2_X1   g017(.A1(G2072), .A2(G2078), .ZN(new_n443));
  NAND3_X1  g018(.A1(new_n443), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT66), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n466), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT67), .B1(new_n468), .B2(new_n463), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n462), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n464), .A2(new_n466), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n462), .ZN(new_n477));
  INV_X1    g052(.A(G137), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n472), .A2(new_n479), .ZN(G160));
  INV_X1    g055(.A(new_n477), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n476), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  AOI22_X1  g058(.A1(G136), .A2(new_n481), .B1(new_n483), .B2(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT68), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n484), .A2(new_n487), .ZN(G162));
  NAND3_X1  g063(.A1(new_n467), .A2(new_n469), .A3(G138), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(KEYINPUT4), .B(G138), .C1(new_n468), .C2(new_n463), .ZN(new_n492));
  NAND2_X1  g067(.A1(G102), .A2(G2104), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(new_n462), .ZN(new_n495));
  OAI21_X1  g070(.A(G126), .B1(new_n468), .B2(new_n463), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n490), .B1(G114), .B2(G2104), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n462), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n491), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  NAND2_X1  g076(.A1(G75), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G62), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n502), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT5), .B(G543), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(new_n508), .A3(G62), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g087(.A(G651), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT71), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n505), .A2(new_n506), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT69), .B(G88), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  OAI21_X1  g095(.A(G543), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n517), .A2(new_n518), .B1(new_n522), .B2(G50), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n513), .A2(new_n514), .A3(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n514), .B1(new_n513), .B2(new_n523), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT72), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n521), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g106(.A(KEYINPUT72), .B(G543), .C1(new_n519), .C2(new_n520), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(KEYINPUT5), .A2(G543), .ZN(new_n534));
  OAI211_X1 g109(.A(G63), .B(G651), .C1(new_n534), .C2(new_n504), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT7), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n538), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n504), .A2(new_n534), .B1(new_n519), .B2(new_n520), .ZN(new_n541));
  INV_X1    g116(.A(G89), .ZN(new_n542));
  OAI211_X1 g117(.A(new_n535), .B(new_n540), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n533), .A2(new_n543), .ZN(G168));
  NAND2_X1  g119(.A1(new_n531), .A2(new_n532), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G52), .ZN(new_n546));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n534), .A2(new_n504), .ZN(new_n548));
  INV_X1    g123(.A(G64), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n550), .A2(G651), .B1(new_n517), .B2(G90), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n546), .A2(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G56), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n548), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G651), .ZN(new_n557));
  XNOR2_X1  g132(.A(KEYINPUT73), .B(G81), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n517), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(G43), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n531), .B2(new_n532), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  OAI211_X1 g143(.A(G53), .B(G543), .C1(new_n519), .C2(new_n520), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n570));
  XNOR2_X1  g145(.A(KEYINPUT6), .B(G651), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n571), .A2(new_n572), .A3(G53), .A4(G543), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n510), .A2(new_n571), .A3(G91), .ZN(new_n575));
  INV_X1    g150(.A(G651), .ZN(new_n576));
  AND2_X1   g151(.A1(G78), .A2(G543), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(new_n510), .B2(G65), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n574), .B(new_n575), .C1(new_n576), .C2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G168), .ZN(G286));
  NAND2_X1  g155(.A1(new_n517), .A2(G87), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n522), .A2(G49), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(G288));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  OR3_X1    g160(.A1(new_n541), .A2(KEYINPUT74), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(KEYINPUT74), .B1(new_n541), .B2(new_n585), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n548), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(new_n522), .B2(G48), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n588), .A2(new_n592), .ZN(G305));
  XNOR2_X1  g168(.A(KEYINPUT76), .B(G47), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n545), .A2(new_n594), .B1(G85), .B2(new_n517), .ZN(new_n595));
  INV_X1    g170(.A(G60), .ZN(new_n596));
  INV_X1    g171(.A(G72), .ZN(new_n597));
  INV_X1    g172(.A(G543), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n548), .A2(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(KEYINPUT75), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n601));
  OAI221_X1 g176(.A(new_n601), .B1(new_n597), .B2(new_n598), .C1(new_n548), .C2(new_n596), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n600), .A2(G651), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n595), .A2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n541), .B2(new_n607), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n510), .A2(new_n571), .A3(KEYINPUT10), .A4(G92), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g185(.A(KEYINPUT72), .B1(new_n571), .B2(G543), .ZN(new_n611));
  INV_X1    g186(.A(new_n532), .ZN(new_n612));
  OAI21_X1  g187(.A(G54), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G66), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n548), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G651), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n610), .A2(new_n613), .A3(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n605), .B1(new_n619), .B2(G868), .ZN(G284));
  OAI21_X1  g195(.A(new_n605), .B1(new_n619), .B2(G868), .ZN(G321));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(G299), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n622), .B2(G168), .ZN(G297));
  OAI21_X1  g199(.A(new_n623), .B1(new_n622), .B2(G168), .ZN(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n619), .B1(new_n626), .B2(G860), .ZN(G148));
  NOR2_X1   g202(.A1(new_n563), .A2(G868), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n618), .A2(G559), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n628), .B1(new_n630), .B2(G868), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT77), .Z(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND3_X1   g208(.A1(new_n467), .A2(new_n469), .A3(new_n474), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT12), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT78), .B(KEYINPUT13), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2100), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n481), .A2(G135), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n483), .A2(G123), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n462), .A2(G111), .ZN(new_n644));
  OAI21_X1  g219(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n642), .B(new_n643), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT79), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT80), .B(G2096), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n641), .A2(new_n649), .ZN(G156));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(new_n655), .A3(KEYINPUT14), .ZN(new_n656));
  XOR2_X1   g231(.A(G1341), .B(G1348), .Z(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2451), .B(G2454), .Z(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(new_n663), .ZN(new_n665));
  AND3_X1   g240(.A1(new_n664), .A2(G14), .A3(new_n665), .ZN(G401));
  XOR2_X1   g241(.A(G2067), .B(G2678), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT82), .ZN(new_n668));
  NOR2_X1   g243(.A1(G2072), .A2(G2078), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n443), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n668), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT18), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n668), .A2(new_n670), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n670), .B(KEYINPUT17), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n675), .B(new_n672), .C1(new_n668), .C2(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n668), .A2(new_n671), .A3(new_n676), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n674), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2096), .B(G2100), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT83), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1956), .B(G2474), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n687), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n686), .A2(new_n687), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n691), .A2(KEYINPUT20), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(KEYINPUT20), .ZN(new_n693));
  OAI221_X1 g268(.A(new_n688), .B1(new_n685), .B2(new_n689), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G1991), .B(G1996), .Z(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1981), .B(G1986), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n696), .A2(new_n698), .ZN(new_n701));
  AND3_X1   g276(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n700), .B1(new_n699), .B2(new_n701), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(G229));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G22), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G166), .B2(new_n705), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n707), .A2(G1971), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(G1971), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n705), .A2(G6), .ZN(new_n710));
  INV_X1    g285(.A(G305), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(new_n705), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT32), .B(G1981), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n705), .A2(G23), .ZN(new_n715));
  INV_X1    g290(.A(G288), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n705), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT33), .B(G1976), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT85), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n717), .B(new_n719), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n708), .A2(new_n709), .A3(new_n714), .A4(new_n720), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G25), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n481), .A2(G131), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n483), .A2(G119), .ZN(new_n727));
  OR2_X1    g302(.A1(G95), .A2(G2105), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n728), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n725), .B1(new_n731), .B2(new_n724), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT35), .B(G1991), .Z(new_n733));
  XOR2_X1   g308(.A(new_n732), .B(new_n733), .Z(new_n734));
  AND2_X1   g309(.A1(new_n705), .A2(G24), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G290), .B2(G16), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(G1986), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n737), .A2(G1986), .ZN(new_n739));
  NOR3_X1   g314(.A1(new_n734), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n722), .A2(new_n723), .A3(new_n740), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT36), .Z(new_n742));
  AOI22_X1  g317(.A1(new_n481), .A2(G141), .B1(G105), .B2(new_n474), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n483), .A2(G129), .ZN(new_n744));
  NAND3_X1  g319(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT26), .Z(new_n746));
  NAND3_X1  g321(.A1(new_n743), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  MUX2_X1   g322(.A(G32), .B(new_n747), .S(G29), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT89), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT27), .B(G1996), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n749), .B(new_n750), .Z(new_n751));
  INV_X1    g326(.A(KEYINPUT24), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n724), .B1(new_n752), .B2(G34), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n752), .B2(G34), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G160), .B2(G29), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G2084), .ZN(new_n756));
  NOR2_X1   g331(.A1(G29), .A2(G33), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n757), .A2(KEYINPUT88), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n757), .A2(KEYINPUT88), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n467), .A2(new_n469), .A3(G127), .ZN(new_n760));
  NAND2_X1  g335(.A1(G115), .A2(G2104), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n462), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT25), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G139), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n765), .B1(new_n477), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n758), .B(new_n759), .C1(new_n768), .C2(G29), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n756), .B1(new_n769), .B2(G2072), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(G2072), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n755), .A2(G2084), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT90), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G16), .B2(G21), .ZN(new_n774));
  NAND2_X1  g349(.A1(G168), .A2(G16), .ZN(new_n775));
  MUX2_X1   g350(.A(new_n773), .B(new_n774), .S(new_n775), .Z(new_n776));
  INV_X1    g351(.A(G1966), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n772), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n724), .A2(G35), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G162), .B2(new_n724), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT29), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n771), .B(new_n778), .C1(new_n781), .C2(G2090), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n751), .A2(new_n770), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n781), .A2(G2090), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n705), .A2(G20), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT23), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n570), .A2(new_n573), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n575), .B1(new_n578), .B2(new_n576), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n786), .B1(new_n789), .B2(new_n705), .ZN(new_n790));
  INV_X1    g365(.A(G1956), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n784), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT96), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n705), .A2(G5), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G171), .B2(new_n705), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT92), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G1961), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT93), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT31), .B(G11), .Z(new_n801));
  INV_X1    g376(.A(G28), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n802), .A2(KEYINPUT30), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT91), .Z(new_n804));
  AOI21_X1  g379(.A(G29), .B1(new_n802), .B2(KEYINPUT30), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n801), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n647), .B2(new_n724), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n724), .A2(G26), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT28), .Z(new_n809));
  OR2_X1    g384(.A1(G104), .A2(G2105), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n810), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n811));
  INV_X1    g386(.A(G140), .ZN(new_n812));
  INV_X1    g387(.A(G128), .ZN(new_n813));
  OAI221_X1 g388(.A(new_n811), .B1(new_n477), .B2(new_n812), .C1(new_n813), .C2(new_n482), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n809), .B1(new_n814), .B2(G29), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT87), .B(G2067), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n807), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n777), .B2(new_n776), .ZN(new_n819));
  NOR2_X1   g394(.A1(G4), .A2(G16), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT86), .Z(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n618), .B2(new_n705), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1348), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n798), .B2(G1961), .ZN(new_n824));
  NAND2_X1  g399(.A1(G164), .A2(G29), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G27), .B2(G29), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT94), .B(G2078), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT95), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n563), .A2(G16), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(G16), .B2(G19), .ZN(new_n830));
  INV_X1    g405(.A(G1341), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n826), .A2(new_n828), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n832), .B(new_n833), .C1(new_n828), .C2(new_n826), .ZN(new_n834));
  NOR3_X1   g409(.A1(new_n819), .A2(new_n824), .A3(new_n834), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n783), .A2(new_n794), .A3(new_n800), .A4(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n742), .A2(new_n836), .ZN(G311));
  OR2_X1    g412(.A1(new_n742), .A2(new_n836), .ZN(G150));
  NAND2_X1  g413(.A1(new_n545), .A2(G55), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n517), .A2(G93), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n839), .B(new_n840), .C1(new_n576), .C2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G860), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT37), .Z(new_n844));
  AOI22_X1  g419(.A1(new_n556), .A2(G651), .B1(new_n517), .B2(new_n558), .ZN(new_n845));
  OAI21_X1  g420(.A(G43), .B1(new_n611), .B2(new_n612), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n845), .A2(new_n846), .A3(KEYINPUT97), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(KEYINPUT98), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT98), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n845), .A2(new_n846), .A3(KEYINPUT97), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT97), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n560), .B2(new_n562), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(new_n842), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n848), .A2(new_n853), .A3(new_n842), .A4(new_n850), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n626), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT38), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n857), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n862));
  INV_X1    g437(.A(G860), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n861), .B2(KEYINPUT39), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n844), .B1(new_n862), .B2(new_n864), .ZN(G145));
  XNOR2_X1  g440(.A(new_n747), .B(new_n768), .ZN(new_n866));
  INV_X1    g441(.A(new_n638), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n481), .A2(G142), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n483), .A2(G130), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n462), .A2(G118), .ZN(new_n870));
  OAI21_X1  g445(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n868), .B(new_n869), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n867), .A2(new_n872), .ZN(new_n874));
  OR3_X1    g449(.A1(new_n866), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n866), .B1(new_n873), .B2(new_n874), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n500), .B(new_n814), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n730), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n875), .A2(new_n879), .A3(new_n876), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n647), .B(G160), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(G162), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(G37), .B1(new_n883), .B2(new_n885), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g464(.A1(new_n857), .A2(new_n629), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n630), .B1(new_n855), .B2(new_n856), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT99), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(new_n618), .B2(new_n789), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n608), .A2(new_n609), .B1(G651), .B2(new_n616), .ZN(new_n896));
  NAND4_X1  g471(.A1(G299), .A2(new_n896), .A3(KEYINPUT99), .A4(new_n613), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n618), .A2(new_n789), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n893), .A2(KEYINPUT100), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(KEYINPUT100), .B1(new_n893), .B2(new_n900), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT41), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n903), .B1(new_n618), .B2(new_n789), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n898), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT101), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n900), .A2(new_n903), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT101), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n898), .A2(new_n908), .A3(new_n904), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n902), .B1(new_n892), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n510), .A2(G62), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n913), .A2(KEYINPUT70), .B1(G75), .B2(G543), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n576), .B1(new_n914), .B2(new_n511), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n517), .A2(new_n518), .ZN(new_n916));
  INV_X1    g491(.A(G50), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n916), .B1(new_n917), .B2(new_n521), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT71), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n919), .A2(new_n524), .A3(G305), .ZN(new_n920));
  AOI21_X1  g495(.A(G305), .B1(new_n919), .B2(new_n524), .ZN(new_n921));
  NAND2_X1  g496(.A1(G290), .A2(new_n716), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n595), .A2(new_n603), .A3(G288), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n920), .A2(new_n921), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n711), .B1(new_n525), .B2(new_n526), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n919), .A2(new_n524), .A3(G305), .ZN(new_n927));
  AOI22_X1  g502(.A1(new_n926), .A2(new_n927), .B1(new_n922), .B2(new_n923), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n912), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n924), .B1(new_n920), .B2(new_n921), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n926), .A2(new_n922), .A3(new_n923), .A4(new_n927), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT102), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT42), .ZN(new_n934));
  OR3_X1    g509(.A1(new_n925), .A2(new_n928), .A3(KEYINPUT42), .ZN(new_n935));
  AND4_X1   g510(.A1(new_n901), .A2(new_n911), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n911), .A2(new_n901), .B1(new_n934), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(G868), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n842), .A2(new_n622), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(G295));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n939), .ZN(G331));
  XOR2_X1   g516(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n898), .A2(new_n908), .A3(new_n904), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n908), .B1(new_n898), .B2(new_n904), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT41), .B1(new_n898), .B2(new_n899), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n545), .A2(G51), .ZN(new_n949));
  INV_X1    g524(.A(new_n543), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n533), .A2(new_n543), .A3(KEYINPUT104), .ZN(new_n952));
  OAI21_X1  g527(.A(G171), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(G168), .A2(new_n948), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT104), .B1(new_n533), .B2(new_n543), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(G301), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n857), .A2(new_n957), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n855), .A2(new_n856), .A3(new_n953), .A4(new_n956), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT105), .B1(new_n947), .B2(new_n960), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT102), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT102), .B1(new_n930), .B2(new_n931), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n856), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n848), .A2(new_n850), .B1(new_n853), .B2(new_n842), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n965), .A2(new_n957), .A3(new_n966), .ZN(new_n967));
  AOI22_X1  g542(.A1(new_n855), .A2(new_n856), .B1(new_n953), .B2(new_n956), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n969), .A2(new_n910), .A3(new_n970), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n895), .A2(new_n897), .B1(new_n789), .B2(new_n618), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n972), .B1(new_n958), .B2(new_n959), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n961), .A2(new_n964), .A3(new_n971), .A4(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G37), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n909), .B1(KEYINPUT41), .B2(new_n972), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n959), .B(new_n958), .C1(new_n978), .C2(new_n945), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n973), .B1(new_n979), .B2(KEYINPUT105), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n964), .B1(new_n980), .B2(new_n971), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n943), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n983));
  INV_X1    g558(.A(new_n975), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n905), .B1(new_n972), .B2(KEYINPUT41), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n958), .A2(new_n985), .A3(new_n959), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n933), .B1(new_n986), .B2(new_n973), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n987), .A2(new_n976), .A3(new_n942), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n983), .B1(new_n984), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n969), .A2(new_n985), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n974), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(G37), .B1(new_n991), .B2(new_n933), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n992), .A2(KEYINPUT106), .A3(new_n975), .A4(new_n942), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n982), .A2(new_n989), .A3(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n977), .A2(new_n981), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n992), .A2(new_n975), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n995), .A2(new_n942), .B1(KEYINPUT43), .B2(new_n996), .ZN(new_n997));
  MUX2_X1   g572(.A(new_n994), .B(new_n997), .S(KEYINPUT44), .Z(G397));
  INV_X1    g573(.A(G1384), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n500), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G40), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n472), .A2(new_n479), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G1996), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n747), .B(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G2067), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n814), .B(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n731), .A2(new_n733), .ZN(new_n1011));
  OR2_X1    g586(.A1(new_n731), .A2(new_n733), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(G290), .B(G1986), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1006), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT108), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1016), .B1(new_n1000), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n498), .B1(new_n462), .B2(new_n494), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1384), .B1(new_n1020), .B2(new_n491), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1021), .A2(KEYINPUT108), .A3(new_n1017), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1000), .A2(KEYINPUT50), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1019), .A2(new_n1022), .A3(new_n1004), .A4(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1348), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1021), .A2(new_n1004), .A3(new_n1009), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n619), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1004), .B1(new_n1021), .B2(KEYINPUT45), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT56), .B(G2072), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n500), .A2(new_n1034), .A3(new_n999), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1035), .B(new_n1004), .C1(new_n1021), .C2(new_n1017), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1032), .A2(new_n1033), .B1(new_n791), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(G299), .B(KEYINPUT57), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT118), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1036), .A2(new_n791), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1033), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1030), .A2(new_n1031), .A3(new_n1043), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1041), .B(new_n1038), .C1(new_n1042), .C2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1029), .A2(new_n1040), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1040), .A2(KEYINPUT61), .A3(new_n1045), .A4(new_n1047), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1026), .A2(KEYINPUT60), .A3(new_n618), .A4(new_n1027), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n1051));
  NOR2_X1   g626(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1042), .A2(new_n1044), .A3(new_n1038), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1049), .A2(new_n1050), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1030), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1021), .A2(KEYINPUT45), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1056), .A2(new_n1057), .A3(new_n1007), .A4(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1058), .A2(new_n1002), .A3(new_n1007), .A4(new_n1004), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT119), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1021), .A2(new_n1004), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(G1341), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1059), .A2(new_n1061), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n563), .A2(KEYINPUT121), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1067), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT60), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n619), .B1(new_n1028), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT60), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1074));
  OAI22_X1  g649(.A1(new_n1070), .A2(new_n1071), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1048), .B1(new_n1055), .B2(new_n1075), .ZN(new_n1076));
  NOR3_X1   g651(.A1(new_n1030), .A2(new_n1031), .A3(G2078), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT53), .ZN(new_n1078));
  XNOR2_X1  g653(.A(KEYINPUT123), .B(G1961), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1024), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1077), .A2(KEYINPUT53), .ZN(new_n1082));
  OAI21_X1  g657(.A(G171), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1077), .A2(KEYINPUT53), .B1(new_n1024), .B2(new_n1079), .ZN(new_n1084));
  OR2_X1    g659(.A1(new_n1077), .A2(KEYINPUT53), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1084), .A2(new_n1085), .A3(G301), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT54), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n777), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1088));
  NOR4_X1   g663(.A1(new_n472), .A2(new_n479), .A3(new_n1003), .A4(G2084), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1019), .A2(new_n1022), .A3(new_n1023), .A4(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n1090), .A3(G168), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G8), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT51), .ZN(new_n1093));
  AOI21_X1  g668(.A(G168), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT51), .ZN(new_n1095));
  OAI211_X1 g670(.A(G8), .B(new_n1091), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1032), .A2(G1971), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT109), .B(G2090), .Z(new_n1099));
  NOR2_X1   g674(.A1(new_n1036), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(G8), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT110), .ZN(new_n1102));
  NAND4_X1  g677(.A1(G303), .A2(new_n1102), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n919), .A2(G8), .A3(new_n524), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT55), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT110), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1101), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n716), .A2(G1976), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1062), .A2(G8), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT111), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1062), .A2(KEYINPUT111), .A3(G8), .A4(new_n1111), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(KEYINPUT52), .A3(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n592), .B1(new_n585), .B2(new_n541), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(G1981), .ZN(new_n1118));
  XOR2_X1   g693(.A(KEYINPUT112), .B(G1981), .Z(new_n1119));
  NAND3_X1  g694(.A1(new_n588), .A2(new_n592), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT113), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT49), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1062), .A2(G8), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT49), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1121), .A2(KEYINPUT113), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(G1976), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT52), .B1(G288), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1124), .A2(new_n1111), .A3(new_n1129), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1116), .A2(new_n1127), .A3(new_n1130), .ZN(new_n1131));
  OAI22_X1  g706(.A1(new_n1024), .A2(new_n1099), .B1(new_n1032), .B2(G1971), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1132), .A2(new_n1108), .A3(G8), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1110), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1087), .A2(new_n1097), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1086), .A2(KEYINPUT54), .ZN(new_n1136));
  AOI21_X1  g711(.A(G301), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT124), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1083), .A2(new_n1086), .A3(new_n1139), .A4(KEYINPUT54), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1076), .A2(new_n1135), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT63), .ZN(new_n1143));
  NAND2_X1  g718(.A1(G168), .A2(G8), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1144), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1145), .A2(KEYINPUT116), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT116), .ZN(new_n1147));
  AOI211_X1 g722(.A(new_n1147), .B(new_n1144), .C1(new_n1088), .C2(new_n1090), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1143), .B1(new_n1134), .B2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1133), .B(KEYINPUT63), .C1(new_n1146), .C2(new_n1148), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1108), .B1(new_n1132), .B2(G8), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1116), .A2(new_n1127), .A3(new_n1130), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT114), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT114), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1116), .A2(new_n1127), .A3(new_n1130), .A4(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1153), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT117), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1152), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AOI211_X1 g735(.A(KEYINPUT117), .B(new_n1153), .C1(new_n1155), .C2(new_n1157), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1150), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1133), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n716), .A2(new_n1128), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n1165), .B(KEYINPUT115), .Z(new_n1166));
  OAI21_X1  g741(.A(new_n1120), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1163), .B1(new_n1124), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1142), .A2(new_n1162), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1093), .A2(new_n1096), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1172), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1137), .A2(new_n1110), .A3(new_n1131), .A4(new_n1133), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(KEYINPUT62), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1170), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  AND4_X1   g753(.A1(new_n1133), .A2(new_n1137), .A3(new_n1131), .A4(new_n1110), .ZN(new_n1179));
  AND4_X1   g754(.A1(new_n1170), .A2(new_n1179), .A3(new_n1177), .A4(new_n1172), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1015), .B1(new_n1169), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1013), .A2(new_n1006), .ZN(new_n1183));
  NOR2_X1   g758(.A1(G290), .A2(G1986), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1006), .A2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1183), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1187), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n1002), .A2(new_n1005), .A3(G1996), .ZN(new_n1189));
  OR2_X1    g764(.A1(new_n1189), .A2(KEYINPUT46), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(KEYINPUT46), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1010), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1006), .B1(new_n1192), .B2(new_n747), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1190), .A2(new_n1191), .A3(new_n1193), .ZN(new_n1194));
  XOR2_X1   g769(.A(new_n1194), .B(KEYINPUT47), .Z(new_n1195));
  NAND2_X1  g770(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1196));
  OAI22_X1  g771(.A1(new_n1196), .A2(new_n1011), .B1(G2067), .B2(new_n814), .ZN(new_n1197));
  AOI211_X1 g772(.A(new_n1188), .B(new_n1195), .C1(new_n1006), .C2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1182), .A2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n1201));
  NOR3_X1   g775(.A1(G401), .A2(G227), .A3(new_n460), .ZN(new_n1202));
  OAI21_X1  g776(.A(new_n1202), .B1(new_n702), .B2(new_n703), .ZN(new_n1203));
  AOI21_X1  g777(.A(new_n1203), .B1(new_n886), .B2(new_n887), .ZN(new_n1204));
  AND3_X1   g778(.A1(new_n994), .A2(new_n1201), .A3(new_n1204), .ZN(new_n1205));
  AOI21_X1  g779(.A(new_n1201), .B1(new_n994), .B2(new_n1204), .ZN(new_n1206));
  NOR2_X1   g780(.A1(new_n1205), .A2(new_n1206), .ZN(G308));
  NAND2_X1  g781(.A1(new_n994), .A2(new_n1204), .ZN(G225));
endmodule


