//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1303,
    new_n1304, new_n1305, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  OAI21_X1  g0010(.A(G50), .B1(G58), .B2(G68), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT65), .Z(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT66), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n222), .A2(new_n223), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n207), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n210), .B(new_n216), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(KEYINPUT73), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  OAI211_X1 g0050(.A(G223), .B(new_n248), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  OAI211_X1 g0051(.A(G226), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G87), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G274), .ZN(new_n262));
  AND2_X1   g0062(.A1(G1), .A2(G13), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n262), .B1(new_n263), .B2(new_n257), .ZN(new_n264));
  INV_X1    g0064(.A(new_n260), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n261), .A2(G232), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AND3_X1   g0066(.A1(new_n256), .A2(G190), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G200), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n268), .B1(new_n256), .B2(new_n266), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n247), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n256), .A2(G190), .A3(new_n266), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n264), .A2(new_n265), .ZN(new_n272));
  INV_X1    g0072(.A(G232), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n258), .A2(new_n260), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(new_n255), .B2(new_n254), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n271), .B(KEYINPUT73), .C1(new_n276), .C2(new_n268), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n270), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT8), .B(G58), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT68), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT8), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G58), .ZN(new_n282));
  OR2_X1    g0082(.A1(new_n282), .A2(KEYINPUT68), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n213), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n288), .B1(new_n259), .B2(G20), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n286), .B1(new_n284), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n288), .ZN(new_n292));
  INV_X1    g0092(.A(G58), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(new_n218), .ZN(new_n294));
  OAI21_X1  g0094(.A(G20), .B1(new_n294), .B2(new_n201), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G159), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(KEYINPUT3), .A2(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(KEYINPUT3), .A2(G33), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(new_n214), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT7), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n249), .A2(new_n250), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n298), .B1(new_n306), .B2(G68), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n292), .B1(new_n307), .B2(KEYINPUT16), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT16), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n218), .B1(new_n303), .B2(new_n305), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n309), .B1(new_n310), .B2(new_n298), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n291), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n278), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT17), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT18), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT7), .B1(new_n304), .B2(new_n214), .ZN(new_n317));
  NOR4_X1   g0117(.A1(new_n249), .A2(new_n250), .A3(new_n302), .A4(G20), .ZN(new_n318));
  OAI21_X1  g0118(.A(G68), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n298), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(KEYINPUT16), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n311), .A2(new_n321), .A3(new_n288), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n290), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n276), .A2(G179), .ZN(new_n324));
  INV_X1    g0124(.A(G169), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n325), .B1(new_n256), .B2(new_n266), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n316), .B1(new_n323), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n323), .A2(new_n316), .A3(new_n328), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n278), .A2(KEYINPUT17), .A3(new_n312), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n315), .A2(new_n330), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n299), .A2(new_n300), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(G232), .A3(G1698), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(G226), .A3(new_n248), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G97), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n255), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT13), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n258), .A2(G274), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n342), .A2(new_n260), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(G238), .B2(new_n261), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n340), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n341), .B1(new_n340), .B2(new_n344), .ZN(new_n346));
  OAI21_X1  g0146(.A(G169), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT14), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n340), .A2(new_n344), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT13), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n340), .A2(new_n344), .A3(new_n341), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT14), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(new_n353), .A3(G169), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n350), .A2(G179), .A3(new_n351), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n348), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n296), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n357), .A2(new_n202), .B1(new_n214), .B2(G68), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n214), .A2(G33), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(new_n220), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n288), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT11), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n289), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT12), .ZN(new_n365));
  INV_X1    g0165(.A(new_n285), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n365), .B1(new_n366), .B2(new_n218), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n285), .A2(KEYINPUT12), .A3(G68), .ZN(new_n368));
  OAI22_X1  g0168(.A1(new_n364), .A2(new_n218), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n361), .A2(new_n362), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n363), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n356), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n352), .A2(G200), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n350), .A2(G190), .A3(new_n351), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(new_n371), .A3(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n272), .B1(new_n221), .B2(new_n274), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n335), .A2(G232), .A3(new_n248), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n335), .A2(G238), .A3(G1698), .ZN(new_n379));
  INV_X1    g0179(.A(G107), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n378), .B(new_n379), .C1(new_n380), .C2(new_n335), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n377), .B1(new_n381), .B2(new_n255), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n382), .A2(G169), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT71), .ZN(new_n385));
  INV_X1    g0185(.A(G179), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n382), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n385), .B1(new_n382), .B2(new_n386), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n384), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n366), .A2(new_n220), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n364), .B2(new_n220), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n214), .A2(new_n220), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT69), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n279), .B(new_n394), .ZN(new_n395));
  OAI211_X1 g0195(.A(KEYINPUT70), .B(new_n393), .C1(new_n395), .C2(new_n357), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT70), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n293), .A2(KEYINPUT8), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n282), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n394), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n279), .A2(KEYINPUT69), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n357), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n397), .B1(new_n402), .B2(new_n392), .ZN(new_n403));
  XOR2_X1   g0203(.A(KEYINPUT15), .B(G87), .Z(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n396), .B(new_n403), .C1(new_n405), .C2(new_n359), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n391), .B1(new_n406), .B2(new_n288), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n389), .A2(new_n407), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n382), .A2(G190), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n382), .A2(new_n268), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n408), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n334), .A2(new_n373), .A3(new_n376), .A4(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G226), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n272), .B1(new_n414), .B2(new_n274), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n335), .A2(G222), .A3(new_n248), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n335), .A2(G223), .A3(G1698), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n416), .B(new_n417), .C1(new_n220), .C2(new_n335), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT67), .ZN(new_n419));
  OR2_X1    g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n258), .B1(new_n418), .B2(new_n419), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n415), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT9), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n285), .A2(G50), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n289), .B2(G50), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n280), .A2(new_n214), .A3(new_n283), .A4(G33), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n296), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n423), .B(new_n425), .C1(new_n428), .C2(new_n292), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n292), .B1(new_n426), .B2(new_n427), .ZN(new_n430));
  INV_X1    g0230(.A(new_n425), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT9), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n422), .A2(G190), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n420), .A2(new_n421), .ZN(new_n434));
  OAI21_X1  g0234(.A(G200), .B1(new_n434), .B2(new_n415), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(KEYINPUT72), .A2(KEYINPUT10), .ZN(new_n437));
  OR2_X1    g0237(.A1(KEYINPUT72), .A2(KEYINPUT10), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n433), .A2(new_n435), .A3(KEYINPUT72), .A4(KEYINPUT10), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n422), .A2(new_n386), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n425), .B1(new_n428), .B2(new_n292), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n441), .B(new_n442), .C1(G169), .C2(new_n422), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n439), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n413), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G283), .ZN(new_n446));
  INV_X1    g0246(.A(G97), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n446), .B(new_n214), .C1(G33), .C2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G116), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G20), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n288), .A2(KEYINPUT79), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT79), .B1(new_n288), .B2(new_n450), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n448), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT20), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(KEYINPUT20), .B(new_n448), .C1(new_n451), .C2(new_n452), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(KEYINPUT80), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n259), .A2(G33), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n285), .A2(new_n458), .A3(new_n213), .A4(new_n287), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G116), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(G116), .B2(new_n366), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT80), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n453), .A2(new_n462), .A3(new_n454), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n457), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  OAI211_X1 g0264(.A(G264), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n465));
  OAI211_X1 g0265(.A(G257), .B(new_n248), .C1(new_n249), .C2(new_n250), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n299), .A2(G303), .A3(new_n300), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n255), .ZN(new_n469));
  INV_X1    g0269(.A(G41), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n259), .B(G45), .C1(new_n470), .C2(KEYINPUT5), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT5), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(G41), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n258), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G270), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT76), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n472), .B2(G41), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n470), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n479));
  INV_X1    g0279(.A(G45), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(G1), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n472), .A2(G41), .ZN(new_n482));
  AND4_X1   g0282(.A1(new_n478), .A2(new_n479), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n264), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n469), .A2(new_n476), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G200), .ZN(new_n486));
  INV_X1    g0286(.A(G190), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n464), .B(new_n486), .C1(new_n487), .C2(new_n485), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT21), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n485), .A2(G169), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n464), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n485), .A2(KEYINPUT21), .A3(G169), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n469), .A2(new_n476), .A3(G179), .A4(new_n484), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n457), .A2(new_n461), .A3(new_n463), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT81), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n496), .B1(new_n494), .B2(new_n495), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n488), .B(new_n491), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(G257), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n501));
  OAI211_X1 g0301(.A(G250), .B(new_n248), .C1(new_n249), .C2(new_n250), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G294), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n255), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n475), .A2(G264), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT84), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT84), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n509), .A2(G179), .A3(new_n484), .A4(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n505), .A2(new_n506), .A3(new_n484), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G169), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n335), .A2(KEYINPUT82), .A3(new_n214), .A4(G87), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT22), .ZN(new_n516));
  AOI21_X1  g0316(.A(KEYINPUT83), .B1(new_n380), .B2(G20), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT23), .ZN(new_n518));
  OR2_X1    g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n518), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n515), .A2(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT24), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n214), .A2(KEYINPUT82), .A3(G87), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n304), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(G33), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n525), .A2(new_n449), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n524), .A2(KEYINPUT22), .B1(new_n214), .B2(new_n526), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n521), .A2(new_n522), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n522), .B1(new_n521), .B2(new_n527), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n288), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n459), .A2(new_n380), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT25), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n285), .B2(G107), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n366), .A2(KEYINPUT25), .A3(new_n380), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n514), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n512), .A2(G190), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n509), .A2(new_n484), .A3(new_n510), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n538), .B1(new_n539), .B2(new_n268), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n537), .B1(new_n536), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(G244), .B(new_n248), .C1(new_n249), .C2(new_n250), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT4), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n446), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G250), .A2(G1698), .ZN(new_n546));
  NAND2_X1  g0346(.A1(KEYINPUT4), .A2(G244), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(new_n547), .B2(G1698), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n545), .B1(new_n335), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n258), .B1(new_n544), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(G257), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n478), .A2(new_n479), .A3(new_n481), .A4(new_n482), .ZN(new_n552));
  OAI22_X1  g0352(.A1(new_n474), .A2(new_n551), .B1(new_n552), .B2(new_n342), .ZN(new_n553));
  NOR3_X1   g0353(.A1(new_n550), .A2(new_n553), .A3(G179), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n544), .A2(new_n549), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n255), .ZN(new_n556));
  INV_X1    g0356(.A(new_n553), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT77), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT77), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n550), .B2(new_n553), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n554), .B1(new_n561), .B2(new_n325), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT6), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n563), .A2(new_n447), .A3(G107), .ZN(new_n564));
  XNOR2_X1  g0364(.A(G97), .B(G107), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n564), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  OAI22_X1  g0366(.A1(new_n566), .A2(new_n214), .B1(new_n220), .B2(new_n357), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n380), .B1(new_n303), .B2(new_n305), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n288), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n459), .A2(G97), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n285), .A2(new_n447), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT74), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT74), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n570), .A2(new_n574), .A3(new_n571), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n562), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(KEYINPUT75), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n558), .A2(G190), .A3(new_n560), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT75), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n569), .A2(new_n576), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n556), .A2(new_n557), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G200), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n579), .A2(new_n580), .A3(new_n582), .A4(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(G250), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n480), .B2(G1), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n259), .A2(new_n262), .A3(G45), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n258), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(G238), .A2(G1698), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n590), .B1(new_n221), .B2(G1698), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n526), .B1(new_n591), .B2(new_n335), .ZN(new_n592));
  OAI211_X1 g0392(.A(G190), .B(new_n589), .C1(new_n592), .C2(new_n258), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT78), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n258), .A2(new_n587), .A3(new_n588), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n219), .A2(new_n248), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n221), .A2(G1698), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n596), .B(new_n597), .C1(new_n249), .C2(new_n250), .ZN(new_n598));
  INV_X1    g0398(.A(new_n526), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n595), .B1(new_n600), .B2(new_n255), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT78), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n601), .A2(new_n602), .A3(G190), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n594), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n258), .B1(new_n598), .B2(new_n599), .ZN(new_n605));
  OAI21_X1  g0405(.A(G200), .B1(new_n605), .B2(new_n595), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n404), .A2(new_n285), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT19), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n214), .B1(new_n338), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(G87), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n610), .A2(new_n447), .A3(new_n380), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n214), .B(G68), .C1(new_n249), .C2(new_n250), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n608), .B1(new_n359), .B2(new_n447), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n607), .B1(new_n615), .B2(new_n288), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n459), .A2(new_n610), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n606), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n325), .B1(new_n605), .B2(new_n595), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n386), .B(new_n589), .C1(new_n592), .C2(new_n258), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n616), .B1(new_n459), .B2(new_n405), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n604), .A2(new_n619), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n578), .A2(new_n585), .A3(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n541), .A2(new_n625), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n445), .A2(new_n500), .A3(new_n626), .ZN(G372));
  NAND2_X1  g0427(.A1(new_n622), .A2(new_n623), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT77), .B1(new_n556), .B2(new_n557), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n550), .A2(new_n553), .A3(new_n559), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n325), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n554), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n569), .A2(new_n576), .A3(new_n581), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n581), .B1(new_n569), .B2(new_n576), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT88), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI211_X1 g0438(.A(new_n607), .B(new_n617), .C1(new_n288), .C2(new_n615), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n606), .A2(KEYINPUT85), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n589), .B1(new_n592), .B2(new_n258), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT85), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(new_n642), .A3(G200), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n639), .A2(new_n640), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT86), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n644), .A2(new_n645), .B1(new_n603), .B2(new_n594), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n639), .A2(new_n640), .A3(new_n643), .A4(KEYINPUT86), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n629), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n562), .B(KEYINPUT88), .C1(new_n635), .C2(new_n634), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n638), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n562), .A2(new_n624), .A3(KEYINPUT26), .A4(new_n577), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n653), .B(KEYINPUT89), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n629), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n578), .B(new_n585), .C1(new_n536), .C2(new_n540), .ZN(new_n656));
  INV_X1    g0456(.A(new_n648), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT87), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n578), .A2(new_n585), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT87), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n540), .A2(new_n536), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n659), .A2(new_n660), .A3(new_n661), .A4(new_n648), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n494), .A2(new_n495), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n491), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n537), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n658), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n655), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n445), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g0468(.A(new_n668), .B(KEYINPUT90), .Z(new_n669));
  INV_X1    g0469(.A(new_n443), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT91), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n389), .B2(new_n407), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n406), .A2(new_n288), .ZN(new_n673));
  INV_X1    g0473(.A(new_n391), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n381), .A2(new_n255), .ZN(new_n676));
  INV_X1    g0476(.A(new_n377), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(new_n386), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT71), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n382), .A2(new_n385), .A3(new_n386), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n383), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n675), .A2(new_n681), .A3(KEYINPUT91), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n672), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n376), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n373), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n278), .A2(KEYINPUT17), .A3(new_n312), .ZN(new_n686));
  AOI21_X1  g0486(.A(KEYINPUT17), .B1(new_n278), .B2(new_n312), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n331), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(new_n329), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n439), .A2(new_n440), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n670), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n669), .A2(new_n694), .ZN(G369));
  INV_X1    g0495(.A(new_n664), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n259), .A2(new_n214), .A3(G13), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n697), .A2(KEYINPUT27), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(KEYINPUT27), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G213), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(G343), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n464), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n696), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n499), .B2(new_n704), .ZN(new_n706));
  XNOR2_X1  g0506(.A(KEYINPUT92), .B(G330), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n703), .B1(new_n530), .B2(new_n535), .ZN(new_n710));
  OAI22_X1  g0510(.A1(new_n541), .A2(new_n710), .B1(new_n537), .B2(new_n703), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n514), .A2(new_n536), .A3(new_n703), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n497), .A2(new_n498), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n702), .B1(new_n714), .B2(new_n491), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(new_n537), .A3(new_n661), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n712), .A2(new_n713), .A3(new_n716), .ZN(G399));
  INV_X1    g0517(.A(new_n208), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G41), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n611), .A2(G116), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(G1), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n212), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(new_n720), .ZN(new_n724));
  XOR2_X1   g0524(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n725));
  XNOR2_X1  g0525(.A(new_n724), .B(new_n725), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n537), .B(new_n491), .C1(new_n497), .C2(new_n498), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n727), .A2(new_n659), .A3(new_n661), .A4(new_n648), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n562), .A2(new_n624), .A3(new_n577), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n628), .B1(new_n729), .B2(KEYINPUT26), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n730), .B1(new_n650), .B2(KEYINPUT26), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n728), .B1(new_n731), .B2(KEYINPUT97), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT97), .ZN(new_n733));
  AOI211_X1 g0533(.A(new_n733), .B(new_n730), .C1(new_n650), .C2(KEYINPUT26), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n703), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT98), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT98), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n737), .B(new_n703), .C1(new_n732), .C2(new_n734), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(KEYINPUT29), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n667), .A2(new_n703), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(KEYINPUT96), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT29), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT96), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n667), .A2(new_n744), .A3(new_n703), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n740), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n630), .A2(new_n631), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT84), .ZN(new_n749));
  AOI21_X1  g0549(.A(KEYINPUT84), .B1(new_n505), .B2(new_n506), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n493), .A2(new_n641), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n748), .A2(KEYINPUT30), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT95), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AND4_X1   g0555(.A1(G179), .A2(new_n469), .A3(new_n476), .A4(new_n484), .ZN(new_n756));
  AND4_X1   g0556(.A1(new_n756), .A2(new_n509), .A3(new_n510), .A4(new_n601), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n757), .A2(KEYINPUT95), .A3(KEYINPUT30), .A4(new_n748), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT94), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT30), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n756), .A2(new_n509), .A3(new_n510), .A4(new_n601), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n761), .B1(new_n762), .B2(new_n561), .ZN(new_n763));
  AND4_X1   g0563(.A1(new_n386), .A2(new_n583), .A3(new_n485), .A4(new_n641), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n539), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n759), .B1(new_n760), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n763), .A2(new_n765), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(KEYINPUT94), .ZN(new_n769));
  OAI211_X1 g0569(.A(KEYINPUT31), .B(new_n702), .C1(new_n767), .C2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n626), .A2(new_n500), .A3(new_n703), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT31), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n768), .B1(new_n755), .B2(new_n758), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n772), .B1(new_n773), .B2(new_n703), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n770), .A2(new_n771), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n707), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n747), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n726), .B1(new_n778), .B2(G1), .ZN(G364));
  AND2_X1   g0579(.A1(new_n214), .A2(G13), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n259), .B1(new_n780), .B2(G45), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n720), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n709), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(new_n707), .B2(new_n706), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n208), .A2(G355), .A3(new_n335), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(G116), .B2(new_n208), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n718), .A2(new_n335), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(new_n480), .B2(new_n212), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n242), .A2(new_n480), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n786), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n214), .B1(KEYINPUT99), .B2(new_n325), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n325), .A2(KEYINPUT99), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n213), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G13), .A2(G33), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G20), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n782), .B1(new_n791), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n214), .A2(new_n386), .ZN(new_n801));
  NOR2_X1   g0601(.A1(G190), .A2(G200), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n801), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n804), .A2(new_n487), .A3(G200), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n335), .B1(new_n220), .B2(new_n803), .C1(new_n806), .C2(new_n293), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n804), .A2(new_n487), .A3(new_n268), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(KEYINPUT100), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n808), .A2(KEYINPUT100), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n807), .B1(new_n813), .B2(G50), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n487), .A2(G179), .A3(G200), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n214), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n447), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n804), .A2(new_n268), .A3(G190), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(G68), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT101), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT32), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n214), .A2(G179), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n802), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n821), .B1(new_n824), .B2(G159), .ZN(new_n825));
  INV_X1    g0625(.A(G159), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n823), .A2(KEYINPUT32), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n822), .A2(new_n487), .A3(G200), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n380), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n822), .A2(G190), .A3(G200), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(new_n610), .ZN(new_n831));
  NOR4_X1   g0631(.A1(new_n825), .A2(new_n827), .A3(new_n829), .A4(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n814), .A2(new_n820), .A3(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n816), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n813), .A2(G326), .B1(G294), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(KEYINPUT102), .ZN(new_n836));
  INV_X1    g0636(.A(G317), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(KEYINPUT33), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n837), .A2(KEYINPUT33), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n818), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(G322), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n841), .B2(new_n806), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(G329), .B2(new_n824), .ZN(new_n843));
  INV_X1    g0643(.A(G311), .ZN(new_n844));
  INV_X1    g0644(.A(G303), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n304), .B1(new_n803), .B2(new_n844), .C1(new_n845), .C2(new_n830), .ZN(new_n846));
  INV_X1    g0646(.A(new_n828), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n846), .B1(G283), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n836), .A2(new_n843), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n835), .A2(KEYINPUT102), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n833), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n800), .B1(new_n851), .B2(new_n794), .ZN(new_n852));
  INV_X1    g0652(.A(new_n797), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n852), .B1(new_n706), .B2(new_n853), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n784), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(G396));
  NAND2_X1  g0656(.A1(new_n675), .A2(new_n702), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n407), .A2(new_n411), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n859), .B(KEYINPUT106), .C1(new_n407), .C2(new_n389), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n683), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT106), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n859), .B(new_n862), .C1(new_n407), .C2(new_n389), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n857), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n742), .A2(new_n745), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n857), .B1(new_n672), .B2(new_n682), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n867), .A2(new_n860), .B1(new_n857), .B2(new_n863), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n667), .A2(new_n703), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n782), .B1(new_n870), .B2(new_n776), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n776), .B2(new_n870), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n794), .A2(new_n795), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n782), .B1(G77), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n803), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n818), .A2(G150), .B1(G159), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g0676(.A(KEYINPUT105), .B(G143), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n876), .B1(new_n806), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n813), .B2(G137), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT34), .ZN(new_n880));
  INV_X1    g0680(.A(G132), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n335), .B1(new_n823), .B2(new_n881), .C1(new_n816), .C2(new_n293), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n202), .A2(new_n830), .B1(new_n828), .B2(new_n218), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n818), .ZN(new_n885));
  XNOR2_X1  g0685(.A(KEYINPUT103), .B(G283), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n885), .A2(new_n886), .B1(new_n803), .B2(new_n449), .ZN(new_n887));
  INV_X1    g0687(.A(G294), .ZN(new_n888));
  OAI22_X1  g0688(.A1(new_n806), .A2(new_n888), .B1(new_n823), .B2(new_n844), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n828), .A2(new_n610), .ZN(new_n890));
  NOR4_X1   g0690(.A1(new_n887), .A2(new_n889), .A3(new_n817), .A4(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n845), .B2(new_n812), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n304), .B1(new_n830), .B2(new_n380), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n893), .B(KEYINPUT104), .Z(new_n894));
  OAI22_X1  g0694(.A1(new_n880), .A2(new_n884), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n874), .B1(new_n895), .B2(new_n794), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n868), .B2(new_n796), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n872), .A2(new_n897), .ZN(G384));
  INV_X1    g0698(.A(new_n566), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n899), .A2(KEYINPUT35), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(KEYINPUT35), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n900), .A2(G116), .A3(new_n215), .A4(new_n901), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n902), .B(KEYINPUT36), .Z(new_n903));
  OAI211_X1 g0703(.A(new_n212), .B(G77), .C1(new_n293), .C2(new_n218), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n202), .A2(G68), .ZN(new_n905));
  AOI211_X1 g0705(.A(new_n259), .B(G13), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n740), .A2(new_n445), .A3(new_n746), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n908), .A2(new_n694), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT110), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n356), .A2(new_n372), .A3(new_n703), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT38), .ZN(new_n913));
  INV_X1    g0713(.A(new_n700), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n323), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n688), .B2(new_n691), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT37), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n323), .B1(new_n328), .B2(new_n914), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n313), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n917), .B1(new_n313), .B2(new_n918), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n913), .B1(new_n916), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n323), .B1(new_n270), .B2(new_n277), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n326), .B1(G179), .B2(new_n276), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT108), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n310), .B2(new_n298), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n319), .A2(KEYINPUT108), .A3(new_n320), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n927), .A2(new_n928), .A3(new_n309), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n308), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n925), .B1(new_n930), .B2(new_n290), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n700), .B1(new_n930), .B2(new_n290), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n924), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n919), .B1(new_n933), .B2(new_n917), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n333), .A2(new_n932), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT38), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT109), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT39), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n923), .A2(new_n936), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n923), .A2(new_n936), .A3(new_n938), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(KEYINPUT109), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n924), .A2(new_n931), .ZN(new_n942));
  INV_X1    g0742(.A(new_n932), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n920), .B1(new_n944), .B2(KEYINPUT37), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n943), .B1(new_n688), .B2(new_n691), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n913), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n938), .B1(new_n947), .B2(new_n936), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n912), .B(new_n939), .C1(new_n941), .C2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n936), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n372), .A2(new_n702), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n373), .A2(new_n376), .A3(new_n951), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n372), .B(new_n702), .C1(new_n684), .C2(new_n356), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI211_X1 g0754(.A(new_n702), .B(new_n865), .C1(new_n655), .C2(new_n666), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n408), .A2(new_n703), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT107), .Z(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n950), .B(new_n954), .C1(new_n955), .C2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n691), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n700), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n949), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n910), .B(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n923), .A2(new_n936), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n954), .A2(new_n868), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n772), .B(new_n703), .C1(new_n759), .C2(new_n766), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT111), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n967), .B1(new_n774), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n759), .A2(new_n766), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n970), .A2(new_n968), .A3(KEYINPUT31), .A4(new_n702), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n771), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n965), .B(new_n966), .C1(new_n969), .C2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n954), .A2(new_n868), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n771), .A2(new_n971), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n970), .A2(KEYINPUT31), .A3(new_n702), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT31), .B1(new_n970), .B2(new_n702), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n976), .B1(new_n977), .B2(KEYINPUT111), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n974), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(KEYINPUT40), .B1(new_n947), .B2(new_n936), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n973), .A2(KEYINPUT40), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n975), .A2(new_n978), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n445), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n981), .B(new_n983), .Z(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n707), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n964), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n259), .B2(new_n780), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n964), .A2(new_n985), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n907), .B1(new_n987), .B2(new_n988), .ZN(G367));
  NOR2_X1   g0789(.A1(new_n788), .A2(new_n238), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n798), .B1(new_n208), .B2(new_n405), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n782), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n335), .B1(new_n293), .B2(new_n830), .C1(new_n885), .C2(new_n826), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n828), .A2(new_n220), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n816), .A2(new_n218), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(G150), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n806), .A2(new_n997), .B1(new_n803), .B2(new_n202), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G137), .B2(new_n824), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n996), .B(new_n999), .C1(new_n812), .C2(new_n877), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n805), .A2(G303), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n837), .B2(new_n823), .C1(new_n885), .C2(new_n888), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT46), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n830), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(G116), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1002), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n1003), .B2(new_n1005), .C1(new_n844), .C2(new_n812), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n886), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n335), .B1(new_n875), .B2(new_n1008), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n447), .B2(new_n828), .C1(new_n380), .C2(new_n816), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1000), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT47), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n992), .B1(new_n1012), .B2(new_n794), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n639), .A2(new_n703), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n628), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n648), .B2(new_n1014), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT112), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n797), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n781), .B(KEYINPUT114), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n716), .B1(new_n711), .B2(new_n715), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(new_n708), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n777), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n716), .A2(new_n713), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n636), .A2(new_n703), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n702), .B1(new_n634), .B2(new_n635), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1025), .B1(new_n659), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT45), .ZN(new_n1029));
  AOI21_X1  g0829(.A(KEYINPUT44), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1024), .A2(KEYINPUT44), .A3(new_n1027), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AND3_X1   g0833(.A1(new_n1029), .A2(new_n712), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n712), .B1(new_n1029), .B2(new_n1033), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1023), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n778), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n719), .B(KEYINPUT41), .Z(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1020), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT43), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1017), .A2(new_n1042), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n716), .A2(new_n1027), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1044), .A2(KEYINPUT42), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n578), .B1(new_n1027), .B2(new_n537), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n703), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1044), .A2(KEYINPUT42), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1045), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT113), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1017), .A2(new_n1042), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1050), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1043), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(KEYINPUT113), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1043), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(new_n1058), .A3(new_n1052), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1055), .A2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n712), .A2(new_n1027), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1060), .B(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1019), .B1(new_n1041), .B2(new_n1063), .ZN(G387));
  INV_X1    g0864(.A(new_n1023), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n777), .A2(new_n1022), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1065), .A2(new_n719), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n721), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n208), .A2(new_n335), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n395), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n202), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT50), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n480), .B1(new_n218), .B2(new_n220), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n1072), .A2(new_n1068), .A3(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n787), .B1(new_n235), .B2(new_n480), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1069), .B1(G107), .B2(new_n208), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n798), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1077), .B(new_n782), .C1(new_n711), .C2(new_n853), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n806), .A2(new_n202), .B1(new_n803), .B2(new_n218), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n304), .B(new_n1079), .C1(G150), .C2(new_n824), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n828), .A2(new_n447), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n830), .A2(new_n220), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1081), .B(new_n1082), .C1(new_n404), .C2(new_n834), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n813), .A2(G159), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n284), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n818), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1080), .A2(new_n1083), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n813), .A2(G322), .B1(G311), .B2(new_n818), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1088), .A2(KEYINPUT115), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(KEYINPUT115), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n805), .A2(G317), .B1(G303), .B2(new_n875), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT48), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n834), .A2(new_n1008), .B1(new_n1004), .B2(G294), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT49), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(KEYINPUT116), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n828), .A2(new_n449), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n335), .B(new_n1100), .C1(G326), .C2(new_n824), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1098), .A2(KEYINPUT116), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1087), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1078), .B1(new_n1104), .B2(new_n794), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1022), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1105), .B1(new_n1106), .B2(new_n1020), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1067), .A2(new_n1107), .ZN(G393));
  AOI21_X1  g0908(.A(new_n720), .B1(new_n1023), .B2(new_n1036), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n1023), .B2(new_n1036), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1036), .A2(new_n1020), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n788), .A2(new_n245), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n798), .B1(new_n208), .B2(new_n447), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n782), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n812), .A2(new_n837), .B1(new_n844), .B2(new_n806), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT52), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n818), .A2(G303), .B1(G294), .B2(new_n875), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n449), .B2(new_n816), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT117), .Z(new_n1119));
  OAI21_X1  g0919(.A(new_n304), .B1(new_n823), .B2(new_n841), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n829), .B(new_n1120), .C1(new_n1004), .C2(new_n1008), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1116), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n812), .A2(new_n997), .B1(new_n826), .B2(new_n806), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT51), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n830), .A2(new_n218), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n890), .B(new_n1125), .C1(G77), .C2(new_n834), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n335), .B1(new_n823), .B2(new_n877), .C1(new_n885), .C2(new_n202), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n1070), .B2(new_n875), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1124), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1122), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1114), .B1(new_n1130), .B2(new_n794), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1027), .A2(new_n797), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1110), .A2(new_n1111), .A3(new_n1133), .ZN(G390));
  INV_X1    g0934(.A(G330), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n975), .B2(new_n978), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n445), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n908), .A2(new_n694), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n865), .B1(new_n736), .B2(new_n738), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1139), .A2(new_n958), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n954), .B1(new_n1136), .B2(new_n868), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n775), .A2(new_n707), .A3(new_n868), .A4(new_n954), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n869), .A2(new_n957), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n954), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n776), .B2(new_n865), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1136), .A2(new_n966), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1140), .A2(new_n1144), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1138), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1136), .A2(new_n966), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1142), .B1(new_n1153), .B2(KEYINPUT118), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n954), .B1(new_n955), .B2(new_n958), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n936), .ZN(new_n1156));
  AOI21_X1  g0956(.A(KEYINPUT38), .B1(new_n934), .B2(new_n935), .ZN(new_n1157));
  OAI21_X1  g0957(.A(KEYINPUT39), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1158), .A2(KEYINPUT109), .A3(new_n940), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1155), .A2(new_n911), .B1(new_n1159), .B2(new_n939), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n954), .B1(new_n1139), .B2(new_n958), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n965), .A2(new_n911), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1154), .B(new_n1160), .C1(new_n1161), .C2(new_n1163), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1148), .A2(KEYINPUT118), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1160), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1152), .B1(new_n1164), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1160), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1154), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1151), .B(new_n1172), .C1(new_n1170), .C2(new_n1165), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1169), .A2(new_n719), .A3(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1164), .A2(new_n1168), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1159), .A2(new_n939), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n795), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n782), .B1(new_n1085), .B2(new_n873), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n813), .A2(G283), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n335), .B(new_n831), .C1(G116), .C2(new_n805), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n834), .A2(G77), .B1(new_n847), .B2(G68), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n885), .A2(new_n380), .B1(new_n823), .B2(new_n888), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G97), .B2(new_n875), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .A4(new_n1183), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n818), .A2(G137), .B1(G125), .B2(new_n824), .ZN(new_n1185));
  INV_X1    g0985(.A(G128), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1185), .B1(new_n881), .B2(new_n806), .C1(new_n812), .C2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n828), .A2(new_n202), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(KEYINPUT54), .B(G143), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n335), .B1(new_n803), .B2(new_n1189), .C1(new_n816), .C2(new_n826), .ZN(new_n1190));
  OR3_X1    g0990(.A1(new_n1187), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1004), .A2(G150), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT53), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1184), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1178), .B1(new_n1194), .B2(new_n794), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1175), .A2(new_n1020), .B1(new_n1177), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1174), .A2(new_n1196), .ZN(G378));
  INV_X1    g0997(.A(KEYINPUT120), .ZN(new_n1198));
  XOR2_X1   g0998(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n444), .A2(new_n442), .A3(new_n914), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT119), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n442), .A2(new_n914), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n439), .A2(new_n440), .A3(new_n443), .A4(new_n1203), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1201), .A2(new_n1202), .A3(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1202), .B1(new_n1201), .B2(new_n1204), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1200), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1201), .A2(new_n1204), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(KEYINPUT119), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1201), .A2(new_n1202), .A3(new_n1204), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1209), .A2(new_n1199), .A3(new_n1210), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1207), .A2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n981), .B2(new_n1135), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1207), .A2(new_n1211), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT40), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n979), .B2(new_n965), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n980), .A2(new_n982), .A3(new_n966), .ZN(new_n1217));
  OAI211_X1 g1017(.A(G330), .B(new_n1214), .C1(new_n1216), .C2(new_n1217), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n962), .A2(new_n1213), .A3(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1146), .B1(new_n869), .B2(new_n957), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1220), .A2(new_n950), .B1(new_n960), .B2(new_n700), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1213), .A2(new_n1218), .B1(new_n1221), .B2(new_n949), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1198), .B1(new_n1219), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1213), .A2(new_n1218), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n963), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n962), .A2(new_n1213), .A3(new_n1218), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1225), .A2(KEYINPUT120), .A3(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1223), .A2(new_n1227), .A3(new_n1020), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n782), .B1(G50), .B2(new_n873), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n304), .B2(new_n470), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n470), .B(new_n304), .C1(new_n885), .C2(new_n447), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n828), .A2(new_n293), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(new_n1232), .A2(new_n995), .A3(new_n1082), .A4(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(G283), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n806), .A2(new_n380), .B1(new_n823), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n404), .B2(new_n875), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1234), .B(new_n1237), .C1(new_n449), .C2(new_n812), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT58), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1231), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n813), .A2(G125), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n1186), .A2(new_n806), .B1(new_n885), .B2(new_n881), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G137), .B2(new_n875), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1189), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n834), .A2(G150), .B1(new_n1004), .B2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1241), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(KEYINPUT59), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n847), .A2(G159), .ZN(new_n1248));
  AOI211_X1 g1048(.A(G33), .B(G41), .C1(new_n824), .C2(G124), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1246), .A2(KEYINPUT59), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n1240), .B1(new_n1239), .B2(new_n1238), .C1(new_n1250), .C2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1229), .B1(new_n1252), .B2(new_n794), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n1214), .B2(new_n796), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1228), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT122), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1138), .B1(new_n1175), .B2(new_n1151), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT121), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1225), .A2(new_n1258), .A3(new_n1226), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1222), .A2(KEYINPUT121), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(KEYINPUT57), .A3(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1256), .B1(new_n1257), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1138), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1173), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1261), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1264), .A2(new_n1265), .A3(KEYINPUT122), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1262), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1223), .A2(new_n1227), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(new_n1263), .B2(new_n1173), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n719), .B1(new_n1269), .B2(KEYINPUT57), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1255), .B1(new_n1267), .B2(new_n1270), .ZN(G375));
  NAND2_X1  g1071(.A1(new_n1138), .A2(new_n1150), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1152), .A2(new_n1040), .A3(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n782), .B1(G68), .B2(new_n873), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n813), .A2(G294), .ZN(new_n1275));
  AOI211_X1 g1075(.A(new_n335), .B(new_n994), .C1(G116), .C2(new_n818), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n834), .A2(new_n404), .B1(new_n1004), .B2(G97), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n806), .A2(new_n1235), .B1(new_n823), .B2(new_n845), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(G107), .B2(new_n875), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .A4(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n813), .A2(G132), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n304), .B1(new_n818), .B2(new_n1244), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n805), .A2(G137), .B1(G150), .B2(new_n875), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1233), .B1(G50), .B2(new_n834), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .A4(new_n1284), .ZN(new_n1285));
  OAI22_X1  g1085(.A1(new_n830), .A2(new_n826), .B1(new_n823), .B2(new_n1186), .ZN(new_n1286));
  XOR2_X1   g1086(.A(new_n1286), .B(KEYINPUT123), .Z(new_n1287));
  OAI21_X1  g1087(.A(new_n1280), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1274), .B1(new_n1288), .B2(new_n794), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1289), .B1(new_n954), .B2(new_n796), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1020), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1290), .B1(new_n1150), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1273), .A2(new_n1293), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(new_n1294), .B(KEYINPUT124), .ZN(G381));
  INV_X1    g1095(.A(G390), .ZN(new_n1296));
  INV_X1    g1096(.A(G384), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1067), .A2(new_n855), .A3(new_n1107), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1296), .A2(new_n1297), .A3(new_n1299), .ZN(new_n1300));
  OR3_X1    g1100(.A1(new_n1300), .A2(G387), .A3(G378), .ZN(new_n1301));
  OR3_X1    g1101(.A1(new_n1301), .A2(G375), .A3(G381), .ZN(G407));
  INV_X1    g1102(.A(G378), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n701), .A2(G213), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  OAI211_X1 g1105(.A(G407), .B(G213), .C1(G375), .C2(new_n1305), .ZN(G409));
  OAI211_X1 g1106(.A(G378), .B(new_n1255), .C1(new_n1267), .C2(new_n1270), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1269), .A2(new_n1040), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1259), .A2(new_n1020), .A3(new_n1260), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1308), .A2(new_n1254), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n1303), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1304), .B1(new_n1307), .B2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1138), .A2(new_n1150), .A3(KEYINPUT60), .ZN(new_n1313));
  AND2_X1   g1113(.A1(new_n1313), .A2(new_n719), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT60), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1272), .B1(new_n1151), .B2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1293), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1297), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1317), .A2(G384), .A3(new_n1293), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1319), .A2(G2897), .A3(new_n1304), .A4(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1304), .A2(G2897), .ZN(new_n1322));
  AOI21_X1  g1122(.A(G384), .B1(new_n1317), .B2(new_n1293), .ZN(new_n1323));
  AOI211_X1 g1123(.A(new_n1292), .B(new_n1297), .C1(new_n1314), .C2(new_n1316), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1322), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(KEYINPUT125), .B1(new_n1321), .B2(new_n1325), .ZN(new_n1326));
  AND3_X1   g1126(.A1(new_n1321), .A2(KEYINPUT125), .A3(new_n1325), .ZN(new_n1327));
  OR3_X1    g1127(.A1(new_n1312), .A2(new_n1326), .A3(new_n1327), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1312), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT63), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1312), .A2(KEYINPUT63), .A3(new_n1329), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(G387), .A2(new_n1296), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(G387), .A2(new_n1296), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n855), .B1(new_n1067), .B2(new_n1107), .ZN(new_n1337));
  OAI22_X1  g1137(.A1(new_n1335), .A2(new_n1336), .B1(new_n1299), .B2(new_n1337), .ZN(new_n1338));
  OR2_X1    g1138(.A1(G387), .A2(new_n1296), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1299), .A2(new_n1337), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1339), .A2(new_n1340), .A3(new_n1334), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1338), .A2(new_n1341), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1342), .A2(KEYINPUT61), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1328), .A2(new_n1332), .A3(new_n1333), .A4(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT62), .ZN(new_n1345));
  AND3_X1   g1145(.A1(new_n1312), .A2(new_n1345), .A3(new_n1329), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT61), .ZN(new_n1347));
  AND2_X1   g1147(.A1(new_n1321), .A2(new_n1325), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1347), .B1(new_n1312), .B2(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1345), .B1(new_n1312), .B2(new_n1329), .ZN(new_n1350));
  NOR3_X1   g1150(.A1(new_n1346), .A2(new_n1349), .A3(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1342), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1344), .B1(new_n1351), .B2(new_n1352), .ZN(G405));
  INV_X1    g1153(.A(KEYINPUT126), .ZN(new_n1354));
  OR3_X1    g1154(.A1(new_n1329), .A2(new_n1354), .A3(KEYINPUT127), .ZN(new_n1355));
  OAI21_X1  g1155(.A(KEYINPUT127), .B1(new_n1329), .B2(new_n1354), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1342), .A2(new_n1355), .A3(new_n1356), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1342), .B1(new_n1356), .B2(new_n1355), .ZN(new_n1359));
  AND2_X1   g1159(.A1(G375), .A2(new_n1303), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1329), .A2(new_n1354), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1307), .A2(new_n1361), .ZN(new_n1362));
  OAI22_X1  g1162(.A1(new_n1358), .A2(new_n1359), .B1(new_n1360), .B2(new_n1362), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1352), .A2(new_n1364), .ZN(new_n1365));
  NOR2_X1   g1165(.A1(new_n1360), .A2(new_n1362), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1365), .A2(new_n1366), .A3(new_n1357), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1363), .A2(new_n1367), .ZN(G402));
endmodule


