//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n550, new_n551, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n616,
    new_n617, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n768, new_n769, new_n771,
    new_n772, new_n774, new_n775, new_n776, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n823, new_n824;
  XNOR2_X1  g000(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G99gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT68), .ZN(new_n205));
  XNOR2_X1  g004(.A(G15gat), .B(G43gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT27), .B(G183gat), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI22_X1  g009(.A1(new_n210), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n211));
  INV_X1    g010(.A(G169gat), .ZN(new_n212));
  INV_X1    g011(.A(G176gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  XOR2_X1   g014(.A(new_n215), .B(KEYINPUT26), .Z(new_n216));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G183gat), .Z(new_n217));
  MUX2_X1   g016(.A(G183gat), .B(new_n217), .S(KEYINPUT27), .Z(new_n218));
  OR2_X1    g017(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n219));
  OAI221_X1 g018(.A(new_n211), .B1(new_n214), .B2(new_n216), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n214), .B1(KEYINPUT23), .B2(new_n215), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(KEYINPUT23), .B2(new_n215), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(KEYINPUT25), .ZN(new_n223));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(KEYINPUT24), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G183gat), .B2(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n217), .A2(new_n209), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n228), .A2(new_n225), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT25), .B1(new_n229), .B2(new_n222), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n220), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G113gat), .ZN(new_n232));
  INV_X1    g031(.A(G120gat), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT1), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(new_n232), .B2(new_n233), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT65), .ZN(new_n236));
  XNOR2_X1  g035(.A(G127gat), .B(G134gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n231), .B(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(G227gat), .A3(G233gat), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT33), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n207), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(new_n243), .B2(new_n242), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n240), .A2(KEYINPUT32), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT67), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n207), .A2(new_n241), .ZN(new_n248));
  OAI22_X1  g047(.A1(new_n245), .A2(new_n247), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n239), .B1(G227gat), .B2(G233gat), .ZN(new_n250));
  OR2_X1    g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n249), .A2(new_n250), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n203), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n249), .A2(new_n250), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n251), .A2(new_n255), .A3(new_n202), .ZN(new_n256));
  INV_X1    g055(.A(G226gat), .ZN(new_n257));
  INV_X1    g056(.A(G233gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n231), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n259), .A2(KEYINPUT29), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n261), .B1(new_n231), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G197gat), .B(G204gat), .ZN(new_n264));
  AND2_X1   g063(.A1(G211gat), .A2(G218gat), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n264), .B1(KEYINPUT22), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G211gat), .B(G218gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(new_n268), .B(KEYINPUT70), .Z(new_n269));
  OR2_X1    g068(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n263), .A2(new_n269), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(G64gat), .B(G92gat), .Z(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT71), .ZN(new_n274));
  XNOR2_X1  g073(.A(G8gat), .B(G36gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(new_n276), .B(KEYINPUT72), .Z(new_n277));
  OAI21_X1  g076(.A(KEYINPUT30), .B1(new_n272), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n272), .A2(new_n276), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n272), .A2(KEYINPUT30), .A3(new_n276), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n281), .A2(KEYINPUT73), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(KEYINPUT73), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n280), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G1gat), .B(G29gat), .ZN(new_n285));
  INV_X1    g084(.A(G85gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT0), .B(G57gat), .ZN(new_n288));
  XOR2_X1   g087(.A(new_n287), .B(new_n288), .Z(new_n289));
  XNOR2_X1  g088(.A(G141gat), .B(G148gat), .ZN(new_n290));
  OR2_X1    g089(.A1(new_n290), .A2(KEYINPUT2), .ZN(new_n291));
  NAND2_X1  g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292));
  OR2_X1    g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n293), .A2(KEYINPUT74), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(KEYINPUT74), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n291), .A2(new_n292), .A3(new_n294), .A4(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(KEYINPUT75), .B(G162gat), .Z(new_n297));
  INV_X1    g096(.A(G155gat), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT2), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n290), .B1(new_n292), .B2(new_n293), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  OR2_X1    g101(.A1(new_n238), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT78), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n303), .A2(new_n304), .A3(KEYINPUT4), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n302), .A2(KEYINPUT3), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n302), .A2(KEYINPUT3), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n308), .A3(new_n238), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n303), .B(KEYINPUT4), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n305), .B(new_n309), .C1(new_n310), .C2(new_n304), .ZN(new_n311));
  NAND2_X1  g110(.A1(G225gat), .A2(G233gat), .ZN(new_n312));
  XOR2_X1   g111(.A(new_n312), .B(KEYINPUT76), .Z(new_n313));
  NOR3_X1   g112(.A1(new_n311), .A2(KEYINPUT5), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT79), .ZN(new_n315));
  OR2_X1    g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n315), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n313), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n310), .A2(new_n309), .A3(new_n319), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n320), .A2(KEYINPUT77), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(KEYINPUT77), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT5), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n238), .B(new_n302), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n323), .B1(new_n324), .B2(new_n313), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n321), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n289), .B1(new_n318), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT6), .ZN(new_n329));
  INV_X1    g128(.A(new_n289), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n316), .A2(new_n330), .A3(new_n326), .A4(new_n317), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n328), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  OAI211_X1 g131(.A(KEYINPUT6), .B(new_n289), .C1(new_n318), .C2(new_n327), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n284), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n269), .B1(KEYINPUT29), .B2(new_n306), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n268), .A2(KEYINPUT29), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n302), .B1(new_n336), .B2(KEYINPUT3), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT82), .B1(new_n338), .B2(KEYINPUT81), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(G22gat), .ZN(new_n340));
  XOR2_X1   g139(.A(G50gat), .B(G78gat), .Z(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G228gat), .A2(G233gat), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n343), .B1(new_n338), .B2(KEYINPUT82), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(G106gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n344), .B(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n342), .B(new_n347), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n254), .A2(new_n256), .A3(new_n334), .A4(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT35), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n270), .A2(new_n271), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n352), .A2(KEYINPUT37), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT85), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n276), .B1(new_n352), .B2(KEYINPUT37), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT38), .ZN(new_n357));
  OR2_X1    g156(.A1(new_n352), .A2(KEYINPUT84), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT37), .ZN(new_n359));
  INV_X1    g158(.A(new_n270), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n359), .B1(new_n360), .B2(KEYINPUT84), .ZN(new_n361));
  AOI211_X1 g160(.A(KEYINPUT38), .B(new_n277), .C1(new_n358), .C2(new_n361), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n362), .A2(new_n354), .B1(new_n272), .B2(new_n276), .ZN(new_n363));
  AND4_X1   g162(.A1(new_n333), .A2(new_n357), .A3(new_n363), .A4(new_n332), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n311), .A2(new_n313), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n330), .B1(new_n365), .B2(KEYINPUT39), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT40), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT39), .B1(new_n324), .B2(new_n313), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n368), .B1(new_n311), .B2(new_n313), .ZN(new_n369));
  OR3_X1    g168(.A1(new_n366), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n284), .A2(new_n328), .A3(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n367), .B1(new_n366), .B2(new_n369), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(KEYINPUT83), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n348), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  OAI22_X1  g173(.A1(new_n364), .A2(new_n374), .B1(new_n334), .B2(new_n348), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n254), .A2(KEYINPUT36), .A3(new_n256), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n254), .A2(new_n256), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT36), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n375), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT86), .B1(new_n351), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n349), .B(KEYINPUT35), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n379), .A2(new_n376), .ZN(new_n383));
  INV_X1    g182(.A(new_n375), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT86), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n382), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT15), .ZN(new_n388));
  XNOR2_X1  g187(.A(G43gat), .B(G50gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT87), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n388), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(KEYINPUT87), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  XOR2_X1   g193(.A(KEYINPUT89), .B(G29gat), .Z(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(G36gat), .ZN(new_n396));
  OR3_X1    g195(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n390), .A2(new_n388), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n394), .A2(new_n396), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT88), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n398), .B1(new_n397), .B2(new_n402), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n396), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(new_n393), .A3(new_n392), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT17), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G15gat), .B(G22gat), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT16), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n410), .B1(new_n411), .B2(G1gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n412), .B(new_n413), .C1(G1gat), .C2(new_n410), .ZN(new_n414));
  NOR2_X1   g213(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n406), .A3(KEYINPUT17), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n409), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G229gat), .A2(G233gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT91), .ZN(new_n420));
  INV_X1    g219(.A(new_n416), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n407), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n418), .A2(KEYINPUT18), .A3(new_n420), .A4(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n420), .B(KEYINPUT13), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n421), .A2(new_n407), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n416), .B1(new_n406), .B2(new_n401), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n417), .A2(new_n416), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT17), .B1(new_n401), .B2(new_n406), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n422), .B(new_n420), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT18), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT92), .ZN(new_n436));
  XNOR2_X1  g235(.A(G113gat), .B(G141gat), .ZN(new_n437));
  INV_X1    g236(.A(G197gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(KEYINPUT11), .B(G169gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(KEYINPUT12), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n430), .B(new_n435), .C1(new_n436), .C2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n423), .A2(new_n436), .A3(new_n428), .ZN(new_n444));
  INV_X1    g243(.A(new_n442), .ZN(new_n445));
  INV_X1    g244(.A(new_n435), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n444), .B(new_n445), .C1(new_n446), .C2(new_n429), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G134gat), .B(G162gat), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT95), .ZN(new_n453));
  NAND2_X1  g252(.A1(G85gat), .A2(G92gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(KEYINPUT7), .ZN(new_n455));
  NAND2_X1  g254(.A1(G99gat), .A2(G106gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT8), .ZN(new_n457));
  OR2_X1    g256(.A1(G85gat), .A2(G92gat), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n457), .A2(KEYINPUT94), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT94), .B1(new_n457), .B2(new_n458), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n455), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  XOR2_X1   g260(.A(G99gat), .B(G106gat), .Z(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n462), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n464), .B(new_n455), .C1(new_n459), .C2(new_n460), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n453), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT7), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n454), .B(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n457), .A2(new_n458), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT94), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT94), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n468), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT95), .B1(new_n473), .B2(new_n464), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n409), .B(new_n417), .C1(new_n466), .C2(new_n474), .ZN(new_n475));
  AND3_X1   g274(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n463), .A2(new_n465), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n474), .B1(new_n477), .B2(KEYINPUT95), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n476), .B1(new_n478), .B2(new_n407), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(G190gat), .B(G218gat), .ZN(new_n481));
  XOR2_X1   g280(.A(new_n481), .B(KEYINPUT96), .Z(new_n482));
  AOI21_X1  g281(.A(new_n452), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n482), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n475), .A2(new_n484), .A3(new_n479), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT98), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT97), .B1(new_n480), .B2(new_n482), .ZN(new_n488));
  OR2_X1    g287(.A1(new_n488), .A2(new_n485), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n485), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n452), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G57gat), .B(G64gat), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G71gat), .B(G78gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n497), .A2(KEYINPUT21), .ZN(new_n498));
  XOR2_X1   g297(.A(G127gat), .B(G155gat), .Z(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n501));
  XNOR2_X1  g300(.A(G183gat), .B(G211gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n500), .B(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n421), .B1(KEYINPUT21), .B2(new_n497), .ZN(new_n505));
  NAND2_X1  g304(.A1(G231gat), .A2(G233gat), .ZN(new_n506));
  XOR2_X1   g305(.A(new_n506), .B(KEYINPUT93), .Z(new_n507));
  XNOR2_X1  g306(.A(new_n505), .B(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(new_n504), .B(new_n508), .Z(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G120gat), .B(G148gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(G176gat), .B(G204gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n513), .B(KEYINPUT100), .Z(new_n514));
  NAND2_X1  g313(.A1(G230gat), .A2(G233gat), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT99), .B1(new_n478), .B2(new_n497), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT10), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n497), .A2(new_n465), .A3(new_n463), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT99), .ZN(new_n520));
  INV_X1    g319(.A(new_n497), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n520), .B(new_n521), .C1(new_n466), .C2(new_n474), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n517), .A2(new_n518), .A3(new_n519), .A4(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n478), .A2(KEYINPUT10), .A3(new_n497), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n516), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n522), .A2(new_n519), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n515), .B1(new_n526), .B2(new_n517), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n514), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT101), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g329(.A(KEYINPUT101), .B(new_n514), .C1(new_n525), .C2(new_n527), .ZN(new_n531));
  OR3_X1    g330(.A1(new_n525), .A2(new_n527), .A3(new_n513), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NOR3_X1   g332(.A1(new_n492), .A2(new_n510), .A3(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n381), .A2(new_n387), .A3(new_n448), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n332), .A2(new_n333), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n537), .B(G1gat), .Z(G1324gat));
  INV_X1    g337(.A(KEYINPUT104), .ZN(new_n539));
  INV_X1    g338(.A(new_n284), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT16), .B(G8gat), .ZN(new_n541));
  OR3_X1    g340(.A1(new_n535), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n539), .B1(new_n542), .B2(KEYINPUT102), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT42), .ZN(new_n544));
  OAI21_X1  g343(.A(G8gat), .B1(new_n535), .B2(new_n540), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT103), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT42), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n547), .B1(new_n542), .B2(new_n539), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n544), .B(new_n546), .C1(new_n543), .C2(new_n548), .ZN(G1325gat));
  NOR2_X1   g348(.A1(new_n535), .A2(new_n377), .ZN(new_n550));
  INV_X1    g349(.A(new_n383), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(G15gat), .ZN(new_n552));
  OAI22_X1  g351(.A1(new_n550), .A2(G15gat), .B1(new_n535), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT105), .ZN(G1326gat));
  NOR2_X1   g353(.A1(new_n535), .A2(new_n348), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT106), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT43), .B(G22gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(G1327gat));
  INV_X1    g357(.A(new_n533), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n492), .A2(new_n510), .A3(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT107), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n381), .A2(new_n387), .A3(new_n448), .A4(new_n561), .ZN(new_n562));
  NOR3_X1   g361(.A1(new_n562), .A2(new_n536), .A3(new_n395), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n563), .B(KEYINPUT45), .Z(new_n564));
  NAND2_X1  g363(.A1(new_n382), .A2(new_n385), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n492), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT44), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n381), .A2(new_n387), .A3(KEYINPUT44), .A4(new_n492), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n536), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n559), .A2(KEYINPUT108), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n559), .A2(KEYINPUT108), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n448), .ZN(new_n576));
  NOR3_X1   g375(.A1(new_n575), .A2(new_n576), .A3(new_n509), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n570), .A2(new_n571), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n395), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n579), .ZN(G1328gat));
  NAND4_X1  g379(.A1(new_n568), .A2(new_n569), .A3(new_n284), .A4(new_n577), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(G36gat), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n540), .A2(G36gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  OR3_X1    g383(.A1(new_n562), .A2(KEYINPUT46), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT46), .B1(new_n562), .B2(new_n584), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n582), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT109), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n582), .A2(new_n585), .A3(KEYINPUT109), .A4(new_n586), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(G1329gat));
  NAND4_X1  g390(.A1(new_n570), .A2(G43gat), .A3(new_n551), .A4(new_n577), .ZN(new_n592));
  INV_X1    g391(.A(G43gat), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n593), .B1(new_n562), .B2(new_n377), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n592), .A2(KEYINPUT47), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT47), .B1(new_n592), .B2(new_n594), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(G1330gat));
  INV_X1    g396(.A(new_n348), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n568), .A2(new_n569), .A3(new_n598), .A4(new_n577), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(G50gat), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT110), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT48), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OR3_X1    g401(.A1(new_n562), .A2(G50gat), .A3(new_n348), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n600), .B(new_n603), .C1(new_n601), .C2(KEYINPUT48), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(G1331gat));
  INV_X1    g406(.A(new_n492), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n608), .A2(new_n576), .A3(new_n509), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n574), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(KEYINPUT111), .Z(new_n611));
  NAND2_X1  g410(.A1(new_n565), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n571), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g414(.A(new_n540), .B(new_n612), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n616));
  NOR2_X1   g415(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(G1333gat));
  INV_X1    g417(.A(G71gat), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n619), .B1(new_n612), .B2(new_n377), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n613), .A2(G71gat), .A3(new_n551), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n621), .A2(KEYINPUT112), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(KEYINPUT112), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n620), .B(new_n625), .C1(new_n622), .C2(new_n623), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(G1334gat));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n598), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G78gat), .ZN(G1335gat));
  NAND4_X1  g430(.A1(new_n565), .A2(new_n576), .A3(new_n510), .A4(new_n492), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT51), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n536), .A2(G85gat), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(new_n533), .A3(new_n635), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n559), .A2(new_n448), .A3(new_n509), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n568), .A2(new_n569), .A3(new_n571), .A4(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(G85gat), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT114), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n636), .A2(KEYINPUT114), .A3(new_n639), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(G1336gat));
  NAND2_X1  g443(.A1(new_n575), .A2(new_n284), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(G92gat), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n634), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n568), .A2(new_n569), .A3(new_n284), .A4(new_n637), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(G92gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT52), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT52), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n647), .A2(new_n652), .A3(new_n649), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(G1337gat));
  NAND3_X1  g453(.A1(new_n570), .A2(new_n551), .A3(new_n637), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(G99gat), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n377), .A2(G99gat), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n634), .A2(new_n533), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(G1338gat));
  NOR3_X1   g458(.A1(new_n348), .A2(G106gat), .A3(new_n574), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n634), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT53), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n568), .A2(new_n569), .A3(new_n598), .A4(new_n637), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(G106gat), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n661), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n660), .B(KEYINPUT115), .Z(new_n666));
  AOI22_X1  g465(.A1(new_n634), .A2(new_n666), .B1(new_n663), .B2(G106gat), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n665), .B1(new_n662), .B2(new_n667), .ZN(G1339gat));
  INV_X1    g467(.A(KEYINPUT55), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n523), .A2(new_n516), .A3(new_n524), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT54), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n670), .A2(new_n525), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n523), .A2(new_n524), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n673), .A2(new_n671), .A3(new_n515), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n513), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n669), .B1(new_n672), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n515), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n523), .A2(new_n516), .A3(new_n524), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n677), .A2(KEYINPUT54), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n513), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n680), .B1(new_n525), .B2(new_n671), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n679), .A2(KEYINPUT55), .A3(new_n681), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n676), .A2(new_n532), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n430), .A2(new_n435), .A3(new_n442), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n420), .B1(new_n418), .B2(new_n422), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n426), .A2(new_n427), .A3(new_n425), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n441), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n683), .A2(new_n492), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT116), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n676), .A2(new_n448), .A3(new_n532), .A4(new_n682), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n533), .A2(new_n688), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n608), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n509), .B1(new_n690), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n609), .A2(new_n533), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n697), .A2(new_n377), .A3(new_n598), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n536), .A2(new_n284), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n576), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT117), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n702), .B2(new_n232), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT117), .B(G113gat), .Z(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(new_n701), .B2(new_n704), .ZN(G1340gat));
  OAI21_X1  g504(.A(G120gat), .B1(new_n700), .B2(new_n574), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n533), .A2(new_n233), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n706), .B1(new_n700), .B2(new_n707), .ZN(G1341gat));
  NOR2_X1   g507(.A1(new_n700), .A2(new_n510), .ZN(new_n709));
  INV_X1    g508(.A(G127gat), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT118), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n709), .B(new_n711), .Z(G1342gat));
  NOR2_X1   g511(.A1(new_n700), .A2(new_n608), .ZN(new_n713));
  INV_X1    g512(.A(G134gat), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n715), .B1(KEYINPUT56), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(KEYINPUT56), .B2(new_n716), .ZN(G1343gat));
  NOR2_X1   g517(.A1(new_n697), .A2(new_n348), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT57), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n383), .A2(new_n699), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT119), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n533), .A2(new_n724), .A3(new_n688), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n691), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n724), .B1(new_n533), .B2(new_n688), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n608), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT120), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n690), .A2(new_n729), .ZN(new_n730));
  OR2_X1    g529(.A1(new_n728), .A2(KEYINPUT120), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n509), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n598), .B1(new_n732), .B2(new_n696), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n723), .B1(KEYINPUT57), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n734), .A2(new_n448), .ZN(new_n735));
  INV_X1    g534(.A(G141gat), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n722), .A2(new_n719), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n448), .A2(new_n736), .ZN(new_n738));
  OAI22_X1  g537(.A1(new_n735), .A2(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1344gat));
  INV_X1    g540(.A(new_n737), .ZN(new_n742));
  INV_X1    g541(.A(G148gat), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n742), .A2(new_n743), .A3(new_n533), .ZN(new_n744));
  AOI211_X1 g543(.A(KEYINPUT59), .B(new_n743), .C1(new_n734), .C2(new_n533), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT59), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT122), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n509), .B1(new_n728), .B2(new_n689), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(new_n696), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n609), .A2(new_n533), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n692), .A2(KEYINPUT119), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n751), .A2(new_n691), .A3(new_n725), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n492), .A2(new_n688), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n752), .A2(new_n608), .B1(new_n683), .B2(new_n753), .ZN(new_n754));
  OAI211_X1 g553(.A(KEYINPUT122), .B(new_n750), .C1(new_n754), .C2(new_n509), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n749), .A2(new_n598), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(KEYINPUT123), .A3(new_n720), .ZN(new_n757));
  OAI211_X1 g556(.A(KEYINPUT57), .B(new_n598), .C1(new_n695), .C2(new_n696), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT123), .B1(new_n756), .B2(new_n720), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n761), .A2(new_n533), .A3(new_n722), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n746), .B1(new_n762), .B2(G148gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n744), .B1(new_n745), .B2(new_n763), .ZN(G1345gat));
  AOI21_X1  g563(.A(G155gat), .B1(new_n742), .B2(new_n509), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n510), .A2(new_n298), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n765), .B1(new_n734), .B2(new_n766), .ZN(G1346gat));
  NAND3_X1  g566(.A1(new_n742), .A2(new_n297), .A3(new_n492), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n734), .A2(new_n492), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n769), .B2(new_n297), .ZN(G1347gat));
  NAND3_X1  g569(.A1(new_n698), .A2(new_n536), .A3(new_n284), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n576), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(new_n212), .ZN(G1348gat));
  NAND2_X1  g572(.A1(new_n698), .A2(new_n536), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n774), .A2(new_n213), .A3(new_n645), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n771), .A2(new_n559), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n775), .B1(new_n776), .B2(new_n213), .ZN(G1349gat));
  NOR2_X1   g576(.A1(new_n771), .A2(new_n510), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n208), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n217), .B2(new_n778), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT60), .ZN(G1350gat));
  NOR2_X1   g580(.A1(new_n771), .A2(new_n608), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT61), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(new_n784), .A3(G190gat), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n784), .B1(new_n783), .B2(G190gat), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n782), .A2(KEYINPUT124), .A3(new_n209), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT124), .B1(new_n782), .B2(new_n209), .ZN(new_n789));
  OAI22_X1  g588(.A1(new_n786), .A2(new_n787), .B1(new_n788), .B2(new_n789), .ZN(G1351gat));
  NOR3_X1   g589(.A1(new_n551), .A2(new_n540), .A3(new_n348), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n791), .A2(KEYINPUT125), .ZN(new_n792));
  INV_X1    g591(.A(new_n697), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n571), .B1(new_n791), .B2(KEYINPUT125), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(new_n438), .A3(new_n448), .ZN(new_n796));
  AOI211_X1 g595(.A(new_n571), .B(new_n540), .C1(new_n379), .C2(new_n376), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n761), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n448), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n796), .B1(new_n800), .B2(new_n438), .ZN(G1352gat));
  NOR2_X1   g600(.A1(new_n559), .A2(G204gat), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n792), .A2(new_n794), .A3(new_n793), .A4(new_n802), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n803), .B(KEYINPUT62), .Z(new_n804));
  NAND2_X1  g603(.A1(new_n798), .A2(new_n575), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(G204gat), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(G1353gat));
  NOR2_X1   g606(.A1(new_n510), .A2(G211gat), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n795), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n509), .B(new_n797), .C1(new_n759), .C2(new_n760), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G211gat), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT126), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT63), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n810), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n812), .B1(new_n811), .B2(new_n813), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n809), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT127), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI211_X1 g619(.A(KEYINPUT127), .B(new_n809), .C1(new_n816), .C2(new_n817), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(G1354gat));
  AOI21_X1  g621(.A(G218gat), .B1(new_n795), .B2(new_n492), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n492), .A2(G218gat), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n823), .B1(new_n798), .B2(new_n824), .ZN(G1355gat));
endmodule


