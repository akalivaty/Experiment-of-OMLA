//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  INV_X1    g000(.A(G134), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT65), .B1(new_n187), .B2(G137), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT11), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n187), .A2(G137), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT11), .ZN(new_n191));
  OAI211_X1 g005(.A(KEYINPUT65), .B(new_n191), .C1(new_n187), .C2(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT67), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G131), .ZN(new_n196));
  OR2_X1    g010(.A1(new_n193), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n193), .A2(new_n198), .A3(G131), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n195), .A2(new_n197), .A3(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT0), .B(G128), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G143), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n201), .B(KEYINPUT64), .C1(new_n203), .C2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  XNOR2_X1  g021(.A(G143), .B(G146), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n200), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G116), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G119), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  XOR2_X1   g030(.A(KEYINPUT71), .B(G119), .Z(new_n217));
  AOI21_X1  g031(.A(new_n216), .B1(new_n217), .B2(G116), .ZN(new_n218));
  XOR2_X1   g032(.A(KEYINPUT2), .B(G113), .Z(new_n219));
  XNOR2_X1  g033(.A(new_n218), .B(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n202), .B(G146), .C1(new_n222), .C2(KEYINPUT1), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n204), .A3(G143), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n225), .B(KEYINPUT70), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n208), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT69), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n208), .A2(new_n230), .A3(new_n227), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n193), .A2(new_n196), .ZN(new_n234));
  OR3_X1    g048(.A1(new_n187), .A2(KEYINPUT68), .A3(G137), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n190), .A2(KEYINPUT68), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n187), .A2(G137), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n235), .B(G131), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n233), .A2(new_n240), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n213), .A2(new_n221), .A3(new_n241), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n193), .A2(new_n198), .A3(G131), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n198), .B1(new_n193), .B2(G131), .ZN(new_n244));
  NOR3_X1   g058(.A1(new_n243), .A2(new_n244), .A3(new_n234), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n241), .B1(new_n245), .B2(new_n211), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT30), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT30), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n213), .A2(new_n248), .A3(new_n241), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n242), .B1(new_n250), .B2(new_n220), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n252), .B(G101), .ZN(new_n253));
  NOR2_X1   g067(.A1(G237), .A2(G953), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G210), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n253), .B(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT74), .B1(new_n251), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT74), .ZN(new_n258));
  INV_X1    g072(.A(new_n256), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n221), .B1(new_n247), .B2(new_n249), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n258), .B(new_n259), .C1(new_n260), .C2(new_n242), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n221), .B1(new_n213), .B2(new_n241), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT28), .B1(new_n242), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n213), .A2(new_n221), .A3(new_n241), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n263), .A2(new_n266), .A3(new_n256), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT73), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n257), .A2(new_n261), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT75), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT29), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n267), .A2(KEYINPUT73), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n269), .A2(new_n270), .A3(new_n271), .A4(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n266), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n275), .B1(new_n263), .B2(KEYINPUT76), .ZN(new_n276));
  INV_X1    g090(.A(new_n262), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n264), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT76), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(new_n279), .A3(KEYINPUT28), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(new_n271), .ZN(new_n282));
  AOI21_X1  g096(.A(G902), .B1(new_n282), .B2(new_n256), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n257), .A2(new_n268), .A3(new_n271), .A4(new_n261), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT75), .B1(new_n284), .B2(new_n272), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n274), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G472), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT32), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n213), .A2(new_n248), .A3(new_n241), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n248), .B1(new_n213), .B2(new_n241), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n220), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(new_n264), .A3(new_n256), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT31), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n291), .A2(KEYINPUT31), .A3(new_n264), .A4(new_n256), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n263), .A2(new_n266), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n259), .ZN(new_n298));
  AOI21_X1  g112(.A(G902), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G472), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT72), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n294), .A2(new_n295), .B1(new_n297), .B2(new_n259), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n303));
  NOR4_X1   g117(.A1(new_n302), .A2(new_n303), .A3(G472), .A4(G902), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n288), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n299), .A2(KEYINPUT32), .A3(new_n300), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n287), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G902), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n214), .A2(G122), .ZN(new_n309));
  INV_X1    g123(.A(G122), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(G116), .ZN(new_n311));
  OAI21_X1  g125(.A(G107), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(G116), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n214), .A2(G122), .ZN(new_n314));
  INV_X1    g128(.A(G107), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n222), .A2(G143), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n202), .A2(G128), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n319), .A3(KEYINPUT13), .ZN(new_n320));
  OR3_X1    g134(.A1(new_n222), .A2(KEYINPUT13), .A3(G143), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G134), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n318), .A2(new_n319), .A3(new_n187), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT89), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT89), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n318), .A2(new_n319), .A3(new_n325), .A4(new_n187), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n317), .A2(new_n322), .A3(new_n324), .A4(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n318), .A2(new_n319), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G134), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n323), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n311), .A2(KEYINPUT14), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n313), .A2(new_n314), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n331), .B(G107), .C1(new_n332), .C2(KEYINPUT14), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n333), .A3(new_n316), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT9), .B(G234), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT80), .ZN(new_n336));
  INV_X1    g150(.A(G953), .ZN(new_n337));
  OR2_X1    g151(.A1(KEYINPUT9), .A2(G234), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n339));
  NAND2_X1  g153(.A1(KEYINPUT9), .A2(G234), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AND4_X1   g155(.A1(G217), .A2(new_n336), .A3(new_n337), .A4(new_n341), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n327), .A2(new_n334), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n342), .B1(new_n327), .B2(new_n334), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n308), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G478), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n346), .B1(KEYINPUT15), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT15), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n345), .A2(new_n349), .A3(G478), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n352), .A2(KEYINPUT90), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(KEYINPUT90), .ZN(new_n354));
  OR2_X1    g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G475), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n254), .A2(G214), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(KEYINPUT87), .A3(G143), .ZN(new_n358));
  OR2_X1    g172(.A1(KEYINPUT87), .A2(G143), .ZN(new_n359));
  NAND2_X1  g173(.A1(KEYINPUT87), .A2(G143), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n359), .A2(G214), .A3(new_n254), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(KEYINPUT18), .A2(G131), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(G125), .B(G140), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n365), .B(new_n204), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n358), .A2(new_n361), .A3(KEYINPUT18), .A4(G131), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n364), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT88), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT88), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n364), .A2(new_n366), .A3(new_n370), .A4(new_n367), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(G113), .B(G122), .ZN(new_n373));
  INV_X1    g187(.A(G104), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n373), .B(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n196), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n362), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT17), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n358), .A2(new_n361), .A3(new_n196), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G125), .ZN(new_n381));
  NOR3_X1   g195(.A1(new_n381), .A2(KEYINPUT16), .A3(G140), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n382), .B1(new_n365), .B2(KEYINPUT16), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n383), .B(new_n204), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n380), .B(new_n384), .C1(new_n378), .C2(new_n379), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n372), .A2(new_n375), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n377), .A2(new_n379), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n383), .A2(G146), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT19), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n365), .B(new_n390), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n388), .B(new_n389), .C1(G146), .C2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n375), .B1(new_n372), .B2(new_n392), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n356), .B(new_n308), .C1(new_n387), .C2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT20), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n372), .A2(new_n392), .ZN(new_n397));
  INV_X1    g211(.A(new_n375), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n386), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n400), .A2(KEYINPUT20), .A3(new_n356), .A4(new_n308), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n375), .B1(new_n372), .B2(new_n385), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n308), .B1(new_n387), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G475), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n396), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  OR2_X1    g219(.A1(new_n355), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(G214), .B1(G237), .B2(G902), .ZN(new_n407));
  INV_X1    g221(.A(G952), .ZN(new_n408));
  AOI211_X1 g222(.A(G953), .B(new_n408), .C1(G234), .C2(G237), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  AOI211_X1 g224(.A(new_n308), .B(new_n337), .C1(G234), .C2(G237), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  XOR2_X1   g226(.A(KEYINPUT21), .B(G898), .Z(new_n413));
  OAI21_X1  g227(.A(new_n410), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT84), .ZN(new_n415));
  XNOR2_X1  g229(.A(KEYINPUT71), .B(G119), .ZN(new_n416));
  OAI211_X1 g230(.A(KEYINPUT5), .B(new_n215), .C1(new_n416), .C2(new_n214), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n217), .A2(G116), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n417), .B(G113), .C1(new_n418), .C2(KEYINPUT5), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n218), .A2(new_n219), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n374), .A2(G107), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n315), .A2(G104), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G101), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT3), .B1(new_n374), .B2(G107), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT3), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n315), .A3(G104), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(new_n428), .A3(new_n422), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT81), .B(G101), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n425), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n415), .B1(new_n421), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n431), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n419), .A2(new_n433), .A3(KEYINPUT84), .A4(new_n420), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n429), .A2(G101), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n436), .A2(KEYINPUT4), .ZN(new_n437));
  XOR2_X1   g251(.A(KEYINPUT81), .B(G101), .Z(new_n438));
  NAND4_X1  g252(.A1(new_n438), .A2(new_n422), .A3(new_n428), .A4(new_n426), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(new_n436), .A3(KEYINPUT4), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT82), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n439), .A2(new_n436), .A3(KEYINPUT82), .A4(KEYINPUT4), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n220), .A2(new_n437), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n435), .A2(new_n444), .ZN(new_n445));
  XOR2_X1   g259(.A(G110), .B(G122), .Z(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n446), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n435), .A2(new_n448), .A3(new_n444), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(KEYINPUT6), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT6), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n445), .A2(new_n451), .A3(new_n446), .ZN(new_n452));
  AOI21_X1  g266(.A(G125), .B1(new_n226), .B2(new_n232), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT85), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n211), .A2(new_n381), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n337), .A2(G224), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT85), .B1(new_n453), .B2(new_n456), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n460), .B1(new_n458), .B2(new_n461), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n450), .A2(new_n452), .A3(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n453), .A2(new_n456), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n459), .A2(KEYINPUT7), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n466), .B(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT86), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n421), .B1(new_n469), .B2(new_n433), .ZN(new_n470));
  AOI211_X1 g284(.A(KEYINPUT86), .B(new_n431), .C1(new_n419), .C2(new_n420), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n446), .B(KEYINPUT8), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(G902), .B1(new_n474), .B2(new_n449), .ZN(new_n475));
  OAI21_X1  g289(.A(G210), .B1(G237), .B2(G902), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n465), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n476), .B1(new_n465), .B2(new_n475), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n407), .B(new_n414), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n406), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G221), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n336), .A2(new_n341), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n482), .B1(new_n483), .B2(new_n308), .ZN(new_n484));
  XNOR2_X1  g298(.A(G110), .B(G140), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n337), .A2(G227), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n485), .B(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT70), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n225), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n225), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT70), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n232), .A2(new_n431), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n208), .A2(new_n230), .A3(new_n227), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n230), .B1(new_n208), .B2(new_n227), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n433), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(KEYINPUT12), .A3(new_n200), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT83), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n200), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT12), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT83), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n497), .A2(new_n503), .A3(KEYINPUT12), .A4(new_n200), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n499), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n442), .A2(new_n212), .A3(new_n437), .A4(new_n443), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n233), .A2(KEYINPUT10), .A3(new_n433), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT10), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n496), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n506), .A2(new_n507), .A3(new_n245), .A4(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n487), .B1(new_n505), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n510), .A2(new_n487), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n506), .A2(new_n507), .A3(new_n509), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n200), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G469), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n511), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n516), .A2(new_n308), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n505), .A2(new_n512), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n514), .A2(new_n510), .ZN(new_n521));
  INV_X1    g335(.A(new_n487), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(G902), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n519), .B1(new_n524), .B2(new_n516), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n484), .B1(new_n518), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n337), .A2(G221), .A3(G234), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT22), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(G137), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G119), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n531), .A2(KEYINPUT71), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n531), .A2(KEYINPUT71), .ZN(new_n533));
  OAI21_X1  g347(.A(G128), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT24), .B(G110), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n531), .A2(G128), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n534), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT77), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT78), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT23), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n543), .B1(new_n534), .B2(new_n538), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT23), .B1(new_n416), .B2(new_n222), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n545), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n537), .B1(new_n217), .B2(G128), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n547), .B(KEYINPUT78), .C1(new_n548), .C2(new_n543), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n546), .A2(new_n549), .A3(G110), .ZN(new_n550));
  INV_X1    g364(.A(new_n384), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n541), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT79), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n547), .B1(new_n548), .B2(new_n543), .ZN(new_n554));
  OAI22_X1  g368(.A1(new_n554), .A2(G110), .B1(new_n536), .B2(new_n548), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n365), .A2(new_n204), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n556), .A3(new_n389), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n552), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n553), .B1(new_n552), .B2(new_n557), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n530), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n552), .A2(new_n557), .A3(new_n529), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(new_n308), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT25), .ZN(new_n563));
  INV_X1    g377(.A(G217), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n564), .B1(G234), .B2(new_n308), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT25), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n560), .A2(new_n566), .A3(new_n308), .A4(new_n561), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n563), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n565), .A2(G902), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n560), .A2(new_n561), .A3(new_n569), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n307), .A2(new_n481), .A3(new_n526), .A4(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(new_n430), .ZN(G3));
  NOR2_X1   g387(.A1(new_n299), .A2(new_n300), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT31), .B1(new_n251), .B2(new_n256), .ZN(new_n575));
  NOR4_X1   g389(.A1(new_n260), .A2(new_n293), .A3(new_n242), .A4(new_n259), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n298), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(new_n300), .A3(new_n308), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n303), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n299), .A2(KEYINPUT72), .A3(new_n300), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n574), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n581), .A2(new_n526), .A3(new_n571), .ZN(new_n582));
  INV_X1    g396(.A(new_n407), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n478), .B2(KEYINPUT91), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n465), .A2(new_n475), .ZN(new_n585));
  INV_X1    g399(.A(new_n476), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT91), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(new_n588), .A3(new_n477), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n414), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT92), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n592), .B1(new_n343), .B2(new_n344), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT33), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n592), .B(KEYINPUT33), .C1(new_n343), .C2(new_n344), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  OAI211_X1 g411(.A(G478), .B(new_n308), .C1(new_n595), .C2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n346), .A2(G478), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n405), .A2(new_n601), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n590), .A2(new_n591), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n582), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT34), .B(G104), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G6));
  AND3_X1   g420(.A1(new_n396), .A2(new_n401), .A3(new_n404), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n355), .A2(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n590), .A2(new_n591), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n582), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT35), .B(G107), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G9));
  NOR2_X1   g426(.A1(new_n558), .A2(new_n559), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n530), .A2(KEYINPUT36), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n613), .B(new_n614), .Z(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n569), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n568), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n617), .A2(new_n526), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n581), .A2(new_n481), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G110), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT93), .B(KEYINPUT37), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G12));
  INV_X1    g436(.A(new_n590), .ZN(new_n623));
  INV_X1    g437(.A(G900), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n409), .B1(new_n411), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n608), .A2(new_n625), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n623), .A2(new_n618), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n307), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G128), .ZN(G30));
  NOR2_X1   g443(.A1(new_n251), .A2(new_n259), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n308), .B1(new_n278), .B2(new_n256), .ZN(new_n631));
  OAI21_X1  g445(.A(G472), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n305), .A2(new_n306), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(new_n625), .B(KEYINPUT39), .Z(new_n634));
  NAND2_X1  g448(.A1(new_n526), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(KEYINPUT40), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n617), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n355), .A2(new_n405), .ZN(new_n638));
  AOI211_X1 g452(.A(new_n583), .B(new_n638), .C1(new_n635), .C2(KEYINPUT40), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT38), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n640), .B1(new_n478), .B2(new_n479), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n587), .A2(KEYINPUT38), .A3(new_n477), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n633), .A2(new_n637), .A3(new_n639), .A4(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G143), .ZN(G45));
  AOI21_X1  g459(.A(new_n590), .B1(new_n568), .B2(new_n616), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n602), .A2(new_n625), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n526), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n307), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G146), .ZN(G48));
  XNOR2_X1  g464(.A(new_n524), .B(G469), .ZN(new_n651));
  INV_X1    g465(.A(new_n484), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n307), .A2(new_n603), .A3(new_n571), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT41), .B(G113), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G15));
  NAND4_X1  g471(.A1(new_n307), .A2(new_n571), .A3(new_n609), .A4(new_n654), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G116), .ZN(G18));
  INV_X1    g473(.A(new_n406), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n653), .A2(new_n591), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n307), .A2(new_n646), .A3(new_n660), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G119), .ZN(G21));
  AOI22_X1  g477(.A1(new_n259), .A2(new_n281), .B1(new_n294), .B2(new_n295), .ZN(new_n664));
  NOR2_X1   g478(.A1(G472), .A2(G902), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(KEYINPUT94), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT94), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n575), .A2(new_n576), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n256), .B1(new_n276), .B2(new_n280), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n668), .B(new_n665), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT95), .B(G472), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n672), .B1(new_n302), .B2(G902), .ZN(new_n673));
  AND4_X1   g487(.A1(new_n571), .A2(new_n667), .A3(new_n671), .A4(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n590), .A2(new_n638), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n674), .A2(new_n675), .A3(new_n661), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G122), .ZN(G24));
  NAND4_X1  g491(.A1(new_n667), .A2(new_n617), .A3(new_n671), .A4(new_n673), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n584), .A2(new_n589), .A3(new_n647), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n678), .A2(new_n679), .A3(new_n653), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n381), .ZN(G27));
  NAND3_X1  g495(.A1(new_n587), .A2(new_n477), .A3(new_n407), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT97), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n587), .A2(KEYINPUT97), .A3(new_n477), .A4(new_n407), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n684), .A2(new_n647), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT96), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n525), .B1(new_n687), .B2(new_n517), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n517), .A2(new_n687), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n652), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n307), .A2(new_n571), .A3(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n571), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n578), .B(KEYINPUT32), .ZN(new_n697));
  AOI211_X1 g511(.A(new_n694), .B(new_n696), .C1(new_n287), .C2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n692), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G131), .ZN(G33));
  NAND2_X1  g515(.A1(new_n684), .A2(new_n685), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n702), .A2(new_n608), .A3(new_n625), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n524), .A2(new_n516), .ZN(new_n704));
  INV_X1    g518(.A(new_n519), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n505), .A2(new_n510), .ZN(new_n707));
  AOI22_X1  g521(.A1(new_n707), .A2(new_n522), .B1(new_n512), .B2(new_n514), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n687), .B1(new_n708), .B2(G469), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n484), .B1(new_n710), .B2(new_n689), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n307), .A2(new_n703), .A3(new_n571), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G134), .ZN(G36));
  INV_X1    g527(.A(new_n581), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT99), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n593), .A2(new_n594), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n347), .B(G902), .C1(new_n717), .C2(new_n596), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n716), .B1(new_n718), .B2(new_n599), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n598), .A2(KEYINPUT99), .A3(new_n600), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n715), .B1(new_n721), .B2(new_n405), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT100), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI211_X1 g538(.A(KEYINPUT100), .B(new_n715), .C1(new_n721), .C2(new_n405), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n607), .A2(KEYINPUT43), .A3(new_n601), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n714), .A2(new_n617), .A3(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n708), .A2(KEYINPUT45), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n733), .B1(new_n511), .B2(new_n515), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n732), .A2(G469), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n705), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT46), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n736), .A2(new_n737), .B1(new_n516), .B2(new_n524), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n735), .A2(KEYINPUT46), .A3(new_n705), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n652), .A3(new_n634), .ZN(new_n741));
  XOR2_X1   g555(.A(new_n741), .B(KEYINPUT98), .Z(new_n742));
  OR2_X1    g556(.A1(new_n729), .A2(new_n730), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT101), .ZN(new_n744));
  INV_X1    g558(.A(new_n702), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n744), .B1(new_n743), .B2(new_n745), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n731), .B(new_n742), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G137), .ZN(G39));
  NOR3_X1   g563(.A1(new_n307), .A2(new_n571), .A3(new_n686), .ZN(new_n750));
  XOR2_X1   g564(.A(new_n750), .B(KEYINPUT102), .Z(new_n751));
  AOI21_X1  g565(.A(KEYINPUT47), .B1(new_n740), .B2(new_n652), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT47), .ZN(new_n753));
  AOI211_X1 g567(.A(new_n753), .B(new_n484), .C1(new_n738), .C2(new_n739), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n751), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G140), .ZN(G42));
  INV_X1    g570(.A(new_n602), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n757), .B1(new_n351), .B2(new_n607), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n480), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n581), .A2(new_n759), .A3(new_n526), .A4(new_n571), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n760), .A2(new_n619), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n572), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT103), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n761), .A2(new_n572), .A3(KEYINPUT103), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n655), .A2(new_n658), .A3(new_n662), .A4(new_n676), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n694), .A2(new_n693), .B1(new_n698), .B2(new_n692), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n711), .A2(new_n647), .A3(new_n684), .A4(new_n685), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT104), .B1(new_n770), .B2(new_n678), .ZN(new_n771));
  INV_X1    g585(.A(new_n686), .ZN(new_n772));
  INV_X1    g586(.A(new_n678), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT104), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n772), .A2(new_n773), .A3(new_n774), .A4(new_n711), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n702), .A2(new_n351), .A3(new_n405), .ZN(new_n777));
  INV_X1    g591(.A(new_n625), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n307), .A2(new_n777), .A3(new_n618), .A4(new_n778), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n776), .A2(new_n779), .A3(new_n712), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n766), .A2(new_n769), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT105), .B1(new_n617), .B2(new_n625), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT105), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n616), .A2(new_n784), .A3(new_n568), .A4(new_n778), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n691), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n633), .A2(new_n675), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n680), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n649), .A2(new_n628), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n789), .A2(KEYINPUT106), .A3(KEYINPUT52), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(new_n789), .B2(KEYINPUT106), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n781), .A2(new_n782), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n766), .A2(new_n769), .A3(new_n780), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n789), .A2(KEYINPUT107), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n680), .B1(new_n307), .B2(new_n627), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT107), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n796), .A2(new_n797), .A3(new_n649), .A4(new_n787), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n795), .A2(KEYINPUT52), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT52), .B1(new_n795), .B2(new_n798), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n794), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n793), .B(KEYINPUT54), .C1(new_n801), .C2(new_n782), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n803));
  INV_X1    g617(.A(new_n765), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT103), .B1(new_n761), .B2(new_n572), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n780), .B(KEYINPUT53), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT108), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n808), .B1(new_n767), .B2(new_n768), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n658), .A2(new_n662), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n655), .A2(new_n676), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n700), .A2(new_n810), .A3(new_n811), .A4(KEYINPUT108), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n807), .A2(new_n792), .A3(new_n809), .A4(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n803), .B(new_n813), .C1(new_n801), .C2(KEYINPUT53), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n802), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT109), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n802), .A2(new_n814), .A3(KEYINPUT109), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n410), .B1(new_n726), .B2(new_n727), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(new_n623), .A3(new_n674), .A4(new_n654), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n745), .A2(new_n654), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n571), .A2(new_n409), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n821), .A2(new_n633), .A3(new_n822), .ZN(new_n823));
  AOI211_X1 g637(.A(new_n408), .B(G953), .C1(new_n823), .C2(new_n757), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n821), .A2(new_n633), .A3(new_n405), .A4(new_n822), .ZN(new_n825));
  INV_X1    g639(.A(new_n601), .ZN(new_n826));
  INV_X1    g640(.A(new_n819), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n821), .A2(new_n827), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n825), .A2(new_n826), .B1(new_n773), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT110), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n830), .B1(new_n752), .B2(new_n754), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n736), .A2(new_n737), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n832), .A2(new_n704), .A3(new_n739), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n753), .B1(new_n833), .B2(new_n484), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n740), .A2(KEYINPUT47), .A3(new_n652), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(KEYINPUT110), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n651), .A2(new_n484), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n831), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n819), .A2(new_n745), .A3(new_n674), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n407), .B1(new_n641), .B2(new_n642), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n819), .A2(new_n654), .A3(new_n674), .A4(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT111), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(KEYINPUT50), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n843), .A2(KEYINPUT50), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n844), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n846), .A2(new_n848), .A3(KEYINPUT112), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT112), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n842), .A2(new_n847), .ZN(new_n851));
  INV_X1    g665(.A(new_n844), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n850), .B1(new_n853), .B2(new_n845), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n829), .B(new_n840), .C1(new_n849), .C2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT113), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n856), .B1(new_n855), .B2(new_n857), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n820), .B(new_n824), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n696), .B1(new_n287), .B2(new_n697), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n828), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n862), .B(KEYINPUT48), .Z(new_n863));
  AND3_X1   g677(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n864), .A2(KEYINPUT114), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(KEYINPUT114), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n865), .A2(new_n839), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n853), .A2(new_n845), .ZN(new_n868));
  AND4_X1   g682(.A1(KEYINPUT51), .A2(new_n867), .A3(new_n868), .A4(new_n829), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n860), .A2(new_n863), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n817), .A2(new_n818), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT115), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n408), .A2(new_n337), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n817), .A2(new_n870), .A3(KEYINPUT115), .A4(new_n818), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n651), .B(KEYINPUT49), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(new_n652), .A3(new_n601), .ZN(new_n878));
  NOR4_X1   g692(.A1(new_n878), .A2(new_n583), .A3(new_n696), .A4(new_n643), .ZN(new_n879));
  INV_X1    g693(.A(new_n633), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n607), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n876), .A2(new_n881), .ZN(G75));
  NOR2_X1   g696(.A1(new_n337), .A2(G952), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n799), .A2(new_n800), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT53), .B1(new_n884), .B2(new_n781), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n809), .A2(new_n812), .ZN(new_n886));
  NOR4_X1   g700(.A1(new_n886), .A2(new_n806), .A3(new_n791), .A4(new_n790), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(new_n308), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(G210), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT56), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n450), .A2(new_n452), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(new_n464), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT55), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n883), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n890), .A2(KEYINPUT116), .ZN(new_n897));
  XNOR2_X1  g711(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT116), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n889), .A2(new_n900), .A3(G210), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n897), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n896), .A2(new_n902), .ZN(G51));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n888), .A2(new_n308), .A3(new_n735), .ZN(new_n905));
  XOR2_X1   g719(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n519), .ZN(new_n907));
  INV_X1    g721(.A(new_n906), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n705), .ZN(new_n909));
  INV_X1    g723(.A(new_n814), .ZN(new_n910));
  INV_X1    g724(.A(new_n800), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n795), .A2(KEYINPUT52), .A3(new_n798), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n782), .B1(new_n913), .B2(new_n794), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n803), .B1(new_n914), .B2(new_n813), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n907), .B(new_n909), .C1(new_n910), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n520), .A2(new_n523), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n905), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n904), .B1(new_n918), .B2(new_n883), .ZN(new_n919));
  INV_X1    g733(.A(new_n883), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT54), .B1(new_n885), .B2(new_n887), .ZN(new_n921));
  AOI22_X1  g735(.A1(new_n921), .A2(new_n814), .B1(new_n705), .B2(new_n908), .ZN(new_n922));
  AOI22_X1  g736(.A1(new_n922), .A2(new_n907), .B1(new_n523), .B2(new_n520), .ZN(new_n923));
  OAI211_X1 g737(.A(KEYINPUT119), .B(new_n920), .C1(new_n923), .C2(new_n905), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n919), .A2(new_n924), .ZN(G54));
  NAND3_X1  g739(.A1(new_n889), .A2(KEYINPUT58), .A3(G475), .ZN(new_n926));
  INV_X1    g740(.A(new_n400), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n928), .A2(new_n929), .A3(new_n883), .ZN(G60));
  NOR2_X1   g744(.A1(new_n595), .A2(new_n597), .ZN(new_n931));
  XNOR2_X1  g745(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n347), .A2(new_n308), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n932), .B(new_n933), .Z(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  AOI211_X1 g749(.A(new_n931), .B(new_n935), .C1(new_n921), .C2(new_n814), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n817), .A2(new_n818), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n934), .ZN(new_n938));
  AOI211_X1 g752(.A(new_n883), .B(new_n936), .C1(new_n938), .C2(new_n931), .ZN(G63));
  NAND2_X1  g753(.A1(new_n914), .A2(new_n813), .ZN(new_n940));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT60), .Z(new_n942));
  XNOR2_X1  g756(.A(new_n615), .B(KEYINPUT121), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n944), .A2(KEYINPUT122), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n940), .A2(new_n942), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n560), .A2(new_n561), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n883), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n944), .A2(KEYINPUT122), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n945), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n945), .A2(KEYINPUT61), .A3(new_n948), .A4(new_n949), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(G66));
  AOI21_X1  g768(.A(new_n337), .B1(new_n413), .B2(G224), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n766), .A2(new_n811), .A3(new_n810), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n955), .B1(new_n956), .B2(new_n337), .ZN(new_n957));
  INV_X1    g771(.A(G898), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n893), .B1(new_n958), .B2(G953), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n957), .B(new_n959), .ZN(G69));
  NAND2_X1  g774(.A1(new_n796), .A2(new_n649), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT123), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n644), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT62), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n755), .A2(new_n748), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n307), .A2(new_n571), .ZN(new_n968));
  NOR4_X1   g782(.A1(new_n968), .A2(new_n635), .A3(new_n702), .A4(new_n758), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n966), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n337), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n250), .B(new_n391), .Z(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n742), .A2(new_n675), .A3(new_n861), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n963), .A2(new_n700), .A3(new_n712), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n967), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n974), .B1(new_n979), .B2(new_n337), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n624), .B2(new_n337), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n337), .B1(G227), .B2(G900), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT124), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n983), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n982), .B(new_n985), .ZN(G72));
  NAND2_X1  g800(.A1(G472), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT63), .Z(new_n988));
  OAI21_X1  g802(.A(new_n988), .B1(new_n971), .B2(new_n956), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT125), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI211_X1 g805(.A(KEYINPUT125), .B(new_n988), .C1(new_n971), .C2(new_n956), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n991), .A2(new_n630), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n257), .A2(new_n292), .A3(new_n261), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n988), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT127), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n793), .B(new_n996), .C1(new_n801), .C2(new_n782), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT126), .ZN(new_n998));
  NOR4_X1   g812(.A1(new_n967), .A2(new_n978), .A3(new_n956), .A4(new_n977), .ZN(new_n999));
  INV_X1    g813(.A(new_n988), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n259), .B(new_n251), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n998), .B1(new_n1001), .B2(new_n920), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n1001), .A2(new_n998), .A3(new_n920), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n993), .B(new_n997), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(G57));
endmodule


