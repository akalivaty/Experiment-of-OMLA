

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U558 ( .A1(G651), .A2(n587), .ZN(n798) );
  NOR2_X2 U559 ( .A1(n523), .A2(G2105), .ZN(n524) );
  NOR2_X1 U560 ( .A1(n971), .A2(n627), .ZN(n629) );
  XNOR2_X1 U561 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U562 ( .A1(n691), .A2(n690), .ZN(n738) );
  BUF_X1 U563 ( .A(n622), .Z(n680) );
  OR2_X1 U564 ( .A1(n738), .A2(n693), .ZN(n694) );
  NAND2_X1 U565 ( .A1(n620), .A2(n619), .ZN(n971) );
  BUF_X1 U566 ( .A(n630), .Z(n544) );
  BUF_X1 U567 ( .A(n705), .Z(n706) );
  INV_X4 U568 ( .A(G2104), .ZN(n523) );
  OR2_X2 U569 ( .A1(n587), .A2(n549), .ZN(n550) );
  XNOR2_X2 U570 ( .A(n541), .B(KEYINPUT84), .ZN(G164) );
  XNOR2_X1 U571 ( .A(n612), .B(n611), .ZN(n613) );
  XNOR2_X1 U572 ( .A(KEYINPUT67), .B(KEYINPUT23), .ZN(n525) );
  INV_X1 U573 ( .A(KEYINPUT26), .ZN(n623) );
  INV_X1 U574 ( .A(KEYINPUT64), .ZN(n628) );
  INV_X1 U575 ( .A(KEYINPUT93), .ZN(n645) );
  NAND2_X1 U576 ( .A1(n665), .A2(n664), .ZN(n667) );
  XNOR2_X1 U577 ( .A(n667), .B(n666), .ZN(n670) );
  INV_X1 U578 ( .A(KEYINPUT96), .ZN(n673) );
  INV_X1 U579 ( .A(KEYINPUT32), .ZN(n688) );
  NAND2_X1 U580 ( .A1(n593), .A2(n703), .ZN(n622) );
  XNOR2_X1 U581 ( .A(KEYINPUT74), .B(KEYINPUT12), .ZN(n611) );
  NOR2_X1 U582 ( .A1(G543), .A2(n549), .ZN(n542) );
  XNOR2_X1 U583 ( .A(n638), .B(KEYINPUT15), .ZN(n919) );
  XNOR2_X1 U584 ( .A(n526), .B(n525), .ZN(n528) );
  NOR2_X2 U585 ( .A1(n534), .A2(n533), .ZN(G160) );
  XNOR2_X1 U586 ( .A(n524), .B(KEYINPUT66), .ZN(n705) );
  NAND2_X1 U587 ( .A1(n705), .A2(G101), .ZN(n526) );
  AND2_X1 U588 ( .A1(G2104), .A2(G2105), .ZN(n899) );
  NAND2_X1 U589 ( .A1(G113), .A2(n899), .ZN(n527) );
  NAND2_X1 U590 ( .A1(n528), .A2(n527), .ZN(n534) );
  NOR2_X1 U591 ( .A1(G2104), .A2(G2105), .ZN(n529) );
  XOR2_X1 U592 ( .A(KEYINPUT17), .B(n529), .Z(n704) );
  NAND2_X1 U593 ( .A1(G137), .A2(n704), .ZN(n532) );
  NAND2_X1 U594 ( .A1(n523), .A2(G2105), .ZN(n530) );
  XNOR2_X2 U595 ( .A(n530), .B(KEYINPUT65), .ZN(n902) );
  NAND2_X1 U596 ( .A1(G125), .A2(n902), .ZN(n531) );
  NAND2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U598 ( .A1(G138), .A2(n704), .ZN(n536) );
  NAND2_X1 U599 ( .A1(G102), .A2(n705), .ZN(n535) );
  NAND2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n540) );
  NAND2_X1 U601 ( .A1(G114), .A2(n899), .ZN(n538) );
  NAND2_X1 U602 ( .A1(G126), .A2(n902), .ZN(n537) );
  NAND2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U604 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U605 ( .A(KEYINPUT0), .B(G543), .Z(n587) );
  NAND2_X1 U606 ( .A1(n798), .A2(G51), .ZN(n546) );
  XOR2_X1 U607 ( .A(G651), .B(KEYINPUT68), .Z(n549) );
  XOR2_X1 U608 ( .A(KEYINPUT1), .B(n542), .Z(n543) );
  XNOR2_X1 U609 ( .A(KEYINPUT70), .B(n543), .ZN(n630) );
  NAND2_X1 U610 ( .A1(G63), .A2(n544), .ZN(n545) );
  NAND2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U612 ( .A(KEYINPUT6), .B(n547), .ZN(n556) );
  NOR2_X2 U613 ( .A1(G651), .A2(G543), .ZN(n795) );
  NAND2_X1 U614 ( .A1(n795), .A2(G89), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n548), .B(KEYINPUT4), .ZN(n552) );
  XNOR2_X2 U616 ( .A(n550), .B(KEYINPUT69), .ZN(n802) );
  NAND2_X1 U617 ( .A1(G76), .A2(n802), .ZN(n551) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(KEYINPUT5), .B(n553), .ZN(n554) );
  XNOR2_X1 U620 ( .A(KEYINPUT77), .B(n554), .ZN(n555) );
  NOR2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U622 ( .A(KEYINPUT7), .B(n557), .Z(G168) );
  NAND2_X1 U623 ( .A1(n798), .A2(G52), .ZN(n559) );
  NAND2_X1 U624 ( .A1(G64), .A2(n544), .ZN(n558) );
  NAND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(KEYINPUT72), .B(n560), .ZN(n565) );
  NAND2_X1 U627 ( .A1(G90), .A2(n795), .ZN(n562) );
  NAND2_X1 U628 ( .A1(G77), .A2(n802), .ZN(n561) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U630 ( .A(KEYINPUT9), .B(n563), .Z(n564) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(G171) );
  INV_X1 U632 ( .A(G171), .ZN(G301) );
  XOR2_X1 U633 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U634 ( .A1(G88), .A2(n795), .ZN(n567) );
  NAND2_X1 U635 ( .A1(G75), .A2(n802), .ZN(n566) );
  NAND2_X1 U636 ( .A1(n567), .A2(n566), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n798), .A2(G50), .ZN(n569) );
  NAND2_X1 U638 ( .A1(G62), .A2(n544), .ZN(n568) );
  NAND2_X1 U639 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U640 ( .A1(n571), .A2(n570), .ZN(G166) );
  INV_X1 U641 ( .A(G166), .ZN(G303) );
  NAND2_X1 U642 ( .A1(G86), .A2(n795), .ZN(n573) );
  NAND2_X1 U643 ( .A1(G48), .A2(n798), .ZN(n572) );
  NAND2_X1 U644 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U645 ( .A1(n802), .A2(G73), .ZN(n574) );
  XOR2_X1 U646 ( .A(KEYINPUT2), .B(n574), .Z(n575) );
  NOR2_X1 U647 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U648 ( .A1(G61), .A2(n544), .ZN(n577) );
  NAND2_X1 U649 ( .A1(n578), .A2(n577), .ZN(G305) );
  NAND2_X1 U650 ( .A1(G85), .A2(n795), .ZN(n580) );
  NAND2_X1 U651 ( .A1(G47), .A2(n798), .ZN(n579) );
  NAND2_X1 U652 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U653 ( .A1(G60), .A2(n544), .ZN(n581) );
  XNOR2_X1 U654 ( .A(KEYINPUT71), .B(n581), .ZN(n582) );
  NOR2_X1 U655 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U656 ( .A1(n802), .A2(G72), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n585), .A2(n584), .ZN(G290) );
  NAND2_X1 U658 ( .A1(G49), .A2(n798), .ZN(n586) );
  XNOR2_X1 U659 ( .A(n586), .B(KEYINPUT80), .ZN(n592) );
  NAND2_X1 U660 ( .A1(G87), .A2(n587), .ZN(n589) );
  NAND2_X1 U661 ( .A1(G74), .A2(G651), .ZN(n588) );
  NAND2_X1 U662 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U663 ( .A1(n544), .A2(n590), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n592), .A2(n591), .ZN(G288) );
  NAND2_X1 U665 ( .A1(G160), .A2(G40), .ZN(n702) );
  INV_X1 U666 ( .A(n702), .ZN(n593) );
  NOR2_X2 U667 ( .A1(G164), .A2(G1384), .ZN(n703) );
  NAND2_X1 U668 ( .A1(G8), .A2(n680), .ZN(n743) );
  NOR2_X1 U669 ( .A1(G1966), .A2(n743), .ZN(n678) );
  XNOR2_X1 U670 ( .A(KEYINPUT31), .B(KEYINPUT95), .ZN(n609) );
  NOR2_X1 U671 ( .A1(G2084), .A2(n680), .ZN(n675) );
  NOR2_X1 U672 ( .A1(n678), .A2(n675), .ZN(n594) );
  NAND2_X1 U673 ( .A1(G8), .A2(n594), .ZN(n595) );
  XOR2_X1 U674 ( .A(KEYINPUT30), .B(n595), .Z(n597) );
  INV_X1 U675 ( .A(G168), .ZN(n596) );
  NAND2_X1 U676 ( .A1(n597), .A2(n596), .ZN(n607) );
  INV_X1 U677 ( .A(n680), .ZN(n657) );
  NOR2_X1 U678 ( .A1(n657), .A2(G1961), .ZN(n598) );
  NOR2_X1 U679 ( .A1(KEYINPUT90), .A2(n598), .ZN(n605) );
  XOR2_X1 U680 ( .A(G2078), .B(KEYINPUT25), .Z(n932) );
  NOR2_X1 U681 ( .A1(n680), .A2(n932), .ZN(n599) );
  XNOR2_X1 U682 ( .A(n599), .B(KEYINPUT91), .ZN(n603) );
  INV_X1 U683 ( .A(KEYINPUT90), .ZN(n600) );
  NOR2_X1 U684 ( .A1(G1961), .A2(n600), .ZN(n601) );
  NAND2_X1 U685 ( .A1(n680), .A2(n601), .ZN(n602) );
  NAND2_X1 U686 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U687 ( .A1(n605), .A2(n604), .ZN(n668) );
  NAND2_X1 U688 ( .A1(n668), .A2(G301), .ZN(n606) );
  NAND2_X1 U689 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U690 ( .A(n609), .B(n608), .ZN(n672) );
  NAND2_X1 U691 ( .A1(G56), .A2(n630), .ZN(n610) );
  XNOR2_X1 U692 ( .A(KEYINPUT14), .B(n610), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n802), .A2(G68), .ZN(n614) );
  NAND2_X1 U694 ( .A1(G81), .A2(n795), .ZN(n612) );
  NAND2_X1 U695 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U696 ( .A(n615), .B(KEYINPUT13), .ZN(n616) );
  NAND2_X1 U697 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U698 ( .A(n618), .B(KEYINPUT75), .ZN(n620) );
  NAND2_X1 U699 ( .A1(G43), .A2(n798), .ZN(n619) );
  INV_X1 U700 ( .A(G1996), .ZN(n621) );
  NOR2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n624) );
  XNOR2_X1 U702 ( .A(n624), .B(n623), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n680), .A2(G1341), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U705 ( .A(n629), .B(n628), .ZN(n647) );
  INV_X1 U706 ( .A(n647), .ZN(n639) );
  NAND2_X1 U707 ( .A1(G79), .A2(n802), .ZN(n637) );
  NAND2_X1 U708 ( .A1(n795), .A2(G92), .ZN(n632) );
  NAND2_X1 U709 ( .A1(G66), .A2(n630), .ZN(n631) );
  NAND2_X1 U710 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n798), .A2(G54), .ZN(n633) );
  XOR2_X1 U712 ( .A(KEYINPUT76), .B(n633), .Z(n634) );
  NOR2_X1 U713 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n637), .A2(n636), .ZN(n638) );
  INV_X1 U715 ( .A(n919), .ZN(n957) );
  NAND2_X1 U716 ( .A1(n639), .A2(n919), .ZN(n640) );
  XNOR2_X1 U717 ( .A(n640), .B(KEYINPUT92), .ZN(n644) );
  NOR2_X1 U718 ( .A1(n657), .A2(G1348), .ZN(n642) );
  NOR2_X1 U719 ( .A1(G2067), .A2(n680), .ZN(n641) );
  NOR2_X1 U720 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U721 ( .A1(n644), .A2(n643), .ZN(n646) );
  XNOR2_X1 U722 ( .A(n646), .B(n645), .ZN(n649) );
  NAND2_X1 U723 ( .A1(n647), .A2(n957), .ZN(n648) );
  NAND2_X1 U724 ( .A1(n649), .A2(n648), .ZN(n661) );
  NAND2_X1 U725 ( .A1(n798), .A2(G53), .ZN(n651) );
  NAND2_X1 U726 ( .A1(G65), .A2(n544), .ZN(n650) );
  NAND2_X1 U727 ( .A1(n651), .A2(n650), .ZN(n655) );
  NAND2_X1 U728 ( .A1(G91), .A2(n795), .ZN(n653) );
  NAND2_X1 U729 ( .A1(G78), .A2(n802), .ZN(n652) );
  NAND2_X1 U730 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U731 ( .A1(n655), .A2(n654), .ZN(n963) );
  NAND2_X1 U732 ( .A1(n657), .A2(G2072), .ZN(n656) );
  XNOR2_X1 U733 ( .A(n656), .B(KEYINPUT27), .ZN(n659) );
  INV_X1 U734 ( .A(G1956), .ZN(n983) );
  NOR2_X1 U735 ( .A1(n983), .A2(n657), .ZN(n658) );
  NOR2_X1 U736 ( .A1(n659), .A2(n658), .ZN(n662) );
  NAND2_X1 U737 ( .A1(n963), .A2(n662), .ZN(n660) );
  NAND2_X1 U738 ( .A1(n661), .A2(n660), .ZN(n665) );
  NOR2_X1 U739 ( .A1(n963), .A2(n662), .ZN(n663) );
  XOR2_X1 U740 ( .A(n663), .B(KEYINPUT28), .Z(n664) );
  XNOR2_X1 U741 ( .A(KEYINPUT94), .B(KEYINPUT29), .ZN(n666) );
  NOR2_X1 U742 ( .A1(n668), .A2(G301), .ZN(n669) );
  NOR2_X1 U743 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U744 ( .A1(n672), .A2(n671), .ZN(n674) );
  XNOR2_X1 U745 ( .A(n674), .B(n673), .ZN(n679) );
  NAND2_X1 U746 ( .A1(G8), .A2(n675), .ZN(n676) );
  NAND2_X1 U747 ( .A1(n679), .A2(n676), .ZN(n677) );
  NOR2_X1 U748 ( .A1(n678), .A2(n677), .ZN(n691) );
  NAND2_X1 U749 ( .A1(n679), .A2(G286), .ZN(n687) );
  INV_X1 U750 ( .A(G8), .ZN(n685) );
  NOR2_X1 U751 ( .A1(G1971), .A2(n743), .ZN(n682) );
  NOR2_X1 U752 ( .A1(G2090), .A2(n680), .ZN(n681) );
  NOR2_X1 U753 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U754 ( .A1(n683), .A2(G303), .ZN(n684) );
  OR2_X1 U755 ( .A1(n685), .A2(n684), .ZN(n686) );
  AND2_X1 U756 ( .A1(n687), .A2(n686), .ZN(n689) );
  NAND2_X1 U757 ( .A1(G166), .A2(G8), .ZN(n692) );
  NOR2_X1 U758 ( .A1(G2090), .A2(n692), .ZN(n693) );
  NAND2_X1 U759 ( .A1(n694), .A2(n743), .ZN(n696) );
  INV_X1 U760 ( .A(KEYINPUT97), .ZN(n695) );
  XNOR2_X1 U761 ( .A(n696), .B(n695), .ZN(n701) );
  NOR2_X1 U762 ( .A1(G1981), .A2(G305), .ZN(n697) );
  XNOR2_X1 U763 ( .A(KEYINPUT24), .B(n697), .ZN(n698) );
  XNOR2_X1 U764 ( .A(KEYINPUT89), .B(n698), .ZN(n699) );
  OR2_X1 U765 ( .A1(n743), .A2(n699), .ZN(n700) );
  NAND2_X1 U766 ( .A1(n701), .A2(n700), .ZN(n737) );
  NOR2_X1 U767 ( .A1(n703), .A2(n702), .ZN(n767) );
  XNOR2_X1 U768 ( .A(KEYINPUT37), .B(G2067), .ZN(n765) );
  BUF_X1 U769 ( .A(n704), .Z(n895) );
  NAND2_X1 U770 ( .A1(G140), .A2(n895), .ZN(n708) );
  NAND2_X1 U771 ( .A1(G104), .A2(n706), .ZN(n707) );
  NAND2_X1 U772 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U773 ( .A(n709), .B(KEYINPUT34), .ZN(n710) );
  XNOR2_X1 U774 ( .A(n710), .B(KEYINPUT85), .ZN(n716) );
  XNOR2_X1 U775 ( .A(KEYINPUT35), .B(KEYINPUT86), .ZN(n714) );
  NAND2_X1 U776 ( .A1(G116), .A2(n899), .ZN(n712) );
  NAND2_X1 U777 ( .A1(G128), .A2(n902), .ZN(n711) );
  NAND2_X1 U778 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U779 ( .A(n714), .B(n713), .ZN(n715) );
  NAND2_X1 U780 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U781 ( .A(KEYINPUT36), .B(n717), .Z(n882) );
  NOR2_X1 U782 ( .A1(n765), .A2(n882), .ZN(n1023) );
  NAND2_X1 U783 ( .A1(n767), .A2(n1023), .ZN(n763) );
  NAND2_X1 U784 ( .A1(G117), .A2(n899), .ZN(n719) );
  NAND2_X1 U785 ( .A1(G129), .A2(n902), .ZN(n718) );
  NAND2_X1 U786 ( .A1(n719), .A2(n718), .ZN(n722) );
  NAND2_X1 U787 ( .A1(G105), .A2(n706), .ZN(n720) );
  XOR2_X1 U788 ( .A(KEYINPUT38), .B(n720), .Z(n721) );
  NOR2_X1 U789 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U790 ( .A(KEYINPUT87), .B(n723), .Z(n725) );
  NAND2_X1 U791 ( .A1(n895), .A2(G141), .ZN(n724) );
  NAND2_X1 U792 ( .A1(n725), .A2(n724), .ZN(n914) );
  NAND2_X1 U793 ( .A1(G1996), .A2(n914), .ZN(n726) );
  XOR2_X1 U794 ( .A(KEYINPUT88), .B(n726), .Z(n734) );
  NAND2_X1 U795 ( .A1(G107), .A2(n899), .ZN(n728) );
  NAND2_X1 U796 ( .A1(G131), .A2(n895), .ZN(n727) );
  NAND2_X1 U797 ( .A1(n728), .A2(n727), .ZN(n732) );
  NAND2_X1 U798 ( .A1(G119), .A2(n902), .ZN(n730) );
  NAND2_X1 U799 ( .A1(G95), .A2(n706), .ZN(n729) );
  NAND2_X1 U800 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U801 ( .A1(n732), .A2(n731), .ZN(n910) );
  INV_X1 U802 ( .A(G1991), .ZN(n756) );
  NOR2_X1 U803 ( .A1(n910), .A2(n756), .ZN(n733) );
  NOR2_X1 U804 ( .A1(n734), .A2(n733), .ZN(n755) );
  XOR2_X1 U805 ( .A(G1986), .B(G290), .Z(n955) );
  NAND2_X1 U806 ( .A1(n755), .A2(n955), .ZN(n735) );
  NAND2_X1 U807 ( .A1(n735), .A2(n767), .ZN(n736) );
  AND2_X1 U808 ( .A1(n763), .A2(n736), .ZN(n747) );
  NAND2_X1 U809 ( .A1(n737), .A2(n747), .ZN(n772) );
  INV_X1 U810 ( .A(n738), .ZN(n741) );
  NOR2_X1 U811 ( .A1(G1971), .A2(G303), .ZN(n739) );
  NOR2_X1 U812 ( .A1(G1976), .A2(G288), .ZN(n962) );
  NOR2_X1 U813 ( .A1(n739), .A2(n962), .ZN(n740) );
  NAND2_X1 U814 ( .A1(n741), .A2(n740), .ZN(n751) );
  NAND2_X1 U815 ( .A1(G1976), .A2(G288), .ZN(n960) );
  INV_X1 U816 ( .A(n960), .ZN(n742) );
  NOR2_X1 U817 ( .A1(n743), .A2(n742), .ZN(n749) );
  NAND2_X1 U818 ( .A1(n962), .A2(KEYINPUT33), .ZN(n744) );
  NOR2_X1 U819 ( .A1(n744), .A2(n743), .ZN(n746) );
  XOR2_X1 U820 ( .A(G1981), .B(G305), .Z(n952) );
  INV_X1 U821 ( .A(n952), .ZN(n745) );
  NOR2_X1 U822 ( .A1(n746), .A2(n745), .ZN(n748) );
  AND2_X1 U823 ( .A1(n748), .A2(n747), .ZN(n752) );
  AND2_X1 U824 ( .A1(n749), .A2(n752), .ZN(n750) );
  AND2_X1 U825 ( .A1(n751), .A2(n750), .ZN(n754) );
  AND2_X1 U826 ( .A1(n752), .A2(KEYINPUT33), .ZN(n753) );
  NOR2_X1 U827 ( .A1(n754), .A2(n753), .ZN(n770) );
  NOR2_X1 U828 ( .A1(G1996), .A2(n914), .ZN(n1016) );
  INV_X1 U829 ( .A(n755), .ZN(n1027) );
  AND2_X1 U830 ( .A1(n756), .A2(n910), .ZN(n757) );
  XNOR2_X1 U831 ( .A(KEYINPUT98), .B(n757), .ZN(n1019) );
  NOR2_X1 U832 ( .A1(G1986), .A2(G290), .ZN(n758) );
  NOR2_X1 U833 ( .A1(n1019), .A2(n758), .ZN(n759) );
  NOR2_X1 U834 ( .A1(n1027), .A2(n759), .ZN(n760) );
  NOR2_X1 U835 ( .A1(n1016), .A2(n760), .ZN(n761) );
  XOR2_X1 U836 ( .A(n761), .B(KEYINPUT99), .Z(n762) );
  XNOR2_X1 U837 ( .A(n762), .B(KEYINPUT39), .ZN(n764) );
  NAND2_X1 U838 ( .A1(n764), .A2(n763), .ZN(n766) );
  NAND2_X1 U839 ( .A1(n765), .A2(n882), .ZN(n1029) );
  NAND2_X1 U840 ( .A1(n766), .A2(n1029), .ZN(n768) );
  NAND2_X1 U841 ( .A1(n768), .A2(n767), .ZN(n769) );
  AND2_X1 U842 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U843 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U844 ( .A(n773), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U845 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U846 ( .A(G132), .ZN(G219) );
  INV_X1 U847 ( .A(G57), .ZN(G237) );
  INV_X1 U848 ( .A(G120), .ZN(G236) );
  NAND2_X1 U849 ( .A1(G7), .A2(G661), .ZN(n774) );
  XNOR2_X1 U850 ( .A(n774), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U851 ( .A(G223), .ZN(n834) );
  NAND2_X1 U852 ( .A1(n834), .A2(G567), .ZN(n775) );
  XOR2_X1 U853 ( .A(KEYINPUT11), .B(n775), .Z(G234) );
  INV_X1 U854 ( .A(G860), .ZN(n780) );
  OR2_X1 U855 ( .A1(n971), .A2(n780), .ZN(G153) );
  NAND2_X1 U856 ( .A1(G868), .A2(G301), .ZN(n777) );
  INV_X1 U857 ( .A(G868), .ZN(n815) );
  NAND2_X1 U858 ( .A1(n957), .A2(n815), .ZN(n776) );
  NAND2_X1 U859 ( .A1(n777), .A2(n776), .ZN(G284) );
  INV_X1 U860 ( .A(n963), .ZN(G299) );
  NOR2_X1 U861 ( .A1(G286), .A2(n815), .ZN(n779) );
  NOR2_X1 U862 ( .A1(G868), .A2(G299), .ZN(n778) );
  NOR2_X1 U863 ( .A1(n779), .A2(n778), .ZN(G297) );
  NAND2_X1 U864 ( .A1(n780), .A2(G559), .ZN(n781) );
  NAND2_X1 U865 ( .A1(n781), .A2(n919), .ZN(n782) );
  XNOR2_X1 U866 ( .A(n782), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U867 ( .A1(G868), .A2(n971), .ZN(n785) );
  NAND2_X1 U868 ( .A1(G868), .A2(n919), .ZN(n783) );
  NOR2_X1 U869 ( .A1(G559), .A2(n783), .ZN(n784) );
  NOR2_X1 U870 ( .A1(n785), .A2(n784), .ZN(G282) );
  NAND2_X1 U871 ( .A1(G111), .A2(n899), .ZN(n787) );
  NAND2_X1 U872 ( .A1(G135), .A2(n895), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U874 ( .A1(n902), .A2(G123), .ZN(n788) );
  XOR2_X1 U875 ( .A(KEYINPUT18), .B(n788), .Z(n789) );
  NOR2_X1 U876 ( .A1(n790), .A2(n789), .ZN(n792) );
  NAND2_X1 U877 ( .A1(G99), .A2(n706), .ZN(n791) );
  NAND2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n1020) );
  XNOR2_X1 U879 ( .A(G2096), .B(n1020), .ZN(n793) );
  NOR2_X1 U880 ( .A1(G2100), .A2(n793), .ZN(n794) );
  XOR2_X1 U881 ( .A(KEYINPUT78), .B(n794), .Z(G156) );
  NAND2_X1 U882 ( .A1(n795), .A2(G93), .ZN(n797) );
  NAND2_X1 U883 ( .A1(G67), .A2(n544), .ZN(n796) );
  NAND2_X1 U884 ( .A1(n797), .A2(n796), .ZN(n801) );
  NAND2_X1 U885 ( .A1(G55), .A2(n798), .ZN(n799) );
  XNOR2_X1 U886 ( .A(KEYINPUT79), .B(n799), .ZN(n800) );
  NOR2_X1 U887 ( .A1(n801), .A2(n800), .ZN(n804) );
  NAND2_X1 U888 ( .A1(n802), .A2(G80), .ZN(n803) );
  NAND2_X1 U889 ( .A1(n804), .A2(n803), .ZN(n816) );
  NAND2_X1 U890 ( .A1(n919), .A2(G559), .ZN(n813) );
  XNOR2_X1 U891 ( .A(n971), .B(n813), .ZN(n805) );
  NOR2_X1 U892 ( .A1(G860), .A2(n805), .ZN(n806) );
  XOR2_X1 U893 ( .A(n816), .B(n806), .Z(G145) );
  XOR2_X1 U894 ( .A(G290), .B(n971), .Z(n807) );
  XNOR2_X1 U895 ( .A(n816), .B(n807), .ZN(n810) );
  XNOR2_X1 U896 ( .A(KEYINPUT19), .B(G305), .ZN(n808) );
  XNOR2_X1 U897 ( .A(n808), .B(G288), .ZN(n809) );
  XOR2_X1 U898 ( .A(n810), .B(n809), .Z(n812) );
  XNOR2_X1 U899 ( .A(G166), .B(n963), .ZN(n811) );
  XNOR2_X1 U900 ( .A(n812), .B(n811), .ZN(n918) );
  XOR2_X1 U901 ( .A(n918), .B(n813), .Z(n814) );
  NAND2_X1 U902 ( .A1(G868), .A2(n814), .ZN(n818) );
  NAND2_X1 U903 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U904 ( .A1(n818), .A2(n817), .ZN(G295) );
  NAND2_X1 U905 ( .A1(G2078), .A2(G2084), .ZN(n819) );
  XOR2_X1 U906 ( .A(KEYINPUT20), .B(n819), .Z(n820) );
  NAND2_X1 U907 ( .A1(G2090), .A2(n820), .ZN(n821) );
  XNOR2_X1 U908 ( .A(KEYINPUT21), .B(n821), .ZN(n822) );
  NAND2_X1 U909 ( .A1(n822), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U910 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U911 ( .A(KEYINPUT73), .B(G82), .ZN(G220) );
  NOR2_X1 U912 ( .A1(G236), .A2(G237), .ZN(n823) );
  NAND2_X1 U913 ( .A1(G69), .A2(n823), .ZN(n824) );
  XNOR2_X1 U914 ( .A(KEYINPUT81), .B(n824), .ZN(n825) );
  NAND2_X1 U915 ( .A1(n825), .A2(G108), .ZN(n930) );
  NAND2_X1 U916 ( .A1(G567), .A2(n930), .ZN(n830) );
  NOR2_X1 U917 ( .A1(G219), .A2(G220), .ZN(n826) );
  XOR2_X1 U918 ( .A(KEYINPUT22), .B(n826), .Z(n827) );
  NOR2_X1 U919 ( .A1(G218), .A2(n827), .ZN(n828) );
  NAND2_X1 U920 ( .A1(G96), .A2(n828), .ZN(n931) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n931), .ZN(n829) );
  NAND2_X1 U922 ( .A1(n830), .A2(n829), .ZN(n831) );
  XOR2_X1 U923 ( .A(KEYINPUT82), .B(n831), .Z(G319) );
  INV_X1 U924 ( .A(G319), .ZN(n924) );
  NAND2_X1 U925 ( .A1(G661), .A2(G483), .ZN(n832) );
  NOR2_X1 U926 ( .A1(n924), .A2(n832), .ZN(n838) );
  NAND2_X1 U927 ( .A1(n838), .A2(G36), .ZN(n833) );
  XOR2_X1 U928 ( .A(KEYINPUT83), .B(n833), .Z(G176) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n834), .ZN(G217) );
  NAND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n835) );
  XNOR2_X1 U931 ( .A(KEYINPUT103), .B(n835), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n836), .A2(G661), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U934 ( .A1(n838), .A2(n837), .ZN(G188) );
  XNOR2_X1 U935 ( .A(G2443), .B(G2451), .ZN(n848) );
  XOR2_X1 U936 ( .A(G2446), .B(G2454), .Z(n840) );
  XNOR2_X1 U937 ( .A(KEYINPUT100), .B(G2435), .ZN(n839) );
  XNOR2_X1 U938 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U939 ( .A(KEYINPUT101), .B(G2438), .Z(n842) );
  XNOR2_X1 U940 ( .A(G1341), .B(G1348), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U942 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U943 ( .A(G2427), .B(G2430), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(n849) );
  NAND2_X1 U946 ( .A1(n849), .A2(G14), .ZN(n850) );
  XOR2_X1 U947 ( .A(KEYINPUT102), .B(n850), .Z(G401) );
  XOR2_X1 U948 ( .A(KEYINPUT106), .B(G2678), .Z(n852) );
  XNOR2_X1 U949 ( .A(KEYINPUT43), .B(G2096), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U951 ( .A(n853), .B(KEYINPUT42), .Z(n855) );
  XNOR2_X1 U952 ( .A(G2067), .B(G2090), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U954 ( .A(G2100), .B(G2084), .Z(n857) );
  XNOR2_X1 U955 ( .A(G2078), .B(G2072), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U957 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U958 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n860) );
  XNOR2_X1 U959 ( .A(n861), .B(n860), .ZN(G227) );
  XOR2_X1 U960 ( .A(KEYINPUT107), .B(G1956), .Z(n863) );
  XNOR2_X1 U961 ( .A(G1976), .B(G1961), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U963 ( .A(n864), .B(KEYINPUT41), .Z(n866) );
  XNOR2_X1 U964 ( .A(G1996), .B(G1991), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U966 ( .A(G1966), .B(G1971), .Z(n868) );
  XNOR2_X1 U967 ( .A(G1986), .B(G1981), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U969 ( .A(n870), .B(n869), .Z(n872) );
  XNOR2_X1 U970 ( .A(G2474), .B(KEYINPUT108), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(G229) );
  XOR2_X1 U972 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n874) );
  NAND2_X1 U973 ( .A1(G124), .A2(n902), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U975 ( .A(n875), .B(KEYINPUT109), .ZN(n877) );
  NAND2_X1 U976 ( .A1(n899), .A2(G112), .ZN(n876) );
  NAND2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n881) );
  NAND2_X1 U978 ( .A1(G136), .A2(n895), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G100), .A2(n706), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U981 ( .A1(n881), .A2(n880), .ZN(G162) );
  XNOR2_X1 U982 ( .A(G160), .B(G164), .ZN(n883) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n1020), .B(n884), .ZN(n894) );
  NAND2_X1 U985 ( .A1(G139), .A2(n895), .ZN(n886) );
  NAND2_X1 U986 ( .A1(G103), .A2(n706), .ZN(n885) );
  NAND2_X1 U987 ( .A1(n886), .A2(n885), .ZN(n892) );
  NAND2_X1 U988 ( .A1(n899), .A2(G115), .ZN(n887) );
  XOR2_X1 U989 ( .A(KEYINPUT113), .B(n887), .Z(n889) );
  NAND2_X1 U990 ( .A1(n902), .A2(G127), .ZN(n888) );
  NAND2_X1 U991 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U992 ( .A(KEYINPUT47), .B(n890), .Z(n891) );
  NOR2_X1 U993 ( .A1(n892), .A2(n891), .ZN(n1010) );
  XNOR2_X1 U994 ( .A(n1010), .B(G162), .ZN(n893) );
  XNOR2_X1 U995 ( .A(n894), .B(n893), .ZN(n916) );
  XOR2_X1 U996 ( .A(KEYINPUT115), .B(KEYINPUT46), .Z(n908) );
  NAND2_X1 U997 ( .A1(G142), .A2(n895), .ZN(n897) );
  NAND2_X1 U998 ( .A1(G106), .A2(n706), .ZN(n896) );
  NAND2_X1 U999 ( .A1(n897), .A2(n896), .ZN(n898) );
  XNOR2_X1 U1000 ( .A(n898), .B(KEYINPUT45), .ZN(n901) );
  NAND2_X1 U1001 ( .A1(G118), .A2(n899), .ZN(n900) );
  NAND2_X1 U1002 ( .A1(n901), .A2(n900), .ZN(n905) );
  NAND2_X1 U1003 ( .A1(G130), .A2(n902), .ZN(n903) );
  XNOR2_X1 U1004 ( .A(KEYINPUT111), .B(n903), .ZN(n904) );
  NOR2_X1 U1005 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(n906), .B(KEYINPUT114), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1008 ( .A(n909), .B(KEYINPUT112), .Z(n912) );
  XNOR2_X1 U1009 ( .A(n910), .B(KEYINPUT48), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1011 ( .A(n914), .B(n913), .Z(n915) );
  XNOR2_X1 U1012 ( .A(n916), .B(n915), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n917), .ZN(G395) );
  XOR2_X1 U1014 ( .A(KEYINPUT116), .B(n918), .Z(n921) );
  XNOR2_X1 U1015 ( .A(n919), .B(G286), .ZN(n920) );
  XNOR2_X1 U1016 ( .A(n921), .B(n920), .ZN(n922) );
  XNOR2_X1 U1017 ( .A(n922), .B(G301), .ZN(n923) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n923), .ZN(G397) );
  OR2_X1 U1019 ( .A1(G401), .A2(n924), .ZN(n927) );
  NOR2_X1 U1020 ( .A1(G227), .A2(G229), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(KEYINPUT49), .B(n925), .ZN(n926) );
  NOR2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(n929) );
  NOR2_X1 U1023 ( .A1(G395), .A2(G397), .ZN(n928) );
  NAND2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(G225) );
  XNOR2_X1 U1025 ( .A(KEYINPUT117), .B(G225), .ZN(G308) );
  INV_X1 U1027 ( .A(G108), .ZN(G238) );
  INV_X1 U1028 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(G325) );
  INV_X1 U1030 ( .A(G325), .ZN(G261) );
  INV_X1 U1031 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1032 ( .A(G1991), .B(G25), .ZN(n942) );
  XOR2_X1 U1033 ( .A(G2072), .B(G33), .Z(n937) );
  XNOR2_X1 U1034 ( .A(G1996), .B(G32), .ZN(n934) );
  XNOR2_X1 U1035 ( .A(n932), .B(G27), .ZN(n933) );
  NOR2_X1 U1036 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1037 ( .A(KEYINPUT120), .B(n935), .ZN(n936) );
  NAND2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n939) );
  XNOR2_X1 U1039 ( .A(G26), .B(G2067), .ZN(n938) );
  NOR2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1041 ( .A(KEYINPUT121), .B(n940), .ZN(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1043 ( .A1(G28), .A2(n943), .ZN(n944) );
  XNOR2_X1 U1044 ( .A(n944), .B(KEYINPUT53), .ZN(n947) );
  XOR2_X1 U1045 ( .A(G2084), .B(G34), .Z(n945) );
  XNOR2_X1 U1046 ( .A(KEYINPUT54), .B(n945), .ZN(n946) );
  NAND2_X1 U1047 ( .A1(n947), .A2(n946), .ZN(n949) );
  XNOR2_X1 U1048 ( .A(G35), .B(G2090), .ZN(n948) );
  NOR2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1050 ( .A(KEYINPUT55), .B(n950), .Z(n951) );
  NOR2_X1 U1051 ( .A1(G29), .A2(n951), .ZN(n1007) );
  XNOR2_X1 U1052 ( .A(G16), .B(KEYINPUT56), .ZN(n977) );
  XNOR2_X1 U1053 ( .A(G1966), .B(G168), .ZN(n953) );
  NAND2_X1 U1054 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1055 ( .A(n954), .B(KEYINPUT57), .ZN(n975) );
  XNOR2_X1 U1056 ( .A(G171), .B(G1961), .ZN(n956) );
  NAND2_X1 U1057 ( .A1(n956), .A2(n955), .ZN(n959) );
  XNOR2_X1 U1058 ( .A(G1348), .B(n957), .ZN(n958) );
  NOR2_X1 U1059 ( .A1(n959), .A2(n958), .ZN(n970) );
  XNOR2_X1 U1060 ( .A(G1971), .B(G166), .ZN(n961) );
  NAND2_X1 U1061 ( .A1(n961), .A2(n960), .ZN(n967) );
  XOR2_X1 U1062 ( .A(n962), .B(KEYINPUT122), .Z(n965) );
  XNOR2_X1 U1063 ( .A(G1956), .B(n963), .ZN(n964) );
  NAND2_X1 U1064 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1065 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1066 ( .A(KEYINPUT123), .B(n968), .Z(n969) );
  NAND2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(G1341), .B(n971), .ZN(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n1005) );
  INV_X1 U1072 ( .A(G16), .ZN(n1003) );
  XOR2_X1 U1073 ( .A(G1966), .B(G21), .Z(n989) );
  XNOR2_X1 U1074 ( .A(G1348), .B(KEYINPUT59), .ZN(n978) );
  XNOR2_X1 U1075 ( .A(n978), .B(G4), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(G1981), .B(G6), .ZN(n980) );
  XNOR2_X1 U1077 ( .A(G19), .B(G1341), .ZN(n979) );
  NOR2_X1 U1078 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1079 ( .A1(n982), .A2(n981), .ZN(n986) );
  XOR2_X1 U1080 ( .A(KEYINPUT124), .B(n983), .Z(n984) );
  XNOR2_X1 U1081 ( .A(G20), .B(n984), .ZN(n985) );
  NOR2_X1 U1082 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1083 ( .A(n987), .B(KEYINPUT60), .ZN(n988) );
  NAND2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1085 ( .A(n990), .B(KEYINPUT125), .ZN(n998) );
  XOR2_X1 U1086 ( .A(G1986), .B(KEYINPUT126), .Z(n991) );
  XNOR2_X1 U1087 ( .A(G24), .B(n991), .ZN(n995) );
  XNOR2_X1 U1088 ( .A(G1976), .B(G23), .ZN(n993) );
  XNOR2_X1 U1089 ( .A(G1971), .B(G22), .ZN(n992) );
  NOR2_X1 U1090 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1091 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1092 ( .A(KEYINPUT58), .B(n996), .Z(n997) );
  NAND2_X1 U1093 ( .A1(n998), .A2(n997), .ZN(n1000) );
  XNOR2_X1 U1094 ( .A(G5), .B(G1961), .ZN(n999) );
  NOR2_X1 U1095 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1096 ( .A(KEYINPUT61), .B(n1001), .ZN(n1002) );
  NAND2_X1 U1097 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1098 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1099 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1100 ( .A1(G11), .A2(n1008), .ZN(n1009) );
  XNOR2_X1 U1101 ( .A(n1009), .B(KEYINPUT127), .ZN(n1038) );
  XNOR2_X1 U1102 ( .A(G2072), .B(n1010), .ZN(n1013) );
  XOR2_X1 U1103 ( .A(G2078), .B(KEYINPUT119), .Z(n1011) );
  XNOR2_X1 U1104 ( .A(G164), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1105 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1106 ( .A(n1014), .B(KEYINPUT50), .ZN(n1032) );
  XOR2_X1 U1107 ( .A(G2090), .B(G162), .Z(n1015) );
  NOR2_X1 U1108 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1109 ( .A(KEYINPUT51), .B(n1017), .Z(n1025) );
  XOR2_X1 U1110 ( .A(G160), .B(G2084), .Z(n1018) );
  NOR2_X1 U1111 ( .A1(n1019), .A2(n1018), .ZN(n1021) );
  NAND2_X1 U1112 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1113 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1114 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1116 ( .A(n1028), .B(KEYINPUT118), .ZN(n1030) );
  NAND2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1118 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1119 ( .A(KEYINPUT52), .B(n1033), .ZN(n1035) );
  INV_X1 U1120 ( .A(KEYINPUT55), .ZN(n1034) );
  NAND2_X1 U1121 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1122 ( .A1(n1036), .A2(G29), .ZN(n1037) );
  NAND2_X1 U1123 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XOR2_X1 U1124 ( .A(KEYINPUT62), .B(n1039), .Z(G311) );
  INV_X1 U1125 ( .A(G311), .ZN(G150) );
endmodule

