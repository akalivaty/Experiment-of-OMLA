

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738;

  XNOR2_X1 U371 ( .A(n400), .B(n442), .ZN(n716) );
  INV_X1 U372 ( .A(G953), .ZN(n726) );
  NOR2_X1 U373 ( .A1(n614), .A2(n710), .ZN(n616) );
  NOR2_X1 U374 ( .A1(n518), .A2(n517), .ZN(n361) );
  XNOR2_X2 U375 ( .A(n383), .B(n452), .ZN(n529) );
  NOR2_X2 U376 ( .A1(n571), .A2(n451), .ZN(n383) );
  AND2_X2 U377 ( .A1(n515), .A2(n665), .ZN(n482) );
  XNOR2_X2 U378 ( .A(KEYINPUT82), .B(KEYINPUT18), .ZN(n435) );
  XOR2_X2 U379 ( .A(G116), .B(G107), .Z(n502) );
  XNOR2_X2 U380 ( .A(n432), .B(n419), .ZN(n462) );
  XNOR2_X2 U381 ( .A(n501), .B(n396), .ZN(n432) );
  NOR2_X1 U382 ( .A1(n634), .A2(n630), .ZN(n574) );
  NOR2_X1 U383 ( .A1(n527), .A2(n526), .ZN(n653) );
  XNOR2_X1 U384 ( .A(n454), .B(G472), .ZN(n663) );
  OR2_X1 U385 ( .A1(n692), .A2(G902), .ZN(n385) );
  XNOR2_X1 U386 ( .A(n462), .B(KEYINPUT97), .ZN(n722) );
  XNOR2_X1 U387 ( .A(KEYINPUT17), .B(KEYINPUT95), .ZN(n436) );
  XNOR2_X1 U388 ( .A(n349), .B(G122), .ZN(n491) );
  XNOR2_X1 U389 ( .A(G113), .B(G104), .ZN(n349) );
  XNOR2_X2 U390 ( .A(G143), .B(G128), .ZN(n501) );
  XNOR2_X2 U391 ( .A(KEYINPUT77), .B(n482), .ZN(n531) );
  XNOR2_X1 U392 ( .A(n412), .B(KEYINPUT38), .ZN(n651) );
  AND2_X1 U393 ( .A1(n380), .A2(n724), .ZN(n605) );
  NOR2_X1 U394 ( .A1(n550), .A2(n391), .ZN(n367) );
  NOR2_X1 U395 ( .A1(n568), .A2(n409), .ZN(n569) );
  XNOR2_X1 U396 ( .A(n410), .B(KEYINPUT87), .ZN(n409) );
  INV_X1 U397 ( .A(KEYINPUT4), .ZN(n396) );
  XOR2_X1 U398 ( .A(KEYINPUT71), .B(G110), .Z(n458) );
  XNOR2_X1 U399 ( .A(n398), .B(n416), .ZN(n442) );
  XNOR2_X1 U400 ( .A(n415), .B(n399), .ZN(n398) );
  INV_X1 U401 ( .A(KEYINPUT94), .ZN(n399) );
  XNOR2_X1 U402 ( .A(n596), .B(n595), .ZN(n603) );
  XNOR2_X1 U403 ( .A(KEYINPUT48), .B(KEYINPUT90), .ZN(n595) );
  NAND2_X1 U404 ( .A1(n364), .A2(n362), .ZN(n596) );
  XNOR2_X1 U405 ( .A(n363), .B(n357), .ZN(n362) );
  NAND2_X1 U406 ( .A1(n651), .A2(n390), .ZN(n388) );
  XNOR2_X1 U407 ( .A(n562), .B(n466), .ZN(n515) );
  XNOR2_X1 U408 ( .A(n465), .B(KEYINPUT65), .ZN(n466) );
  XNOR2_X1 U409 ( .A(n538), .B(n537), .ZN(n539) );
  INV_X1 U410 ( .A(KEYINPUT45), .ZN(n537) );
  XNOR2_X1 U411 ( .A(n394), .B(n393), .ZN(n392) );
  INV_X1 U412 ( .A(G140), .ZN(n393) );
  XNOR2_X1 U413 ( .A(KEYINPUT68), .B(KEYINPUT10), .ZN(n394) );
  XNOR2_X1 U414 ( .A(G119), .B(G137), .ZN(n468) );
  XOR2_X1 U415 ( .A(KEYINPUT88), .B(KEYINPUT8), .Z(n472) );
  XNOR2_X1 U416 ( .A(n491), .B(n401), .ZN(n400) );
  XNOR2_X1 U417 ( .A(n502), .B(n441), .ZN(n401) );
  XOR2_X1 U418 ( .A(KEYINPUT16), .B(KEYINPUT75), .Z(n441) );
  XNOR2_X1 U419 ( .A(n556), .B(n555), .ZN(n679) );
  XNOR2_X1 U420 ( .A(n359), .B(n378), .ZN(n511) );
  INV_X1 U421 ( .A(KEYINPUT34), .ZN(n378) );
  XNOR2_X1 U422 ( .A(n381), .B(n356), .ZN(n518) );
  NOR2_X1 U423 ( .A1(n529), .A2(n382), .ZN(n381) );
  NAND2_X1 U424 ( .A1(n653), .A2(n660), .ZN(n382) );
  INV_X1 U425 ( .A(n397), .ZN(n412) );
  XNOR2_X1 U426 ( .A(n549), .B(KEYINPUT30), .ZN(n550) );
  XNOR2_X1 U427 ( .A(n384), .B(n370), .ZN(n546) );
  INV_X1 U428 ( .A(KEYINPUT98), .ZN(n370) );
  NOR2_X1 U429 ( .A1(G902), .A2(n453), .ZN(n454) );
  XNOR2_X1 U430 ( .A(G119), .B(G101), .ZN(n415) );
  NOR2_X1 U431 ( .A1(n586), .A2(n365), .ZN(n364) );
  INV_X1 U432 ( .A(n639), .ZN(n365) );
  XOR2_X1 U433 ( .A(G146), .B(G113), .Z(n421) );
  XNOR2_X1 U434 ( .A(G143), .B(G131), .ZN(n485) );
  NOR2_X1 U435 ( .A1(G953), .A2(G237), .ZN(n488) );
  INV_X1 U436 ( .A(G137), .ZN(n417) );
  NAND2_X1 U437 ( .A1(G234), .A2(G237), .ZN(n446) );
  XNOR2_X1 U438 ( .A(n554), .B(KEYINPUT111), .ZN(n655) );
  NAND2_X1 U439 ( .A1(n375), .A2(n484), .ZN(n374) );
  NOR2_X1 U440 ( .A1(n529), .A2(n372), .ZN(n371) );
  INV_X1 U441 ( .A(n376), .ZN(n372) );
  AND2_X1 U442 ( .A1(n514), .A2(n660), .ZN(n665) );
  XNOR2_X1 U443 ( .A(n458), .B(n351), .ZN(n459) );
  XNOR2_X1 U444 ( .A(G101), .B(G146), .ZN(n456) );
  XOR2_X1 U445 ( .A(G107), .B(G104), .Z(n457) );
  INV_X1 U446 ( .A(n641), .ZN(n408) );
  NAND2_X1 U447 ( .A1(n350), .A2(n406), .ZN(n395) );
  INV_X1 U448 ( .A(n642), .ZN(n406) );
  NAND2_X1 U449 ( .A1(n389), .A2(n386), .ZN(n604) );
  NAND2_X1 U450 ( .A1(n368), .A2(n387), .ZN(n386) );
  NOR2_X1 U451 ( .A1(n550), .A2(n388), .ZN(n387) );
  XNOR2_X1 U452 ( .A(n475), .B(n405), .ZN(n708) );
  XNOR2_X1 U453 ( .A(n470), .B(n723), .ZN(n405) );
  BUF_X1 U454 ( .A(n696), .Z(n706) );
  XNOR2_X1 U455 ( .A(n440), .B(n433), .ZN(n403) );
  NOR2_X1 U456 ( .A1(G952), .A2(n726), .ZN(n710) );
  NOR2_X1 U457 ( .A1(n679), .A2(n570), .ZN(n564) );
  XNOR2_X1 U458 ( .A(n553), .B(KEYINPUT40), .ZN(n736) );
  NAND2_X1 U459 ( .A1(n604), .A2(n630), .ZN(n553) );
  INV_X1 U460 ( .A(KEYINPUT35), .ZN(n512) );
  XNOR2_X1 U461 ( .A(n361), .B(KEYINPUT32), .ZN(n735) );
  NOR2_X1 U462 ( .A1(n567), .A2(n412), .ZN(n411) );
  AND2_X1 U463 ( .A1(n524), .A2(n519), .ZN(n623) );
  NOR2_X1 U464 ( .A1(n530), .A2(n369), .ZN(n619) );
  XNOR2_X1 U465 ( .A(KEYINPUT83), .B(n607), .ZN(n350) );
  AND2_X1 U466 ( .A1(G227), .A2(n726), .ZN(n351) );
  AND2_X1 U467 ( .A1(G210), .A2(n444), .ZN(n352) );
  XNOR2_X1 U468 ( .A(n547), .B(KEYINPUT80), .ZN(n551) );
  AND2_X1 U469 ( .A1(n373), .A2(n371), .ZN(n353) );
  AND2_X1 U470 ( .A1(n373), .A2(n376), .ZN(n354) );
  XOR2_X1 U471 ( .A(KEYINPUT69), .B(G469), .Z(n355) );
  XOR2_X1 U472 ( .A(KEYINPUT22), .B(KEYINPUT74), .Z(n356) );
  XNOR2_X1 U473 ( .A(KEYINPUT91), .B(KEYINPUT46), .ZN(n357) );
  XNOR2_X1 U474 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n358) );
  XNOR2_X1 U475 ( .A(n463), .B(n464), .ZN(n692) );
  NAND2_X1 U476 ( .A1(n353), .A2(n377), .ZN(n359) );
  NOR2_X2 U477 ( .A1(n710), .A2(n700), .ZN(n702) );
  XNOR2_X1 U478 ( .A(n360), .B(KEYINPUT44), .ZN(n536) );
  NOR2_X2 U479 ( .A1(n523), .A2(n734), .ZN(n360) );
  XNOR2_X2 U480 ( .A(n540), .B(n539), .ZN(n380) );
  NOR2_X2 U481 ( .A1(n710), .A2(n689), .ZN(n690) );
  NOR2_X2 U482 ( .A1(n605), .A2(KEYINPUT2), .ZN(n611) );
  NAND2_X1 U483 ( .A1(n696), .A2(G210), .ZN(n688) );
  NAND2_X1 U484 ( .A1(n380), .A2(n608), .ZN(n645) );
  NAND2_X1 U485 ( .A1(n736), .A2(n737), .ZN(n363) );
  XNOR2_X1 U486 ( .A(n402), .B(n716), .ZN(n686) );
  NOR2_X2 U487 ( .A1(n603), .A2(n407), .ZN(n724) );
  NAND2_X1 U488 ( .A1(n366), .A2(n552), .ZN(n389) );
  NAND2_X1 U489 ( .A1(n368), .A2(n367), .ZN(n366) );
  INV_X1 U490 ( .A(n551), .ZN(n368) );
  INV_X1 U491 ( .A(n546), .ZN(n369) );
  NAND2_X1 U492 ( .A1(n354), .A2(n377), .ZN(n680) );
  OR2_X2 U493 ( .A1(n531), .A2(n374), .ZN(n373) );
  INV_X1 U494 ( .A(n587), .ZN(n375) );
  NAND2_X1 U495 ( .A1(n587), .A2(n379), .ZN(n376) );
  NAND2_X1 U496 ( .A1(n531), .A2(n379), .ZN(n377) );
  INV_X1 U497 ( .A(n484), .ZN(n379) );
  NOR2_X1 U498 ( .A1(n380), .A2(KEYINPUT2), .ZN(n644) );
  NAND2_X1 U499 ( .A1(n380), .A2(n726), .ZN(n714) );
  XNOR2_X1 U500 ( .A(n439), .B(n434), .ZN(n404) );
  XNOR2_X1 U501 ( .A(n404), .B(n403), .ZN(n402) );
  XNOR2_X2 U502 ( .A(n513), .B(n512), .ZN(n734) );
  INV_X1 U503 ( .A(n514), .ZN(n557) );
  NAND2_X1 U504 ( .A1(n562), .A2(n665), .ZN(n384) );
  XNOR2_X2 U505 ( .A(n385), .B(n355), .ZN(n562) );
  NOR2_X1 U506 ( .A1(n551), .A2(n550), .ZN(n566) );
  INV_X1 U507 ( .A(n552), .ZN(n390) );
  INV_X1 U508 ( .A(n651), .ZN(n391) );
  XNOR2_X2 U509 ( .A(n392), .B(n467), .ZN(n723) );
  NOR2_X1 U510 ( .A1(n603), .A2(n395), .ZN(n608) );
  NAND2_X1 U511 ( .A1(n397), .A2(n650), .ZN(n592) );
  XNOR2_X2 U512 ( .A(n443), .B(n352), .ZN(n397) );
  NOR2_X1 U513 ( .A1(n602), .A2(n397), .ZN(n642) );
  OR2_X1 U514 ( .A1(n642), .A2(n408), .ZN(n407) );
  INV_X1 U515 ( .A(n410), .ZN(n627) );
  NAND2_X1 U516 ( .A1(n566), .A2(n411), .ZN(n410) );
  XNOR2_X1 U517 ( .A(n686), .B(n358), .ZN(n687) );
  XNOR2_X1 U518 ( .A(KEYINPUT59), .B(KEYINPUT123), .ZN(n413) );
  OR2_X1 U519 ( .A1(n574), .A2(n534), .ZN(n414) );
  NAND2_X1 U520 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U521 ( .A(n436), .B(n435), .ZN(n438) );
  XNOR2_X1 U522 ( .A(n418), .B(n417), .ZN(n419) );
  INV_X1 U523 ( .A(n559), .ZN(n545) );
  XNOR2_X1 U524 ( .A(n460), .B(n459), .ZN(n461) );
  INV_X1 U525 ( .A(KEYINPUT41), .ZN(n555) );
  INV_X1 U526 ( .A(KEYINPUT1), .ZN(n465) );
  XNOR2_X1 U527 ( .A(n697), .B(n413), .ZN(n698) );
  INV_X1 U528 ( .A(KEYINPUT63), .ZN(n615) );
  XOR2_X1 U529 ( .A(KEYINPUT113), .B(KEYINPUT62), .Z(n431) );
  XOR2_X1 U530 ( .A(KEYINPUT70), .B(KEYINPUT3), .Z(n416) );
  XNOR2_X1 U531 ( .A(G131), .B(G134), .ZN(n418) );
  XOR2_X1 U532 ( .A(n442), .B(n462), .Z(n429) );
  NAND2_X1 U533 ( .A1(n488), .A2(G210), .ZN(n420) );
  XNOR2_X1 U534 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U535 ( .A(n422), .B(KEYINPUT100), .Z(n427) );
  XOR2_X1 U536 ( .A(KEYINPUT79), .B(KEYINPUT5), .Z(n424) );
  XNOR2_X1 U537 ( .A(KEYINPUT99), .B(KEYINPUT78), .ZN(n423) );
  XNOR2_X1 U538 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U539 ( .A(n425), .B(G116), .ZN(n426) );
  XNOR2_X1 U540 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U541 ( .A(n429), .B(n428), .ZN(n453) );
  XNOR2_X1 U542 ( .A(n453), .B(KEYINPUT114), .ZN(n430) );
  XNOR2_X1 U543 ( .A(n431), .B(n430), .ZN(n613) );
  INV_X1 U544 ( .A(n432), .ZN(n434) );
  INV_X1 U545 ( .A(KEYINPUT93), .ZN(n433) );
  NAND2_X1 U546 ( .A1(G224), .A2(n726), .ZN(n437) );
  XNOR2_X1 U547 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X2 U548 ( .A(G146), .B(G125), .Z(n467) );
  XNOR2_X1 U549 ( .A(n458), .B(n467), .ZN(n440) );
  XNOR2_X1 U550 ( .A(G902), .B(KEYINPUT15), .ZN(n606) );
  NAND2_X1 U551 ( .A1(n686), .A2(n606), .ZN(n443) );
  OR2_X1 U552 ( .A1(G237), .A2(G902), .ZN(n444) );
  NAND2_X1 U553 ( .A1(G214), .A2(n444), .ZN(n650) );
  XOR2_X1 U554 ( .A(KEYINPUT19), .B(KEYINPUT66), .Z(n445) );
  XNOR2_X1 U555 ( .A(n592), .B(n445), .ZN(n571) );
  XOR2_X1 U556 ( .A(KEYINPUT14), .B(KEYINPUT96), .Z(n447) );
  XOR2_X1 U557 ( .A(n447), .B(n446), .Z(n448) );
  NAND2_X1 U558 ( .A1(G952), .A2(n448), .ZN(n678) );
  NOR2_X1 U559 ( .A1(G953), .A2(n678), .ZN(n544) );
  AND2_X1 U560 ( .A1(n448), .A2(G953), .ZN(n449) );
  NAND2_X1 U561 ( .A1(G902), .A2(n449), .ZN(n541) );
  NOR2_X1 U562 ( .A1(n541), .A2(G898), .ZN(n450) );
  NOR2_X1 U563 ( .A1(n544), .A2(n450), .ZN(n451) );
  INV_X1 U564 ( .A(KEYINPUT0), .ZN(n452) );
  XNOR2_X1 U565 ( .A(KEYINPUT105), .B(KEYINPUT6), .ZN(n455) );
  XNOR2_X1 U566 ( .A(n455), .B(n663), .ZN(n587) );
  XNOR2_X1 U567 ( .A(n457), .B(n456), .ZN(n460) );
  XOR2_X1 U568 ( .A(n461), .B(KEYINPUT81), .Z(n464) );
  XNOR2_X1 U569 ( .A(n722), .B(G140), .ZN(n463) );
  XOR2_X1 U570 ( .A(G110), .B(G128), .Z(n469) );
  XNOR2_X1 U571 ( .A(n469), .B(n468), .ZN(n470) );
  XOR2_X1 U572 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n474) );
  NAND2_X1 U573 ( .A1(G234), .A2(n726), .ZN(n471) );
  XNOR2_X1 U574 ( .A(n472), .B(n471), .ZN(n506) );
  NAND2_X1 U575 ( .A1(G221), .A2(n506), .ZN(n473) );
  XNOR2_X1 U576 ( .A(n474), .B(n473), .ZN(n475) );
  NOR2_X1 U577 ( .A1(G902), .A2(n708), .ZN(n479) );
  NAND2_X1 U578 ( .A1(G234), .A2(n606), .ZN(n476) );
  XNOR2_X1 U579 ( .A(KEYINPUT20), .B(n476), .ZN(n480) );
  NAND2_X1 U580 ( .A1(n480), .A2(G217), .ZN(n477) );
  XNOR2_X1 U581 ( .A(n477), .B(KEYINPUT25), .ZN(n478) );
  XNOR2_X1 U582 ( .A(n479), .B(n478), .ZN(n514) );
  NAND2_X1 U583 ( .A1(n480), .A2(G221), .ZN(n481) );
  XOR2_X1 U584 ( .A(KEYINPUT21), .B(n481), .Z(n660) );
  XNOR2_X1 U585 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n483) );
  XNOR2_X1 U586 ( .A(n483), .B(KEYINPUT106), .ZN(n484) );
  XNOR2_X1 U587 ( .A(KEYINPUT13), .B(G475), .ZN(n494) );
  XOR2_X1 U588 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n486) );
  XNOR2_X1 U589 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U590 ( .A(n723), .B(n487), .Z(n490) );
  NAND2_X1 U591 ( .A1(G214), .A2(n488), .ZN(n489) );
  XNOR2_X1 U592 ( .A(n490), .B(n489), .ZN(n492) );
  XOR2_X1 U593 ( .A(n492), .B(n491), .Z(n697) );
  NOR2_X1 U594 ( .A1(G902), .A2(n697), .ZN(n493) );
  XNOR2_X1 U595 ( .A(n494), .B(n493), .ZN(n527) );
  XOR2_X1 U596 ( .A(KEYINPUT104), .B(KEYINPUT9), .Z(n496) );
  XNOR2_X1 U597 ( .A(G134), .B(KEYINPUT7), .ZN(n495) );
  XNOR2_X1 U598 ( .A(n496), .B(n495), .ZN(n500) );
  XOR2_X1 U599 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n498) );
  XNOR2_X1 U600 ( .A(G122), .B(KEYINPUT103), .ZN(n497) );
  XNOR2_X1 U601 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U602 ( .A(n500), .B(n499), .Z(n505) );
  INV_X1 U603 ( .A(n501), .ZN(n503) );
  XNOR2_X1 U604 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U605 ( .A(n505), .B(n504), .ZN(n508) );
  NAND2_X1 U606 ( .A1(G217), .A2(n506), .ZN(n507) );
  XOR2_X1 U607 ( .A(n508), .B(n507), .Z(n704) );
  NOR2_X1 U608 ( .A1(G902), .A2(n704), .ZN(n509) );
  XOR2_X1 U609 ( .A(G478), .B(n509), .Z(n526) );
  NAND2_X1 U610 ( .A1(n527), .A2(n526), .ZN(n567) );
  INV_X1 U611 ( .A(n567), .ZN(n510) );
  AND2_X2 U612 ( .A1(n511), .A2(n510), .ZN(n513) );
  BUF_X1 U613 ( .A(n515), .Z(n664) );
  AND2_X1 U614 ( .A1(n557), .A2(n664), .ZN(n516) );
  NAND2_X1 U615 ( .A1(n587), .A2(n516), .ZN(n517) );
  INV_X1 U616 ( .A(n735), .ZN(n521) );
  NOR2_X1 U617 ( .A1(n664), .A2(n518), .ZN(n524) );
  INV_X1 U618 ( .A(n663), .ZN(n560) );
  NOR2_X1 U619 ( .A1(n560), .A2(n514), .ZN(n519) );
  INV_X1 U620 ( .A(n623), .ZN(n520) );
  XNOR2_X1 U621 ( .A(n522), .B(KEYINPUT92), .ZN(n523) );
  AND2_X1 U622 ( .A1(n524), .A2(n587), .ZN(n525) );
  NAND2_X1 U623 ( .A1(n525), .A2(n514), .ZN(n617) );
  INV_X1 U624 ( .A(n526), .ZN(n528) );
  NOR2_X1 U625 ( .A1(n527), .A2(n528), .ZN(n634) );
  NAND2_X1 U626 ( .A1(n528), .A2(n527), .ZN(n588) );
  INV_X1 U627 ( .A(n588), .ZN(n630) );
  INV_X1 U628 ( .A(n529), .ZN(n532) );
  NAND2_X1 U629 ( .A1(n663), .A2(n532), .ZN(n530) );
  NOR2_X1 U630 ( .A1(n663), .A2(n531), .ZN(n671) );
  NAND2_X1 U631 ( .A1(n671), .A2(n532), .ZN(n533) );
  XNOR2_X1 U632 ( .A(KEYINPUT31), .B(n533), .ZN(n635) );
  NOR2_X1 U633 ( .A1(n619), .A2(n635), .ZN(n534) );
  AND2_X1 U634 ( .A1(n617), .A2(n414), .ZN(n535) );
  NAND2_X1 U635 ( .A1(n536), .A2(n535), .ZN(n540) );
  INV_X1 U636 ( .A(KEYINPUT64), .ZN(n538) );
  XOR2_X1 U637 ( .A(KEYINPUT73), .B(KEYINPUT39), .Z(n552) );
  NOR2_X1 U638 ( .A1(G900), .A2(n541), .ZN(n542) );
  XOR2_X1 U639 ( .A(KEYINPUT107), .B(n542), .Z(n543) );
  NOR2_X1 U640 ( .A1(n544), .A2(n543), .ZN(n559) );
  NAND2_X1 U641 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U642 ( .A1(n650), .A2(n560), .ZN(n548) );
  XNOR2_X1 U643 ( .A(n548), .B(KEYINPUT110), .ZN(n549) );
  NAND2_X1 U644 ( .A1(n650), .A2(n651), .ZN(n554) );
  NAND2_X1 U645 ( .A1(n655), .A2(n653), .ZN(n556) );
  NAND2_X1 U646 ( .A1(n557), .A2(n660), .ZN(n558) );
  NOR2_X1 U647 ( .A1(n559), .A2(n558), .ZN(n590) );
  AND2_X1 U648 ( .A1(n560), .A2(n590), .ZN(n561) );
  XNOR2_X1 U649 ( .A(KEYINPUT28), .B(n561), .ZN(n563) );
  NAND2_X1 U650 ( .A1(n563), .A2(n562), .ZN(n570) );
  XOR2_X1 U651 ( .A(KEYINPUT42), .B(n564), .Z(n737) );
  NAND2_X1 U652 ( .A1(n574), .A2(KEYINPUT47), .ZN(n565) );
  XOR2_X1 U653 ( .A(KEYINPUT86), .B(n565), .Z(n568) );
  XNOR2_X1 U654 ( .A(n569), .B(KEYINPUT84), .ZN(n585) );
  NOR2_X1 U655 ( .A1(n571), .A2(n570), .ZN(n628) );
  NAND2_X1 U656 ( .A1(KEYINPUT76), .A2(n628), .ZN(n573) );
  INV_X1 U657 ( .A(KEYINPUT85), .ZN(n581) );
  AND2_X1 U658 ( .A1(n581), .A2(KEYINPUT47), .ZN(n572) );
  NAND2_X1 U659 ( .A1(n573), .A2(n572), .ZN(n580) );
  INV_X1 U660 ( .A(n574), .ZN(n654) );
  XNOR2_X1 U661 ( .A(KEYINPUT76), .B(n654), .ZN(n576) );
  INV_X1 U662 ( .A(KEYINPUT47), .ZN(n575) );
  NAND2_X1 U663 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U664 ( .A1(n577), .A2(n581), .ZN(n578) );
  NAND2_X1 U665 ( .A1(n578), .A2(n628), .ZN(n579) );
  NAND2_X1 U666 ( .A1(n580), .A2(n579), .ZN(n583) );
  NOR2_X1 U667 ( .A1(KEYINPUT47), .A2(n581), .ZN(n582) );
  NOR2_X1 U668 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U669 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U670 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U671 ( .A1(n590), .A2(n589), .ZN(n598) );
  XNOR2_X1 U672 ( .A(KEYINPUT112), .B(n598), .ZN(n591) );
  NOR2_X1 U673 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U674 ( .A(n593), .B(KEYINPUT36), .ZN(n594) );
  NAND2_X1 U675 ( .A1(n594), .A2(n664), .ZN(n639) );
  XOR2_X1 U676 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n597) );
  XNOR2_X1 U677 ( .A(KEYINPUT108), .B(n597), .ZN(n601) );
  NOR2_X1 U678 ( .A1(n664), .A2(n598), .ZN(n599) );
  NAND2_X1 U679 ( .A1(n599), .A2(n650), .ZN(n600) );
  XOR2_X1 U680 ( .A(n601), .B(n600), .Z(n602) );
  NAND2_X1 U681 ( .A1(n604), .A2(n634), .ZN(n641) );
  INV_X1 U682 ( .A(n606), .ZN(n609) );
  NAND2_X1 U683 ( .A1(KEYINPUT2), .A2(n641), .ZN(n607) );
  NAND2_X1 U684 ( .A1(n609), .A2(n645), .ZN(n610) );
  NOR2_X4 U685 ( .A1(n611), .A2(n610), .ZN(n696) );
  NAND2_X1 U686 ( .A1(n696), .A2(G472), .ZN(n612) );
  XNOR2_X1 U687 ( .A(n613), .B(n612), .ZN(n614) );
  XNOR2_X1 U688 ( .A(n616), .B(n615), .ZN(G57) );
  XNOR2_X1 U689 ( .A(G101), .B(n617), .ZN(G3) );
  NAND2_X1 U690 ( .A1(n619), .A2(n630), .ZN(n618) );
  XNOR2_X1 U691 ( .A(n618), .B(G104), .ZN(G6) );
  XOR2_X1 U692 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n621) );
  NAND2_X1 U693 ( .A1(n619), .A2(n634), .ZN(n620) );
  XNOR2_X1 U694 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U695 ( .A(G107), .B(n622), .ZN(G9) );
  XOR2_X1 U696 ( .A(n623), .B(G110), .Z(G12) );
  XOR2_X1 U697 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n625) );
  NAND2_X1 U698 ( .A1(n628), .A2(n634), .ZN(n624) );
  XNOR2_X1 U699 ( .A(n625), .B(n624), .ZN(n626) );
  XOR2_X1 U700 ( .A(G128), .B(n626), .Z(G30) );
  XOR2_X1 U701 ( .A(G143), .B(n627), .Z(G45) );
  NAND2_X1 U702 ( .A1(n628), .A2(n630), .ZN(n629) );
  XNOR2_X1 U703 ( .A(n629), .B(G146), .ZN(G48) );
  XOR2_X1 U704 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n632) );
  NAND2_X1 U705 ( .A1(n635), .A2(n630), .ZN(n631) );
  XNOR2_X1 U706 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U707 ( .A(G113), .B(n633), .ZN(G15) );
  NAND2_X1 U708 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U709 ( .A(n636), .B(KEYINPUT118), .ZN(n637) );
  XNOR2_X1 U710 ( .A(G116), .B(n637), .ZN(G18) );
  XOR2_X1 U711 ( .A(G125), .B(KEYINPUT37), .Z(n638) );
  XNOR2_X1 U712 ( .A(n639), .B(n638), .ZN(G27) );
  XOR2_X1 U713 ( .A(G134), .B(KEYINPUT119), .Z(n640) );
  XNOR2_X1 U714 ( .A(n641), .B(n640), .ZN(G36) );
  XOR2_X1 U715 ( .A(G140), .B(n642), .Z(n643) );
  XNOR2_X1 U716 ( .A(KEYINPUT120), .B(n643), .ZN(G42) );
  XNOR2_X1 U717 ( .A(n644), .B(KEYINPUT89), .ZN(n646) );
  NAND2_X1 U718 ( .A1(n646), .A2(n645), .ZN(n648) );
  NOR2_X1 U719 ( .A1(KEYINPUT2), .A2(n724), .ZN(n647) );
  NOR2_X1 U720 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U721 ( .A1(G953), .A2(n649), .ZN(n684) );
  OR2_X1 U722 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U723 ( .A1(n653), .A2(n652), .ZN(n657) );
  NAND2_X1 U724 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U726 ( .A(KEYINPUT122), .B(n658), .Z(n659) );
  NOR2_X1 U727 ( .A1(n680), .A2(n659), .ZN(n675) );
  NOR2_X1 U728 ( .A1(n660), .A2(n514), .ZN(n661) );
  XNOR2_X1 U729 ( .A(n661), .B(KEYINPUT49), .ZN(n662) );
  NAND2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n668) );
  NOR2_X1 U731 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U732 ( .A(n666), .B(KEYINPUT50), .ZN(n667) );
  NOR2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U734 ( .A(KEYINPUT121), .B(n669), .Z(n670) );
  NOR2_X1 U735 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U736 ( .A(KEYINPUT51), .B(n672), .Z(n673) );
  NOR2_X1 U737 ( .A1(n679), .A2(n673), .ZN(n674) );
  NOR2_X1 U738 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U739 ( .A(n676), .B(KEYINPUT52), .ZN(n677) );
  NOR2_X1 U740 ( .A1(n678), .A2(n677), .ZN(n682) );
  NOR2_X1 U741 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U742 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U743 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U744 ( .A(KEYINPUT53), .B(n685), .Z(G75) );
  XNOR2_X1 U745 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U746 ( .A(n690), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U747 ( .A1(n706), .A2(G469), .ZN(n694) );
  XOR2_X1 U748 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n691) );
  XNOR2_X1 U749 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U750 ( .A(n694), .B(n693), .ZN(n695) );
  NOR2_X1 U751 ( .A1(n710), .A2(n695), .ZN(G54) );
  NAND2_X1 U752 ( .A1(n696), .A2(G475), .ZN(n699) );
  XNOR2_X1 U753 ( .A(n699), .B(n698), .ZN(n700) );
  XOR2_X1 U754 ( .A(KEYINPUT67), .B(KEYINPUT60), .Z(n701) );
  XNOR2_X1 U755 ( .A(n702), .B(n701), .ZN(G60) );
  NAND2_X1 U756 ( .A1(G478), .A2(n706), .ZN(n703) );
  XNOR2_X1 U757 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U758 ( .A1(n710), .A2(n705), .ZN(G63) );
  NAND2_X1 U759 ( .A1(G217), .A2(n706), .ZN(n707) );
  XNOR2_X1 U760 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U761 ( .A1(n710), .A2(n709), .ZN(G66) );
  NAND2_X1 U762 ( .A1(G953), .A2(G224), .ZN(n711) );
  XNOR2_X1 U763 ( .A(KEYINPUT61), .B(n711), .ZN(n712) );
  NAND2_X1 U764 ( .A1(n712), .A2(G898), .ZN(n713) );
  XNOR2_X1 U765 ( .A(n713), .B(KEYINPUT124), .ZN(n715) );
  NAND2_X1 U766 ( .A1(n715), .A2(n714), .ZN(n721) );
  XOR2_X1 U767 ( .A(G110), .B(n716), .Z(n718) );
  NOR2_X1 U768 ( .A1(G898), .A2(n726), .ZN(n717) );
  NOR2_X1 U769 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U770 ( .A(KEYINPUT125), .B(n719), .Z(n720) );
  XNOR2_X1 U771 ( .A(n721), .B(n720), .ZN(G69) );
  XNOR2_X1 U772 ( .A(n722), .B(n723), .ZN(n728) );
  INV_X1 U773 ( .A(n728), .ZN(n725) );
  XNOR2_X1 U774 ( .A(n725), .B(n724), .ZN(n727) );
  NAND2_X1 U775 ( .A1(n727), .A2(n726), .ZN(n733) );
  XNOR2_X1 U776 ( .A(G227), .B(KEYINPUT126), .ZN(n729) );
  XNOR2_X1 U777 ( .A(n729), .B(n728), .ZN(n730) );
  NAND2_X1 U778 ( .A1(G900), .A2(n730), .ZN(n731) );
  NAND2_X1 U779 ( .A1(n731), .A2(G953), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n733), .A2(n732), .ZN(G72) );
  XOR2_X1 U781 ( .A(n734), .B(G122), .Z(G24) );
  XOR2_X1 U782 ( .A(n735), .B(G119), .Z(G21) );
  XNOR2_X1 U783 ( .A(n736), .B(G131), .ZN(G33) );
  XOR2_X1 U784 ( .A(G137), .B(n737), .Z(n738) );
  XNOR2_X1 U785 ( .A(KEYINPUT127), .B(n738), .ZN(G39) );
endmodule

