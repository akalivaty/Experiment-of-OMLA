//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n203), .A2(G1gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT86), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n205), .A2(new_n208), .A3(G8gat), .ZN(new_n209));
  INV_X1    g008(.A(G8gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n204), .B(new_n207), .C1(KEYINPUT86), .C2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  XOR2_X1   g012(.A(G43gat), .B(G50gat), .Z(new_n214));
  NOR2_X1   g013(.A1(G29gat), .A2(G36gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT14), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(KEYINPUT85), .B(G36gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT15), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n214), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n215), .B(KEYINPUT14), .ZN(new_n223));
  INV_X1    g022(.A(new_n219), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n223), .B1(G29gat), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT15), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT17), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n225), .A2(KEYINPUT15), .A3(new_n214), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n228), .B1(new_n227), .B2(new_n229), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n202), .B(new_n213), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G229gat), .A2(G233gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n232), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n212), .B1(new_n235), .B2(new_n230), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n227), .A2(new_n229), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT87), .B1(new_n237), .B2(new_n212), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n233), .B(new_n234), .C1(new_n236), .C2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT88), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n213), .B1(new_n231), .B2(new_n232), .ZN(new_n241));
  INV_X1    g040(.A(new_n238), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT88), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n243), .A2(new_n244), .A3(new_n234), .A4(new_n233), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT18), .B1(new_n240), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n237), .B(new_n212), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n234), .B(KEYINPUT13), .Z(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT18), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n250), .B1(new_n239), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  OAI211_X1 g052(.A(KEYINPUT89), .B(new_n250), .C1(new_n239), .C2(new_n251), .ZN(new_n254));
  XNOR2_X1  g053(.A(G113gat), .B(G141gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT11), .ZN(new_n256));
  INV_X1    g055(.A(G169gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G197gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT12), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n247), .A2(new_n253), .A3(new_n262), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n254), .B(new_n261), .C1(new_n246), .C2(new_n252), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(G1gat), .B(G29gat), .Z(new_n267));
  XNOR2_X1  g066(.A(G57gat), .B(G85gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT75), .B(KEYINPUT0), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n269), .B(new_n270), .Z(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G155gat), .B(G162gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G141gat), .ZN(new_n275));
  INV_X1    g074(.A(G148gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT2), .ZN(new_n278));
  NAND2_X1  g077(.A1(G141gat), .A2(G148gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n274), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G155gat), .ZN(new_n282));
  INV_X1    g081(.A(G162gat), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT2), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n273), .A2(new_n277), .A3(new_n284), .A4(new_n279), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT3), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT3), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n281), .A2(new_n285), .A3(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(G127gat), .B(G134gat), .Z(new_n290));
  XNOR2_X1  g089(.A(G113gat), .B(G120gat), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n290), .B1(KEYINPUT1), .B2(new_n291), .ZN(new_n292));
  XOR2_X1   g091(.A(G113gat), .B(G120gat), .Z(new_n293));
  INV_X1    g092(.A(KEYINPUT1), .ZN(new_n294));
  XNOR2_X1  g093(.A(G127gat), .B(G134gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n287), .A2(new_n289), .A3(new_n297), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n292), .A2(new_n296), .A3(new_n281), .A4(new_n285), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT4), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n292), .A2(new_n296), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n281), .A2(new_n285), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n303), .A3(KEYINPUT4), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n298), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G225gat), .A2(G233gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT39), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n297), .A2(new_n286), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n311), .A2(new_n299), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n310), .B1(new_n312), .B2(new_n307), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n272), .B1(new_n309), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n306), .A2(new_n310), .A3(new_n308), .ZN(new_n315));
  AND3_X1   g114(.A1(new_n314), .A2(KEYINPUT40), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT40), .B1(new_n314), .B2(new_n315), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT5), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n305), .A2(KEYINPUT76), .A3(new_n318), .A4(new_n307), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT76), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n298), .A2(new_n304), .A3(new_n307), .A4(new_n301), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n320), .B1(new_n321), .B2(KEYINPUT5), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n299), .B(KEYINPUT4), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n324), .A2(new_n325), .A3(new_n307), .A4(new_n298), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n321), .A2(KEYINPUT73), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT74), .B1(new_n312), .B2(new_n307), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n307), .B1(new_n311), .B2(new_n299), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n318), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n326), .A2(new_n327), .A3(new_n328), .A4(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n271), .B1(new_n323), .B2(new_n332), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n316), .A2(new_n317), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT25), .ZN(new_n335));
  INV_X1    g134(.A(G176gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n257), .A2(new_n336), .A3(KEYINPUT23), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(G169gat), .B2(G176gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n337), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(G183gat), .A2(G190gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT64), .ZN(new_n345));
  NAND3_X1  g144(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n345), .B1(new_n344), .B2(new_n346), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n335), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n337), .A2(new_n340), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT65), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT65), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n353), .A3(new_n340), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n339), .A2(KEYINPUT25), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n356), .B1(new_n346), .B2(new_n344), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n350), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G183gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT27), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT27), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G183gat), .ZN(new_n363));
  INV_X1    g162(.A(G190gat), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n361), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT66), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT28), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(G169gat), .A2(G176gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NOR3_X1   g169(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n343), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n365), .A2(new_n366), .A3(KEYINPUT28), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT29), .B1(new_n359), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G226gat), .ZN(new_n377));
  INV_X1    g176(.A(G233gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G197gat), .B(G204gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT22), .ZN(new_n382));
  XNOR2_X1  g181(.A(G211gat), .B(G218gat), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(G211gat), .ZN(new_n386));
  INV_X1    g185(.A(G218gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n383), .B(new_n381), .C1(KEYINPUT22), .C2(new_n388), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n350), .A2(new_n358), .B1(new_n374), .B2(new_n373), .ZN(new_n391));
  INV_X1    g190(.A(new_n379), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n380), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G8gat), .B(G36gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(G64gat), .B(G92gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT71), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT70), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n401), .B(new_n392), .C1(new_n391), .C2(KEYINPUT29), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n359), .A2(new_n375), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n379), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT29), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n344), .A2(new_n346), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT64), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n408), .A2(new_n347), .A3(new_n341), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n409), .A2(new_n335), .B1(new_n357), .B2(new_n355), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n373), .A2(new_n374), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n406), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n401), .B1(new_n412), .B2(new_n392), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n400), .B(new_n390), .C1(new_n405), .C2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT70), .B1(new_n376), .B2(new_n379), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n416), .A2(new_n402), .A3(new_n404), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n400), .B1(new_n417), .B2(new_n390), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n395), .B(new_n399), .C1(new_n415), .C2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT72), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT30), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n395), .B1(new_n415), .B2(new_n418), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n398), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n421), .B1(new_n419), .B2(new_n420), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n334), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n289), .A2(new_n406), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n390), .ZN(new_n429));
  OR2_X1    g228(.A1(new_n389), .A2(KEYINPUT79), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n389), .A2(KEYINPUT79), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n385), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT3), .B1(new_n432), .B2(new_n406), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n429), .B1(new_n433), .B2(new_n303), .ZN(new_n434));
  NAND2_X1  g233(.A1(G228gat), .A2(G233gat), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n435), .B1(new_n428), .B2(new_n390), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n288), .B1(new_n390), .B2(KEYINPUT29), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n286), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n434), .A2(new_n435), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT81), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(KEYINPUT80), .A2(G22gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(G78gat), .B(G106gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT31), .B(G50gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G22gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n439), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n449), .B2(KEYINPUT81), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n439), .B(new_n448), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n447), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n390), .B1(new_n405), .B2(new_n413), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT71), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n394), .B1(new_n456), .B2(new_n414), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT37), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n398), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n458), .B(new_n395), .C1(new_n415), .C2(new_n418), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT38), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n323), .A2(new_n332), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n272), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n323), .A2(new_n332), .A3(new_n271), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT78), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n468), .B1(new_n464), .B2(new_n465), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n333), .A2(KEYINPUT78), .A3(KEYINPUT6), .ZN(new_n470));
  AND4_X1   g269(.A1(new_n467), .A2(new_n469), .A3(new_n419), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n462), .A2(new_n471), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n399), .A2(KEYINPUT38), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n390), .B1(new_n380), .B2(new_n393), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT82), .ZN(new_n475));
  INV_X1    g274(.A(new_n390), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n416), .A2(new_n476), .A3(new_n402), .A4(new_n404), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT82), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n478), .B(new_n390), .C1(new_n380), .C2(new_n393), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n473), .B1(new_n480), .B2(KEYINPUT37), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n481), .A2(new_n460), .A3(KEYINPUT83), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT83), .B1(new_n481), .B2(new_n460), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n427), .B(new_n454), .C1(new_n472), .C2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT72), .B1(new_n457), .B2(new_n399), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n486), .A2(new_n421), .B1(new_n423), .B2(new_n398), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n333), .A2(KEYINPUT78), .A3(KEYINPUT6), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT78), .B1(new_n333), .B2(KEYINPUT6), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n467), .A2(KEYINPUT77), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT77), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n464), .A2(new_n492), .A3(new_n465), .A4(new_n466), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n490), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n426), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n487), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n443), .A2(new_n450), .B1(new_n452), .B2(new_n447), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT68), .ZN(new_n499));
  NAND2_X1  g298(.A1(G227gat), .A2(G233gat), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n391), .A2(new_n302), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT67), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(new_n403), .B2(new_n297), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n403), .A2(new_n503), .A3(new_n297), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n500), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT32), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n499), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G15gat), .B(G43gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT69), .ZN(new_n511));
  XOR2_X1   g310(.A(G71gat), .B(G99gat), .Z(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT67), .B1(new_n391), .B2(new_n302), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n506), .B1(new_n514), .B2(new_n501), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n515), .A2(G227gat), .A3(G233gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT33), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n516), .A2(KEYINPUT68), .A3(KEYINPUT32), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n509), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n505), .A2(new_n500), .A3(new_n506), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT34), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n516), .B(KEYINPUT32), .C1(new_n517), .C2(new_n513), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n520), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n523), .B1(new_n520), .B2(new_n524), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT36), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n520), .A2(new_n524), .ZN(new_n528));
  INV_X1    g327(.A(new_n523), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT36), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n520), .A2(new_n523), .A3(new_n524), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n485), .A2(new_n498), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n454), .A2(new_n530), .A3(new_n532), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT35), .B1(new_n496), .B2(new_n536), .ZN(new_n537));
  NOR3_X1   g336(.A1(new_n497), .A2(new_n525), .A3(new_n526), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n425), .A2(new_n426), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT35), .B1(new_n490), .B2(new_n467), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT84), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n535), .A2(new_n542), .A3(KEYINPUT84), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n266), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G183gat), .B(G211gat), .Z(new_n548));
  XNOR2_X1  g347(.A(G127gat), .B(G155gat), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n549), .B(KEYINPUT20), .Z(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT90), .ZN(new_n552));
  XNOR2_X1  g351(.A(G57gat), .B(G64gat), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G71gat), .B(G78gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT21), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(KEYINPUT91), .B(KEYINPUT19), .Z(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n561), .A2(new_n562), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n551), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n565), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n567), .A2(new_n550), .A3(new_n563), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n555), .B(new_n556), .Z(new_n569));
  AOI21_X1  g368(.A(new_n212), .B1(KEYINPUT21), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n566), .A2(new_n568), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n571), .B1(new_n566), .B2(new_n568), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n548), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n566), .A2(new_n568), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n570), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n566), .A2(new_n568), .A3(new_n571), .ZN(new_n577));
  INV_X1    g376(.A(new_n548), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  AND2_X1   g379(.A1(G232gat), .A2(G233gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n581), .A2(KEYINPUT41), .ZN(new_n582));
  NAND2_X1  g381(.A1(G99gat), .A2(G106gat), .ZN(new_n583));
  INV_X1    g382(.A(G85gat), .ZN(new_n584));
  INV_X1    g383(.A(G92gat), .ZN(new_n585));
  AOI22_X1  g384(.A1(KEYINPUT8), .A2(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT7), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n587), .B1(new_n584), .B2(new_n585), .ZN(new_n588));
  NAND3_X1  g387(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G99gat), .B(G106gat), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n590), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT92), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n594), .B1(new_n231), .B2(new_n232), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n590), .B(new_n591), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT92), .ZN(new_n597));
  AOI22_X1  g396(.A1(new_n597), .A2(new_n237), .B1(KEYINPUT41), .B2(new_n581), .ZN(new_n598));
  XNOR2_X1  g397(.A(G190gat), .B(G218gat), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n595), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n600), .B1(new_n595), .B2(new_n598), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n582), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n597), .B1(new_n235), .B2(new_n230), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n581), .A2(KEYINPUT41), .ZN(new_n606));
  INV_X1    g405(.A(new_n237), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n606), .B1(new_n607), .B2(new_n594), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n599), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n582), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(new_n610), .A3(new_n601), .ZN(new_n611));
  XOR2_X1   g410(.A(G134gat), .B(G162gat), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n604), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n613), .B1(new_n604), .B2(new_n611), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G230gat), .A2(G233gat), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n597), .A2(KEYINPUT10), .A3(new_n569), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n569), .B(new_n593), .C1(KEYINPUT93), .C2(new_n592), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n592), .A2(KEYINPUT93), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n596), .B1(new_n557), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT94), .B(KEYINPUT10), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n620), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n618), .B1(new_n619), .B2(new_n624), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n620), .A2(new_n622), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n626), .A2(new_n617), .ZN(new_n627));
  XOR2_X1   g426(.A(G120gat), .B(G148gat), .Z(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT95), .ZN(new_n629));
  XNOR2_X1  g428(.A(G176gat), .B(G204gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  OR3_X1    g431(.A1(new_n625), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT96), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n632), .B1(new_n625), .B2(new_n627), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  OAI211_X1 g435(.A(KEYINPUT96), .B(new_n632), .C1(new_n625), .C2(new_n627), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n580), .A2(new_n616), .A3(KEYINPUT97), .A4(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n580), .A2(new_n616), .A3(new_n638), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n547), .B1(new_n640), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(new_n494), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT98), .B(G1gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(G1324gat));
  INV_X1    g447(.A(KEYINPUT42), .ZN(new_n649));
  INV_X1    g448(.A(new_n645), .ZN(new_n650));
  INV_X1    g449(.A(new_n539), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT16), .B(G8gat), .Z(new_n652));
  AND4_X1   g451(.A1(new_n649), .A2(new_n650), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n649), .B1(new_n654), .B2(G8gat), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(G1325gat));
  OAI21_X1  g456(.A(G15gat), .B1(new_n645), .B2(new_n534), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n525), .A2(new_n526), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n660), .A2(G15gat), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n658), .B1(new_n645), .B2(new_n661), .ZN(G1326gat));
  NOR2_X1   g461(.A1(new_n645), .A2(new_n454), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT43), .B(G22gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1327gat));
  INV_X1    g464(.A(new_n580), .ZN(new_n666));
  INV_X1    g465(.A(new_n611), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n610), .B1(new_n609), .B2(new_n601), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n612), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n604), .A2(new_n611), .A3(new_n613), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n666), .A2(new_n671), .A3(new_n638), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT99), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n535), .A2(KEYINPUT84), .A3(new_n542), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT84), .B1(new_n535), .B2(new_n542), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n265), .B(new_n673), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n676), .A2(G29gat), .A3(new_n494), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(KEYINPUT45), .Z(new_n678));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n616), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n680), .B1(new_n674), .B2(new_n675), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n543), .A2(new_n671), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n679), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n494), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n638), .B(KEYINPUT100), .Z(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n687), .A2(new_n266), .A3(new_n580), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n684), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n678), .B1(new_n218), .B2(new_n689), .ZN(G1328gat));
  INV_X1    g489(.A(KEYINPUT101), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n539), .A2(new_n224), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n676), .B2(new_n693), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n547), .A2(KEYINPUT101), .A3(new_n673), .A4(new_n692), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n696), .A2(KEYINPUT46), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n684), .A2(new_n651), .A3(new_n688), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n224), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n696), .A2(KEYINPUT102), .A3(KEYINPUT46), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT102), .B1(new_n696), .B2(KEYINPUT46), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n697), .B(new_n699), .C1(new_n700), .C2(new_n701), .ZN(G1329gat));
  NOR3_X1   g501(.A1(new_n676), .A2(G43gat), .A3(new_n660), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT47), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n704), .A2(KEYINPUT103), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n704), .A2(KEYINPUT103), .ZN(new_n707));
  INV_X1    g506(.A(new_n534), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n681), .A2(new_n708), .A3(new_n683), .A4(new_n688), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G43gat), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n706), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n707), .B1(new_n706), .B2(new_n710), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(G1330gat));
  NAND4_X1  g512(.A1(new_n681), .A2(new_n497), .A3(new_n683), .A4(new_n688), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(G50gat), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n716));
  AOI21_X1  g515(.A(KEYINPUT48), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  OR3_X1    g516(.A1(new_n676), .A2(G50gat), .A3(new_n454), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n715), .B(new_n718), .C1(new_n716), .C2(KEYINPUT48), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(G1331gat));
  NAND2_X1  g521(.A1(new_n580), .A2(new_n616), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n686), .A2(new_n265), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n543), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n685), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g527(.A(new_n539), .B(new_n725), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n729));
  NOR2_X1   g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1333gat));
  NOR3_X1   g530(.A1(new_n725), .A2(G71gat), .A3(new_n660), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n726), .A2(new_n708), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n732), .B1(G71gat), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1334gat));
  NOR2_X1   g535(.A1(new_n725), .A2(new_n454), .ZN(new_n737));
  XNOR2_X1  g536(.A(KEYINPUT106), .B(G78gat), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1335gat));
  NOR2_X1   g538(.A1(new_n265), .A2(new_n580), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n543), .A2(KEYINPUT51), .A3(new_n671), .A4(new_n740), .ZN(new_n741));
  OR2_X1    g540(.A1(new_n741), .A2(KEYINPUT107), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(KEYINPUT107), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n543), .A2(new_n671), .A3(new_n740), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n742), .A2(new_n743), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT108), .ZN(new_n748));
  INV_X1    g547(.A(new_n638), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n685), .A2(new_n584), .A3(new_n749), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n265), .A2(new_n580), .A3(new_n638), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n684), .A2(new_n685), .A3(new_n751), .ZN(new_n752));
  OAI22_X1  g551(.A1(new_n748), .A2(new_n750), .B1(new_n584), .B2(new_n752), .ZN(G1336gat));
  NOR3_X1   g552(.A1(new_n686), .A2(new_n539), .A3(G92gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n747), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n681), .A2(new_n651), .A3(new_n683), .A4(new_n751), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT52), .B1(new_n756), .B2(G92gat), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n754), .B(KEYINPUT109), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n760), .B1(new_n746), .B2(new_n741), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n761), .B1(G92gat), .B2(new_n756), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n758), .B1(new_n759), .B2(new_n762), .ZN(G1337gat));
  NAND3_X1  g562(.A1(new_n684), .A2(new_n708), .A3(new_n751), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G99gat), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n660), .A2(G99gat), .A3(new_n638), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT110), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n748), .B2(new_n767), .ZN(G1338gat));
  NOR3_X1   g567(.A1(new_n686), .A2(G106gat), .A3(new_n454), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n747), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n681), .A2(new_n497), .A3(new_n683), .A4(new_n751), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G106gat), .ZN(new_n772));
  XOR2_X1   g571(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n773));
  NAND3_X1  g572(.A1(new_n770), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n771), .A2(new_n775), .A3(G106gat), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n775), .B1(new_n771), .B2(G106gat), .ZN(new_n777));
  INV_X1    g576(.A(new_n769), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n778), .B1(new_n746), .B2(new_n741), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n774), .B1(new_n780), .B2(new_n781), .ZN(G1339gat));
  INV_X1    g581(.A(new_n625), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n619), .A2(new_n624), .A3(new_n618), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(KEYINPUT54), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n631), .B1(new_n625), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT55), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n785), .A2(KEYINPUT55), .A3(new_n787), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(new_n633), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n791), .B1(new_n263), .B2(new_n264), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n246), .A2(new_n252), .A3(new_n261), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n248), .A2(new_n249), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n233), .B1(new_n236), .B2(new_n238), .ZN(new_n795));
  INV_X1    g594(.A(new_n234), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n794), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n795), .A2(KEYINPUT113), .A3(new_n796), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n260), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n793), .A2(new_n801), .A3(new_n638), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n616), .B1(new_n792), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n261), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n247), .A2(new_n253), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n799), .A2(new_n800), .ZN(new_n806));
  INV_X1    g605(.A(new_n260), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(new_n808), .A3(KEYINPUT114), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n810), .B1(new_n793), .B2(new_n801), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n790), .A2(new_n633), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(new_n788), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n809), .A2(new_n811), .A3(new_n671), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n580), .B1(new_n803), .B2(new_n814), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n723), .A2(new_n265), .A3(new_n749), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n651), .A2(new_n494), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n538), .ZN(new_n821));
  OAI21_X1  g620(.A(G113gat), .B1(new_n821), .B2(new_n266), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n821), .B(KEYINPUT115), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n266), .A2(G113gat), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(G1340gat));
  OR2_X1    g624(.A1(new_n638), .A2(G120gat), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n820), .A2(new_n538), .A3(new_n687), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(new_n828), .A3(G120gat), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n828), .B1(new_n827), .B2(G120gat), .ZN(new_n831));
  OAI22_X1  g630(.A1(new_n823), .A2(new_n826), .B1(new_n830), .B2(new_n831), .ZN(G1341gat));
  NOR2_X1   g631(.A1(new_n821), .A2(new_n666), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(G127gat), .Z(G1342gat));
  NAND2_X1  g633(.A1(new_n820), .A2(new_n671), .ZN(new_n835));
  NAND2_X1  g634(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n538), .A2(new_n836), .ZN(new_n837));
  OR3_X1    g636(.A1(new_n835), .A2(KEYINPUT117), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT117), .B1(new_n835), .B2(new_n837), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n840), .B(new_n841), .ZN(G1343gat));
  NOR2_X1   g641(.A1(new_n708), .A2(new_n454), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n820), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n265), .A2(new_n275), .ZN(new_n846));
  XOR2_X1   g645(.A(new_n846), .B(KEYINPUT118), .Z(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n818), .A2(new_n534), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n850), .B1(new_n817), .B2(new_n454), .ZN(new_n851));
  OAI211_X1 g650(.A(KEYINPUT57), .B(new_n497), .C1(new_n815), .C2(new_n816), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n849), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n853), .A2(new_n265), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n848), .B1(new_n854), .B2(new_n275), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT58), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n857), .B(new_n848), .C1(new_n854), .C2(new_n275), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(G1344gat));
  NOR3_X1   g658(.A1(new_n844), .A2(G148gat), .A3(new_n638), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT119), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n265), .B1(new_n643), .B2(new_n639), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT121), .B1(new_n616), .B2(new_n791), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n671), .A2(new_n813), .A3(new_n865), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n864), .A2(new_n811), .A3(new_n809), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n803), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n863), .B1(new_n868), .B2(new_n666), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n850), .B1(new_n869), .B2(new_n454), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n852), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n849), .B(KEYINPUT120), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n872), .A2(new_n749), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n276), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n862), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n853), .A2(new_n749), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n875), .A3(G148gat), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n874), .A2(new_n862), .A3(new_n875), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n861), .B1(new_n879), .B2(new_n880), .ZN(G1345gat));
  NAND3_X1  g680(.A1(new_n845), .A2(new_n282), .A3(new_n580), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n853), .A2(new_n580), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(new_n282), .ZN(G1346gat));
  NAND2_X1  g683(.A1(new_n843), .A2(new_n283), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT123), .B1(new_n835), .B2(new_n885), .ZN(new_n886));
  OR3_X1    g685(.A1(new_n835), .A2(KEYINPUT123), .A3(new_n885), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n853), .A2(new_n671), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n886), .B(new_n887), .C1(new_n888), .C2(new_n283), .ZN(G1347gat));
  NOR2_X1   g688(.A1(new_n539), .A2(new_n685), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n538), .B(new_n890), .C1(new_n815), .C2(new_n816), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n266), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(new_n257), .ZN(G1348gat));
  OAI21_X1  g692(.A(G176gat), .B1(new_n891), .B2(new_n686), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n749), .A2(new_n336), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n891), .B2(new_n895), .ZN(G1349gat));
  INV_X1    g695(.A(KEYINPUT125), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(KEYINPUT60), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n817), .A2(new_n685), .A3(new_n539), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n900), .A2(KEYINPUT124), .A3(new_n538), .A4(new_n580), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n902), .B1(new_n891), .B2(new_n666), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n360), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n891), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n906), .A2(new_n361), .A3(new_n363), .A4(new_n580), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n897), .A2(KEYINPUT60), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n899), .B1(new_n905), .B2(new_n910), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n904), .A2(new_n909), .A3(new_n898), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n911), .A2(new_n912), .ZN(G1350gat));
  NAND2_X1  g712(.A1(new_n906), .A2(new_n671), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(new_n915), .A3(G190gat), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n915), .B1(new_n914), .B2(G190gat), .ZN(new_n918));
  OAI22_X1  g717(.A1(new_n917), .A2(new_n918), .B1(G190gat), .B2(new_n914), .ZN(G1351gat));
  NAND2_X1  g718(.A1(new_n900), .A2(new_n843), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(G197gat), .B1(new_n921), .B2(new_n265), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n534), .A2(new_n890), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n923), .B1(new_n870), .B2(new_n852), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n266), .A2(new_n259), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(G1352gat));
  NOR3_X1   g725(.A1(new_n920), .A2(G204gat), .A3(new_n638), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT62), .ZN(new_n928));
  INV_X1    g727(.A(new_n924), .ZN(new_n929));
  OAI21_X1  g728(.A(G204gat), .B1(new_n929), .B2(new_n686), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1353gat));
  INV_X1    g730(.A(new_n923), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n868), .A2(new_n666), .ZN(new_n933));
  INV_X1    g732(.A(new_n863), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT57), .B1(new_n935), .B2(new_n497), .ZN(new_n936));
  INV_X1    g735(.A(new_n852), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n580), .B(new_n932), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n938), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n938), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n938), .A2(G211gat), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT63), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n941), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n921), .A2(new_n386), .A3(new_n580), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1354gat));
  AND2_X1   g747(.A1(new_n924), .A2(KEYINPUT127), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n671), .B1(new_n924), .B2(KEYINPUT127), .ZN(new_n950));
  OAI21_X1  g749(.A(G218gat), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n921), .A2(new_n387), .A3(new_n671), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1355gat));
endmodule


