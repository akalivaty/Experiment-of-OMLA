//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 0 0 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n789, new_n790, new_n791, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010, new_n1011;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT78), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  AND2_X1   g004(.A1(G226gat), .A2(G233gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT29), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(KEYINPUT68), .ZN(new_n211));
  NOR2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT23), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(KEYINPUT25), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G169gat), .ZN(new_n215));
  INV_X1    g014(.A(G176gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT66), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n220));
  NOR3_X1   g019(.A1(new_n212), .A2(new_n220), .A3(KEYINPUT23), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT24), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT24), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n226), .A2(G183gat), .A3(G190gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n223), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  NOR3_X1   g027(.A1(new_n214), .A2(new_n222), .A3(new_n228), .ZN(new_n229));
  AND2_X1   g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n230), .B1(KEYINPUT23), .B2(new_n212), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(new_n219), .B2(new_n221), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT67), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT67), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n234), .B(new_n231), .C1(new_n219), .C2(new_n221), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n223), .B(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n225), .A2(new_n227), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n233), .A2(new_n235), .A3(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n241));
  AOI21_X1  g040(.A(new_n229), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT26), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n212), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n210), .B1(new_n212), .B2(new_n243), .ZN(new_n246));
  OAI211_X1 g045(.A(KEYINPUT69), .B(new_n224), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G183gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT27), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT27), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G183gat), .ZN(new_n251));
  INV_X1    g050(.A(G190gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  OR2_X1    g052(.A1(new_n253), .A2(KEYINPUT28), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(KEYINPUT28), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n247), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n217), .A2(KEYINPUT26), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n257), .A2(new_n210), .A3(new_n244), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT69), .B1(new_n258), .B2(new_n224), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n209), .B1(new_n242), .B2(new_n260), .ZN(new_n261));
  OR2_X1    g060(.A1(new_n256), .A2(new_n259), .ZN(new_n262));
  INV_X1    g061(.A(new_n241), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n232), .A2(KEYINPUT67), .B1(new_n238), .B2(new_n237), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n263), .B1(new_n264), .B2(new_n235), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n262), .B(new_n207), .C1(new_n265), .C2(new_n229), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G197gat), .B(G204gat), .ZN(new_n268));
  AND2_X1   g067(.A1(G211gat), .A2(G218gat), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n268), .B1(KEYINPUT22), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G211gat), .B(G218gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT76), .ZN(new_n274));
  INV_X1    g073(.A(new_n272), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n261), .A2(new_n275), .A3(new_n266), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n273), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n267), .A2(KEYINPUT76), .A3(new_n272), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n277), .A2(KEYINPUT77), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT77), .B1(new_n277), .B2(new_n278), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n205), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G225gat), .A2(G233gat), .ZN(new_n282));
  INV_X1    g081(.A(G113gat), .ZN(new_n283));
  INV_X1    g082(.A(G120gat), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT1), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G127gat), .B(G134gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT70), .B(G120gat), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n285), .B(new_n286), .C1(new_n287), .C2(new_n283), .ZN(new_n288));
  AND2_X1   g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(G155gat), .A2(G162gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G141gat), .B(G148gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT2), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n293), .B1(G155gat), .B2(G162gat), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n291), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G134gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G127gat), .ZN(new_n297));
  INV_X1    g096(.A(G127gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G134gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n283), .A2(new_n284), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT1), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n302), .B1(G113gat), .B2(G120gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n300), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G141gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G148gat), .ZN(new_n306));
  INV_X1    g105(.A(G148gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G141gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G155gat), .B(G162gat), .ZN(new_n310));
  INV_X1    g109(.A(G155gat), .ZN(new_n311));
  INV_X1    g110(.A(G162gat), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT2), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n309), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n288), .A2(new_n295), .A3(new_n304), .A4(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n315), .B(KEYINPUT4), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n309), .A2(new_n310), .A3(new_n313), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n310), .B1(new_n313), .B2(new_n309), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT3), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n295), .A2(new_n314), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n288), .A2(new_n304), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT79), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n295), .A2(new_n314), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n326), .A2(KEYINPUT3), .B1(new_n304), .B2(new_n288), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT79), .B1(new_n327), .B2(new_n321), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n282), .B(new_n316), .C1(new_n325), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n322), .A2(new_n326), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n315), .ZN(new_n331));
  INV_X1    g130(.A(new_n282), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT5), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(G1gat), .B(G29gat), .Z(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(KEYINPUT0), .ZN(new_n338));
  XNOR2_X1  g137(.A(G57gat), .B(G85gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n300), .A2(new_n303), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT70), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n342), .A2(G120gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n284), .A2(KEYINPUT70), .ZN(new_n344));
  OAI21_X1  g143(.A(G113gat), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n285), .B1(new_n283), .B2(new_n284), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n341), .A2(new_n345), .B1(new_n346), .B2(new_n300), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n347), .A2(KEYINPUT4), .A3(new_n295), .A4(new_n314), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n315), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n323), .A2(new_n324), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n327), .A2(KEYINPUT79), .A3(new_n321), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT5), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(new_n355), .A3(new_n282), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n336), .A2(new_n340), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT6), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n340), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n329), .A2(KEYINPUT5), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n334), .B1(new_n354), .B2(new_n282), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n340), .B1(new_n336), .B2(new_n356), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT6), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n205), .B1(new_n277), .B2(new_n278), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT30), .ZN(new_n369));
  INV_X1    g168(.A(new_n205), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n276), .A2(new_n274), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n275), .B1(new_n261), .B2(new_n266), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n278), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n370), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT30), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n281), .A2(new_n367), .A3(new_n369), .A4(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(G228gat), .A2(G233gat), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n320), .B1(new_n272), .B2(KEYINPUT29), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(new_n326), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n379), .B1(new_n381), .B2(KEYINPUT81), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n321), .A2(new_n208), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n272), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n381), .B(new_n384), .C1(KEYINPUT81), .C2(new_n379), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AND2_X1   g187(.A1(KEYINPUT83), .A2(G22gat), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  XOR2_X1   g189(.A(G78gat), .B(G106gat), .Z(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT31), .B(G50gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n393), .B1(new_n388), .B2(new_n389), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  AND3_X1   g194(.A1(new_n386), .A2(KEYINPUT82), .A3(new_n387), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT82), .B1(new_n386), .B2(new_n387), .ZN(new_n397));
  INV_X1    g196(.A(G22gat), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n398), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n393), .B(KEYINPUT80), .Z(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n395), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n378), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT36), .ZN(new_n406));
  AND2_X1   g205(.A1(G227gat), .A2(G233gat), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n347), .B1(new_n242), .B2(new_n260), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n262), .B(new_n322), .C1(new_n265), .C2(new_n229), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n410), .A2(KEYINPUT75), .A3(KEYINPUT34), .ZN(new_n411));
  XOR2_X1   g210(.A(KEYINPUT75), .B(KEYINPUT34), .Z(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n411), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G15gat), .B(G43gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(KEYINPUT72), .ZN(new_n416));
  XNOR2_X1  g215(.A(G71gat), .B(G99gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n408), .A2(new_n407), .A3(new_n409), .ZN(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT71), .B(KEYINPUT33), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT73), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n420), .A2(KEYINPUT32), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n423), .B1(new_n422), .B2(new_n424), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OR2_X1    g226(.A1(new_n419), .A2(new_n421), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n420), .A2(KEYINPUT32), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT74), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n420), .A2(KEYINPUT74), .A3(KEYINPUT32), .A4(new_n428), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n414), .B1(new_n427), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n420), .A2(new_n421), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n424), .A2(new_n435), .A3(new_n418), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT73), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n437), .A2(new_n433), .A3(new_n438), .A4(new_n414), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n406), .B1(new_n434), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n437), .A2(new_n433), .A3(new_n438), .ZN(new_n442));
  INV_X1    g241(.A(new_n414), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n444), .A2(KEYINPUT36), .A3(new_n439), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT38), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT37), .B1(new_n279), .B2(new_n280), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n277), .A2(new_n278), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT37), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n370), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n447), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT85), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n363), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n365), .A2(KEYINPUT85), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n359), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT86), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n359), .A2(new_n454), .A3(KEYINPUT86), .A4(new_n455), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(new_n366), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n450), .B1(new_n373), .B2(new_n374), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n205), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n372), .A2(KEYINPUT87), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n276), .B1(new_n372), .B2(KEYINPUT87), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT37), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(new_n447), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n375), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n452), .A2(new_n460), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n336), .A2(new_n356), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT85), .B1(new_n469), .B2(new_n360), .ZN(new_n470));
  AOI211_X1 g269(.A(new_n453), .B(new_n340), .C1(new_n336), .C2(new_n356), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n354), .A2(new_n282), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT39), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n360), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n331), .A2(new_n332), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT84), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n478), .B1(new_n477), .B2(new_n476), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n475), .B(KEYINPUT40), .C1(new_n473), .C2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n475), .B1(new_n473), .B2(new_n479), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT40), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n472), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n377), .A2(new_n369), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT77), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n486), .B1(new_n373), .B2(new_n374), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n277), .A2(KEYINPUT77), .A3(new_n278), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n370), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n484), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n403), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n405), .B(new_n446), .C1(new_n468), .C2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n444), .A2(new_n403), .A3(new_n439), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n281), .A2(new_n369), .A3(new_n377), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n459), .A2(new_n366), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT86), .B1(new_n472), .B2(new_n359), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(KEYINPUT35), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT35), .B1(new_n493), .B2(new_n378), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n492), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G113gat), .B(G141gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G169gat), .B(G197gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(new_n508), .B(KEYINPUT12), .Z(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G229gat), .A2(G233gat), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G43gat), .B(G50gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT15), .ZN(new_n514));
  XNOR2_X1  g313(.A(KEYINPUT91), .B(G43gat), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n515), .A2(G50gat), .ZN(new_n516));
  XOR2_X1   g315(.A(KEYINPUT92), .B(G50gat), .Z(new_n517));
  INV_X1    g316(.A(G43gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT15), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(KEYINPUT90), .B(G29gat), .Z(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G36gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(G29gat), .A2(G36gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT89), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT89), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(G29gat), .B2(G36gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n524), .A2(new_n526), .A3(KEYINPUT14), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n526), .A2(KEYINPUT14), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n522), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n514), .B1(new_n520), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n529), .A2(new_n514), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G15gat), .B(G22gat), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT16), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n533), .B1(new_n534), .B2(G1gat), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(G1gat), .B2(new_n533), .ZN(new_n536));
  INV_X1    g335(.A(G8gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n532), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT17), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n530), .A2(new_n540), .A3(new_n531), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT93), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n530), .A2(new_n531), .A3(KEYINPUT93), .A4(new_n540), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n536), .B(G8gat), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n546), .B1(new_n532), .B2(KEYINPUT17), .ZN(new_n547));
  AOI211_X1 g346(.A(new_n512), .B(new_n539), .C1(new_n545), .C2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n510), .B1(new_n548), .B2(KEYINPUT18), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n529), .A2(new_n514), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n522), .A2(new_n527), .A3(new_n528), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT15), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n515), .A2(G50gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT92), .B(G50gat), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n554), .A2(G43gat), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n552), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n550), .B1(new_n557), .B2(new_n514), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT93), .B1(new_n558), .B2(new_n540), .ZN(new_n559));
  INV_X1    g358(.A(new_n544), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n547), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n546), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n561), .A2(KEYINPUT18), .A3(new_n511), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n532), .A2(new_n538), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT94), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n511), .B(KEYINPUT13), .Z(new_n567));
  NAND3_X1  g366(.A1(new_n532), .A2(KEYINPUT94), .A3(new_n538), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT96), .B1(new_n549), .B2(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n563), .A2(new_n569), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT96), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n561), .A2(new_n511), .A3(new_n562), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT18), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n509), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n572), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n574), .A2(new_n575), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n579), .B1(new_n570), .B2(KEYINPUT95), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT95), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n581), .B1(new_n563), .B2(new_n569), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n509), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(G57gat), .B(G64gat), .Z(new_n585));
  INV_X1    g384(.A(KEYINPUT9), .ZN(new_n586));
  INV_X1    g385(.A(G71gat), .ZN(new_n587));
  INV_X1    g386(.A(G78gat), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n585), .A2(KEYINPUT97), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n587), .A2(new_n588), .ZN(new_n592));
  NOR2_X1   g391(.A1(G71gat), .A2(G78gat), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n590), .B(new_n591), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G57gat), .B(G64gat), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT97), .ZN(new_n596));
  OAI22_X1  g395(.A1(new_n595), .A2(new_n596), .B1(new_n592), .B2(new_n593), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(new_n589), .A3(new_n585), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n599), .A2(KEYINPUT21), .ZN(new_n600));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(G127gat), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT21), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n597), .B(new_n590), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n538), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n603), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(G155gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(G183gat), .B(G211gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n607), .B(new_n611), .ZN(new_n612));
  AND2_X1   g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n613), .A2(KEYINPUT41), .ZN(new_n614));
  XNOR2_X1  g413(.A(G134gat), .B(G162gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G99gat), .B(G106gat), .Z(new_n618));
  OR2_X1    g417(.A1(KEYINPUT99), .A2(G92gat), .ZN(new_n619));
  INV_X1    g418(.A(G85gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(KEYINPUT99), .A2(G92gat), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G85gat), .A2(G92gat), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT7), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(KEYINPUT98), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G99gat), .A2(G106gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT8), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n622), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT7), .B1(new_n623), .B2(KEYINPUT98), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT98), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n630), .B1(G85gat), .B2(G92gat), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n618), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n628), .A2(new_n632), .A3(new_n618), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n558), .A2(new_n636), .B1(KEYINPUT41), .B2(new_n613), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n636), .B1(new_n532), .B2(KEYINPUT17), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n545), .A2(new_n638), .A3(KEYINPUT100), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT100), .B1(new_n545), .B2(new_n638), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n637), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(G190gat), .B(G218gat), .Z(new_n643));
  AND2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n617), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n642), .A2(new_n643), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n642), .A2(new_n643), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n616), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n612), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n605), .B1(new_n635), .B2(new_n634), .ZN(new_n652));
  INV_X1    g451(.A(new_n628), .ZN(new_n653));
  INV_X1    g452(.A(new_n618), .ZN(new_n654));
  INV_X1    g453(.A(new_n632), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n599), .A2(new_n656), .A3(new_n633), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n652), .A2(new_n657), .A3(KEYINPUT101), .ZN(new_n658));
  INV_X1    g457(.A(G230gat), .ZN(new_n659));
  INV_X1    g458(.A(G233gat), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n605), .B(new_n662), .C1(new_n635), .C2(new_n634), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n658), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G120gat), .B(G148gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(G176gat), .B(G204gat), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n665), .B(new_n666), .Z(new_n667));
  INV_X1    g466(.A(KEYINPUT10), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n657), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n658), .A2(new_n663), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n669), .B1(new_n670), .B2(new_n668), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n664), .B(new_n667), .C1(new_n671), .C2(new_n661), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT102), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT10), .B1(new_n658), .B2(new_n663), .ZN(new_n674));
  OAI22_X1  g473(.A1(new_n674), .A2(new_n669), .B1(new_n659), .B2(new_n660), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n675), .A2(new_n676), .A3(new_n664), .A4(new_n667), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n667), .B1(new_n675), .B2(new_n664), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(KEYINPUT103), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n678), .A2(new_n683), .A3(new_n680), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n651), .A2(new_n685), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n503), .A2(new_n584), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n367), .B(KEYINPUT104), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g489(.A1(new_n687), .A2(new_n494), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(new_n537), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT105), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT16), .B(G8gat), .Z(new_n694));
  NAND2_X1  g493(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT42), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n696), .ZN(G1325gat));
  INV_X1    g496(.A(G15gat), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n434), .A2(new_n440), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n687), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n444), .A2(KEYINPUT36), .A3(new_n439), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT36), .B1(new_n444), .B2(new_n439), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n441), .A2(KEYINPUT106), .A3(new_n445), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n687), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n700), .B1(new_n708), .B2(new_n698), .ZN(G1326gat));
  NAND2_X1  g508(.A1(new_n687), .A2(new_n404), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT107), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT43), .B(G22gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  AOI21_X1  g512(.A(new_n650), .B1(new_n492), .B2(new_n502), .ZN(new_n714));
  INV_X1    g513(.A(new_n584), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n715), .A2(new_n685), .A3(new_n612), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n688), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n717), .A2(new_n521), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n646), .A2(new_n649), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n503), .A2(KEYINPUT44), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n450), .B1(new_n487), .B2(new_n488), .ZN(new_n724));
  OAI21_X1  g523(.A(KEYINPUT38), .B1(new_n724), .B2(new_n462), .ZN(new_n725));
  INV_X1    g524(.A(new_n466), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n368), .B1(new_n726), .B2(new_n451), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n498), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n404), .B1(new_n494), .B2(new_n484), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n730), .A2(new_n704), .A3(new_n405), .A4(new_n705), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n650), .B1(new_n731), .B2(new_n502), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n723), .B(new_n716), .C1(KEYINPUT44), .C2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n521), .B1(new_n733), .B2(new_n718), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n721), .A2(new_n734), .ZN(G1328gat));
  INV_X1    g534(.A(new_n494), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n717), .A2(G36gat), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT46), .ZN(new_n738));
  OAI21_X1  g537(.A(G36gat), .B1(new_n733), .B2(new_n736), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(G1329gat));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n741));
  INV_X1    g540(.A(new_n378), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n444), .A2(new_n403), .A3(new_n439), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI22_X1  g543(.A1(new_n744), .A2(KEYINPUT35), .B1(new_n495), .B2(new_n499), .ZN(new_n745));
  AOI22_X1  g544(.A1(new_n728), .A2(new_n729), .B1(new_n378), .B2(new_n404), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n745), .B1(new_n706), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n741), .B1(new_n747), .B2(new_n650), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n748), .A2(new_n707), .A3(new_n716), .A4(new_n723), .ZN(new_n749));
  INV_X1    g548(.A(new_n515), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n717), .ZN(new_n752));
  INV_X1    g551(.A(new_n699), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(new_n750), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT47), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n755), .A2(KEYINPUT47), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n515), .B1(new_n749), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n731), .A2(new_n502), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT44), .B1(new_n762), .B2(new_n722), .ZN(new_n763));
  AOI211_X1 g562(.A(new_n741), .B(new_n650), .C1(new_n492), .C2(new_n502), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n765), .A2(KEYINPUT109), .A3(new_n707), .A4(new_n716), .ZN(new_n766));
  AOI211_X1 g565(.A(KEYINPUT110), .B(new_n759), .C1(new_n761), .C2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n760), .B1(new_n733), .B2(new_n706), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n766), .A2(new_n769), .A3(new_n750), .ZN(new_n770));
  INV_X1    g569(.A(new_n759), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n768), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n758), .B1(new_n767), .B2(new_n772), .ZN(G1330gat));
  OR2_X1    g572(.A1(new_n717), .A2(KEYINPUT111), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n403), .B1(new_n717), .B2(KEYINPUT111), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n517), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n733), .A2(new_n403), .A3(new_n554), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT48), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(G1331gat));
  INV_X1    g579(.A(new_n685), .ZN(new_n781));
  NOR4_X1   g580(.A1(new_n747), .A2(new_n584), .A3(new_n651), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n688), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n494), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n786));
  XOR2_X1   g585(.A(KEYINPUT49), .B(G64gat), .Z(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n785), .B2(new_n787), .ZN(G1333gat));
  AOI21_X1  g587(.A(new_n587), .B1(new_n782), .B2(new_n707), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n753), .A2(G71gat), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n789), .B1(new_n782), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g591(.A1(new_n782), .A2(new_n404), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g593(.A1(new_n612), .A2(new_n584), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(new_n781), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n723), .B(new_n797), .C1(KEYINPUT44), .C2(new_n732), .ZN(new_n798));
  OAI21_X1  g597(.A(G85gat), .B1(new_n798), .B2(new_n718), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n732), .A2(new_n795), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n800), .A2(KEYINPUT51), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(KEYINPUT51), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n685), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n688), .A2(new_n620), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n799), .B1(new_n803), .B2(new_n804), .ZN(G1336gat));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n619), .A2(new_n621), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n807), .B1(new_n798), .B2(new_n736), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n736), .A2(G92gat), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n806), .B(new_n808), .C1(new_n803), .C2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812));
  NOR2_X1   g611(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n800), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n813), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n732), .B2(new_n795), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n685), .B(new_n809), .C1(new_n814), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n808), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n812), .B1(new_n818), .B2(KEYINPUT52), .ZN(new_n819));
  AOI211_X1 g618(.A(KEYINPUT113), .B(new_n806), .C1(new_n817), .C2(new_n808), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n811), .B1(new_n819), .B2(new_n820), .ZN(G1337gat));
  OAI21_X1  g620(.A(G99gat), .B1(new_n798), .B2(new_n706), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n753), .A2(G99gat), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(new_n803), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n824), .B(new_n825), .ZN(G1338gat));
  NAND3_X1  g625(.A1(new_n765), .A2(new_n404), .A3(new_n797), .ZN(new_n827));
  XNOR2_X1  g626(.A(KEYINPUT115), .B(G106gat), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n781), .A2(G106gat), .A3(new_n403), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n801), .A2(new_n802), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n814), .A2(new_n816), .ZN(new_n834));
  AOI22_X1  g633(.A1(new_n834), .A2(new_n831), .B1(new_n827), .B2(new_n828), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n835), .B2(new_n830), .ZN(G1339gat));
  NOR3_X1   g635(.A1(new_n651), .A2(new_n685), .A3(new_n584), .ZN(new_n837));
  INV_X1    g636(.A(new_n561), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n512), .B1(new_n838), .B2(new_n539), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n566), .A2(new_n568), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n567), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n508), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n549), .A2(new_n570), .A3(KEYINPUT96), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n573), .B1(new_n572), .B2(new_n576), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n845), .B1(new_n682), .B2(new_n684), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n670), .A2(new_n668), .ZN(new_n848));
  INV_X1    g647(.A(new_n669), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n849), .A3(new_n661), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n850), .A2(new_n675), .A3(KEYINPUT54), .ZN(new_n851));
  INV_X1    g650(.A(new_n667), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n852), .B1(new_n675), .B2(KEYINPUT54), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n847), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n671), .A2(new_n661), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n667), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n850), .A2(new_n675), .A3(KEYINPUT54), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(KEYINPUT55), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n854), .A2(new_n859), .A3(new_n678), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n860), .B1(new_n578), .B2(new_n583), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n650), .B1(new_n846), .B2(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n650), .A2(new_n845), .A3(new_n860), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n612), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n837), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n867), .A2(new_n718), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n868), .A2(new_n495), .ZN(new_n869));
  AOI21_X1  g668(.A(G113gat), .B1(new_n869), .B2(new_n584), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n718), .A2(new_n494), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n699), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT116), .B1(new_n867), .B2(new_n404), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n854), .A2(new_n859), .A3(new_n678), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n584), .A2(new_n874), .ZN(new_n875));
  AOI22_X1  g674(.A1(new_n571), .A2(new_n577), .B1(new_n508), .B2(new_n841), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n683), .B1(new_n678), .B2(new_n680), .ZN(new_n877));
  AOI211_X1 g676(.A(KEYINPUT103), .B(new_n679), .C1(new_n673), .C2(new_n677), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n722), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n866), .B1(new_n880), .B2(new_n863), .ZN(new_n881));
  INV_X1    g680(.A(new_n837), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n883), .A2(new_n884), .A3(new_n403), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n872), .B1(new_n873), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n715), .A2(new_n283), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n870), .B1(new_n886), .B2(new_n887), .ZN(G1340gat));
  INV_X1    g687(.A(new_n886), .ZN(new_n889));
  OAI21_X1  g688(.A(G120gat), .B1(new_n889), .B2(new_n781), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n869), .A2(new_n287), .A3(new_n685), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1341gat));
  OAI21_X1  g691(.A(G127gat), .B1(new_n889), .B2(new_n866), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n869), .A2(new_n298), .A3(new_n612), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1342gat));
  NAND4_X1  g694(.A1(new_n868), .A2(new_n296), .A3(new_n495), .A4(new_n722), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT56), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n296), .B1(new_n886), .B2(new_n722), .ZN(new_n898));
  OAI21_X1  g697(.A(KEYINPUT117), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT56), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n896), .B(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n898), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT117), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n899), .A2(new_n904), .ZN(G1343gat));
  AND2_X1   g704(.A1(new_n706), .A2(new_n871), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n883), .A2(new_n404), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT57), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n403), .B1(new_n881), .B2(new_n882), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(KEYINPUT57), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n906), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(G141gat), .B1(new_n912), .B2(new_n715), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n914), .A2(KEYINPUT58), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n706), .A2(new_n404), .ZN(new_n916));
  NOR4_X1   g715(.A1(new_n867), .A2(new_n916), .A3(new_n494), .A4(new_n718), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n715), .A2(G141gat), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n917), .A2(new_n918), .B1(new_n914), .B2(KEYINPUT58), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n913), .A2(new_n915), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n915), .B1(new_n913), .B2(new_n919), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n920), .A2(new_n921), .ZN(G1344gat));
  NAND3_X1  g721(.A1(new_n917), .A2(new_n307), .A3(new_n685), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n923), .B(KEYINPUT119), .Z(new_n924));
  NOR2_X1   g723(.A1(new_n912), .A2(new_n781), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n925), .A2(KEYINPUT59), .A3(new_n307), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT59), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT120), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n928), .B1(new_n910), .B2(KEYINPUT57), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n908), .B1(new_n867), .B2(new_n403), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n907), .A2(new_n928), .A3(new_n908), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n931), .A2(new_n685), .A3(new_n906), .A4(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n927), .B1(new_n933), .B2(G148gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n924), .B1(new_n926), .B2(new_n934), .ZN(G1345gat));
  OAI21_X1  g734(.A(G155gat), .B1(new_n912), .B2(new_n866), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n917), .A2(new_n311), .A3(new_n612), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1346gat));
  NAND3_X1  g737(.A1(new_n917), .A2(new_n312), .A3(new_n722), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT121), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n940), .B1(new_n912), .B2(new_n650), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G162gat), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n912), .A2(new_n940), .A3(new_n650), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n939), .B1(new_n942), .B2(new_n943), .ZN(G1347gat));
  NOR4_X1   g743(.A1(new_n867), .A2(new_n736), .A3(new_n493), .A4(new_n688), .ZN(new_n945));
  AOI21_X1  g744(.A(G169gat), .B1(new_n945), .B2(new_n584), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n688), .A2(new_n736), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(new_n699), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n948), .B1(new_n873), .B2(new_n885), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n715), .A2(new_n215), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(G1348gat));
  AOI21_X1  g750(.A(new_n216), .B1(new_n949), .B2(new_n685), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n945), .A2(new_n216), .A3(new_n685), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n952), .A2(new_n953), .ZN(G1349gat));
  AOI21_X1  g753(.A(new_n248), .B1(new_n949), .B2(new_n612), .ZN(new_n955));
  AND4_X1   g754(.A1(new_n249), .A2(new_n945), .A3(new_n251), .A4(new_n612), .ZN(new_n956));
  OR3_X1    g755(.A1(new_n955), .A2(new_n956), .A3(KEYINPUT60), .ZN(new_n957));
  OAI21_X1  g756(.A(KEYINPUT60), .B1(new_n955), .B2(new_n956), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1350gat));
  NAND2_X1  g758(.A1(new_n873), .A2(new_n885), .ZN(new_n960));
  INV_X1    g759(.A(new_n948), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n960), .A2(new_n722), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(G190gat), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT122), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n962), .A2(KEYINPUT122), .A3(G190gat), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n965), .A2(KEYINPUT61), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(KEYINPUT122), .B1(new_n962), .B2(G190gat), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n650), .A2(G190gat), .ZN(new_n970));
  AOI22_X1  g769(.A1(new_n968), .A2(new_n969), .B1(new_n945), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n967), .A2(new_n971), .ZN(G1351gat));
  NOR4_X1   g771(.A1(new_n867), .A2(new_n916), .A3(new_n736), .A4(new_n688), .ZN(new_n973));
  AOI21_X1  g772(.A(G197gat), .B1(new_n973), .B2(new_n584), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n931), .A2(new_n932), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT123), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n931), .A2(KEYINPUT123), .A3(new_n932), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n584), .A2(G197gat), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n706), .A2(new_n947), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT124), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n706), .A2(KEYINPUT124), .A3(new_n947), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n985), .A2(KEYINPUT125), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(KEYINPUT125), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n980), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n974), .B1(new_n979), .B2(new_n988), .ZN(G1352gat));
  AOI21_X1  g788(.A(new_n781), .B1(new_n986), .B2(new_n987), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n977), .A2(new_n990), .A3(new_n978), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n991), .A2(G204gat), .ZN(new_n992));
  INV_X1    g791(.A(G204gat), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n973), .A2(new_n993), .A3(new_n685), .ZN(new_n994));
  XOR2_X1   g793(.A(new_n994), .B(KEYINPUT62), .Z(new_n995));
  NAND2_X1  g794(.A1(new_n992), .A2(new_n995), .ZN(G1353gat));
  AOI21_X1  g795(.A(new_n866), .B1(new_n983), .B2(new_n984), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n931), .A2(new_n932), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n998), .A2(G211gat), .ZN(new_n999));
  NOR2_X1   g798(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g800(.A(new_n998), .B(G211gat), .C1(KEYINPUT126), .C2(KEYINPUT63), .ZN(new_n1002));
  NAND2_X1  g801(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g803(.A(G211gat), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n973), .A2(new_n1005), .A3(new_n612), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1004), .A2(new_n1006), .ZN(G1354gat));
  AOI21_X1  g806(.A(G218gat), .B1(new_n973), .B2(new_n722), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n722), .A2(G218gat), .ZN(new_n1009));
  XNOR2_X1  g808(.A(new_n1009), .B(KEYINPUT127), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n1010), .B1(new_n986), .B2(new_n987), .ZN(new_n1011));
  AOI21_X1  g810(.A(new_n1008), .B1(new_n979), .B2(new_n1011), .ZN(G1355gat));
endmodule


