//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT22), .B(G137), .ZN(new_n191));
  INV_X1    g005(.A(G221), .ZN(new_n192));
  INV_X1    g006(.A(G234), .ZN(new_n193));
  NOR3_X1   g007(.A1(new_n192), .A2(new_n193), .A3(G953), .ZN(new_n194));
  XOR2_X1   g008(.A(new_n191), .B(new_n194), .Z(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT67), .B(G119), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT75), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G119), .ZN(new_n200));
  AOI22_X1  g014(.A1(new_n197), .A2(G128), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G119), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT67), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT67), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G119), .ZN(new_n205));
  AND4_X1   g019(.A1(new_n198), .A2(new_n203), .A3(new_n205), .A4(G128), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT76), .B1(new_n201), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT24), .B(G110), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n203), .A2(new_n205), .A3(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n200), .A2(new_n198), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n197), .A2(new_n198), .A3(G128), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT76), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n207), .A2(new_n208), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT77), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n217), .B1(new_n197), .B2(G128), .ZN(new_n218));
  INV_X1    g032(.A(G110), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n199), .A2(KEYINPUT23), .A3(G119), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n218), .A2(new_n219), .A3(new_n209), .A4(new_n220), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n215), .A2(new_n216), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n216), .B1(new_n215), .B2(new_n221), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT16), .ZN(new_n224));
  INV_X1    g038(.A(G140), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(new_n225), .A3(G125), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(G125), .ZN(new_n227));
  INV_X1    g041(.A(G125), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G140), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g044(.A(G146), .B(new_n226), .C1(new_n230), .C2(new_n224), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(G146), .B2(new_n230), .ZN(new_n232));
  NOR3_X1   g046(.A1(new_n222), .A2(new_n223), .A3(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n226), .B1(new_n230), .B2(new_n224), .ZN(new_n234));
  INV_X1    g048(.A(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n231), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n218), .A2(new_n209), .A3(new_n220), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n237), .B1(new_n238), .B2(new_n219), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n208), .B1(new_n207), .B2(new_n214), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n196), .B1(new_n233), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n223), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n215), .A2(new_n216), .A3(new_n221), .ZN(new_n244));
  INV_X1    g058(.A(new_n232), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n241), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(new_n195), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n242), .A2(new_n188), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT25), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n242), .A2(new_n248), .A3(KEYINPUT25), .A4(new_n188), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n190), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n242), .A2(new_n248), .ZN(new_n254));
  NOR3_X1   g068(.A1(new_n254), .A2(G902), .A3(new_n189), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(G214), .B1(G237), .B2(G902), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n203), .A2(new_n205), .A3(G116), .ZN(new_n258));
  INV_X1    g072(.A(G116), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G119), .ZN(new_n260));
  INV_X1    g074(.A(G113), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT2), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT2), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G113), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n258), .A2(new_n260), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT68), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n258), .A2(new_n265), .A3(KEYINPUT68), .A4(new_n260), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G104), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT3), .B1(new_n271), .B2(G107), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT3), .ZN(new_n273));
  INV_X1    g087(.A(G107), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(new_n274), .A3(G104), .ZN(new_n275));
  INV_X1    g089(.A(G101), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n271), .A2(G107), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n272), .A2(new_n275), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n271), .A2(G107), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n274), .A2(G104), .ZN(new_n280));
  OAI21_X1  g094(.A(G101), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT5), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n203), .A2(new_n205), .A3(new_n284), .A4(G116), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n285), .A2(G113), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n258), .A2(KEYINPUT5), .A3(new_n260), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n270), .A2(new_n283), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n258), .A2(new_n260), .ZN(new_n290));
  INV_X1    g104(.A(new_n265), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n268), .A2(new_n269), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n272), .A2(new_n275), .A3(new_n277), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT4), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n294), .A3(G101), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n293), .A2(G101), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n278), .A2(KEYINPUT4), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n289), .B1(new_n292), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(G110), .B(G122), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n289), .B(new_n300), .C1(new_n292), .C2(new_n298), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n303), .A3(KEYINPUT6), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n235), .A2(G143), .ZN(new_n305));
  INV_X1    g119(.A(G143), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G146), .ZN(new_n307));
  AND2_X1   g121(.A1(KEYINPUT0), .A2(G128), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(G143), .B(G146), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT0), .B(G128), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n309), .B(G125), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT1), .ZN(new_n313));
  AND4_X1   g127(.A1(new_n313), .A2(new_n305), .A3(new_n307), .A4(G128), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT1), .B1(new_n306), .B2(G146), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n315), .A2(G128), .B1(new_n305), .B2(new_n307), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n312), .B1(new_n317), .B2(G125), .ZN(new_n318));
  INV_X1    g132(.A(G953), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G224), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n318), .B(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT6), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n299), .A2(new_n322), .A3(new_n301), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n304), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n320), .A2(KEYINPUT7), .ZN(new_n325));
  OR2_X1    g139(.A1(new_n318), .A2(new_n325), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n303), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n287), .A2(KEYINPUT81), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n286), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n287), .A2(KEYINPUT81), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n270), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n283), .ZN(new_n332));
  XOR2_X1   g146(.A(new_n300), .B(KEYINPUT8), .Z(new_n333));
  AOI22_X1  g147(.A1(new_n268), .A2(new_n269), .B1(new_n286), .B2(new_n287), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n333), .B1(new_n334), .B2(new_n282), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n315), .A2(G128), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n305), .A2(new_n307), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n310), .A2(G128), .A3(new_n315), .ZN(new_n339));
  AOI21_X1  g153(.A(G125), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n312), .ZN(new_n341));
  OAI211_X1 g155(.A(KEYINPUT7), .B(new_n320), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT82), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n318), .A2(KEYINPUT82), .A3(KEYINPUT7), .A4(new_n320), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n332), .A2(new_n335), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(G902), .B1(new_n327), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(G210), .B1(G237), .B2(G902), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n324), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n348), .B1(new_n324), .B2(new_n347), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n257), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n193), .A2(KEYINPUT9), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT9), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G234), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n352), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n355), .B1(new_n352), .B2(new_n354), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n192), .B1(new_n359), .B2(new_n188), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n317), .A2(new_n282), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n278), .B(new_n281), .C1(new_n314), .C2(new_n316), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT64), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT11), .ZN(new_n366));
  INV_X1    g180(.A(G137), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n365), .A2(new_n366), .A3(new_n367), .A4(G134), .ZN(new_n368));
  INV_X1    g182(.A(G134), .ZN(new_n369));
  OAI22_X1  g183(.A1(new_n369), .A2(G137), .B1(KEYINPUT64), .B2(KEYINPUT11), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n369), .A2(G137), .B1(KEYINPUT64), .B2(KEYINPUT11), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G131), .ZN(new_n374));
  INV_X1    g188(.A(G131), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n375), .A3(new_n372), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n364), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT12), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n364), .A2(KEYINPUT12), .A3(new_n377), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT10), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n363), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n386), .B(new_n295), .C1(new_n296), .C2(new_n297), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n338), .A2(new_n339), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n283), .A2(new_n388), .A3(KEYINPUT10), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n384), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n371), .A2(new_n375), .A3(new_n372), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n375), .B1(new_n371), .B2(new_n372), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT80), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT80), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n374), .A2(new_n394), .A3(new_n376), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n390), .A2(new_n397), .ZN(new_n398));
  XOR2_X1   g212(.A(G110), .B(G140), .Z(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(KEYINPUT79), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n319), .A2(G227), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n400), .B(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n382), .A2(new_n398), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n384), .A2(new_n387), .A3(new_n389), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n405), .A2(new_n377), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n396), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n402), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AOI211_X1 g222(.A(G469), .B(G902), .C1(new_n404), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n405), .A2(new_n377), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n398), .A2(new_n410), .A3(new_n403), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n380), .A2(new_n381), .B1(new_n390), .B2(new_n397), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n411), .B(G469), .C1(new_n412), .C2(new_n403), .ZN(new_n413));
  INV_X1    g227(.A(G469), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(new_n188), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n361), .B1(new_n409), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT85), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n419), .B1(new_n259), .B2(G122), .ZN(new_n420));
  INV_X1    g234(.A(G122), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(KEYINPUT85), .A3(G116), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n420), .A2(new_n422), .B1(new_n259), .B2(G122), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n199), .A2(G143), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n306), .A2(G128), .ZN(new_n425));
  OAI21_X1  g239(.A(G134), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n306), .A2(G128), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n199), .A2(G143), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n428), .A3(new_n369), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n274), .A2(new_n423), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n420), .A2(new_n422), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n259), .A2(G122), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT14), .ZN(new_n433));
  OR3_X1    g247(.A1(new_n421), .A2(KEYINPUT14), .A3(G116), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G107), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n430), .A2(new_n436), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n431), .A2(new_n274), .A3(new_n432), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n274), .B1(new_n431), .B2(new_n432), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n429), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT13), .B1(new_n306), .B2(G128), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n427), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n442), .A2(KEYINPUT86), .B1(KEYINPUT13), .B2(new_n424), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT86), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n444), .A3(new_n427), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n369), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n437), .B1(new_n440), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT87), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n187), .A2(G953), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n448), .B1(new_n359), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n352), .A2(new_n354), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT78), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n356), .A3(new_n449), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(KEYINPUT87), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT88), .B1(new_n447), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n429), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n431), .A2(new_n432), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G107), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n423), .A2(new_n274), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n442), .A2(KEYINPUT86), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n424), .A2(KEYINPUT13), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n445), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G134), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT88), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n359), .A2(new_n448), .A3(new_n449), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n453), .A2(KEYINPUT87), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n466), .A2(new_n467), .A3(new_n470), .A4(new_n437), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n447), .A2(new_n455), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n456), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G478), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(KEYINPUT15), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n473), .A2(new_n188), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n476), .B1(new_n473), .B2(new_n188), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(KEYINPUT18), .A2(G131), .ZN(new_n480));
  OR2_X1    g294(.A1(KEYINPUT69), .A2(G237), .ZN(new_n481));
  NAND2_X1  g295(.A1(KEYINPUT69), .A2(G237), .ZN(new_n482));
  AOI21_X1  g296(.A(G953), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(G143), .A3(G214), .ZN(new_n484));
  AND2_X1   g298(.A1(KEYINPUT69), .A2(G237), .ZN(new_n485));
  NOR2_X1   g299(.A1(KEYINPUT69), .A2(G237), .ZN(new_n486));
  OAI211_X1 g300(.A(G214), .B(new_n319), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n306), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n480), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n484), .A2(new_n488), .A3(new_n480), .ZN(new_n491));
  XNOR2_X1  g305(.A(G125), .B(G140), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(new_n235), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n490), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  XOR2_X1   g308(.A(G113), .B(G122), .Z(new_n495));
  XOR2_X1   g309(.A(KEYINPUT84), .B(G104), .Z(new_n496));
  XOR2_X1   g310(.A(new_n495), .B(new_n496), .Z(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n484), .A2(new_n488), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(G131), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT17), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n484), .A2(new_n488), .A3(new_n375), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n237), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n499), .A2(KEYINPUT17), .A3(G131), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n494), .B(new_n498), .C1(new_n503), .C2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT19), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n492), .B(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n231), .B1(new_n509), .B2(G146), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n510), .B1(new_n500), .B2(new_n502), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n491), .A2(new_n493), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n512), .A2(new_n489), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n497), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n507), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT20), .ZN(new_n516));
  NOR2_X1   g330(.A1(G475), .A2(G902), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n519));
  INV_X1    g333(.A(new_n517), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n520), .B1(new_n507), .B2(new_n514), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n518), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n507), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(new_n504), .A3(new_n505), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n498), .B1(new_n525), .B2(new_n494), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n188), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(G475), .ZN(new_n528));
  INV_X1    g342(.A(G952), .ZN(new_n529));
  AOI211_X1 g343(.A(G953), .B(new_n529), .C1(G234), .C2(G237), .ZN(new_n530));
  AOI211_X1 g344(.A(new_n188), .B(new_n319), .C1(G234), .C2(G237), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT21), .B(G898), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n479), .A2(new_n522), .A3(new_n528), .A4(new_n534), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n351), .A2(new_n418), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT74), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n369), .A2(G137), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n367), .A2(G134), .ZN(new_n539));
  OAI21_X1  g353(.A(G131), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n376), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT66), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT66), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n376), .A2(new_n543), .A3(new_n540), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n388), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n386), .B1(new_n391), .B2(new_n392), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT65), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(KEYINPUT65), .B(new_n386), .C1(new_n391), .C2(new_n392), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n545), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT30), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n290), .A2(new_n291), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n270), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n388), .A2(new_n376), .A3(new_n540), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n546), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(new_n551), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n552), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n483), .A2(G210), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT26), .B(G101), .ZN(new_n563));
  OR2_X1    g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n563), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n556), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n292), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n559), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT31), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n556), .A2(new_n554), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n557), .B1(new_n550), .B2(new_n551), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n572), .B1(new_n573), .B2(new_n554), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n574), .A2(KEYINPUT31), .A3(new_n566), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT72), .ZN(new_n576));
  XOR2_X1   g390(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT65), .B1(new_n377), .B2(new_n386), .ZN(new_n579));
  INV_X1    g393(.A(new_n549), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n292), .B1(new_n581), .B2(new_n545), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n576), .B(new_n578), .C1(new_n582), .C2(new_n572), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n572), .B1(new_n550), .B2(new_n554), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT72), .B1(new_n584), .B2(new_n577), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT28), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n568), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n583), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n566), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n571), .A2(new_n575), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(G472), .A2(G902), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT32), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT32), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n569), .A2(new_n570), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT31), .B1(new_n574), .B2(new_n566), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n587), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n584), .A2(new_n577), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n598), .B1(new_n599), .B2(new_n576), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n566), .B1(new_n600), .B2(new_n585), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n594), .B(new_n591), .C1(new_n597), .C2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n593), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(G472), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n559), .A2(new_n568), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT29), .B1(new_n605), .B2(new_n589), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n583), .A2(new_n585), .A3(new_n566), .A4(new_n587), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n292), .B1(new_n546), .B2(new_n555), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT28), .B1(new_n572), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT29), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n564), .B2(new_n565), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n587), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n613), .A2(KEYINPUT73), .A3(new_n188), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT73), .B1(new_n613), .B2(new_n188), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n604), .B1(new_n608), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n537), .B1(new_n603), .B2(new_n618), .ZN(new_n619));
  AOI211_X1 g433(.A(KEYINPUT74), .B(new_n617), .C1(new_n593), .C2(new_n602), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n256), .B(new_n536), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n471), .A2(new_n472), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n461), .A2(new_n465), .B1(new_n436), .B2(new_n430), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n467), .B1(new_n625), .B2(new_n470), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n623), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n437), .B(KEYINPUT89), .C1(new_n440), .C2(new_n446), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT90), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n470), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n629), .B1(new_n450), .B2(new_n454), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n631), .A2(KEYINPUT89), .B1(new_n466), .B2(new_n437), .ZN(new_n632));
  OAI21_X1  g446(.A(KEYINPUT33), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n474), .A2(G902), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n627), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT91), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n627), .A2(new_n633), .A3(KEYINPUT91), .A4(new_n634), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n473), .A2(new_n188), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n474), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n637), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n522), .A2(new_n528), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n257), .B(new_n534), .C1(new_n349), .C2(new_n350), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n645), .B(KEYINPUT92), .Z(new_n646));
  NOR3_X1   g460(.A1(new_n253), .A2(new_n418), .A3(new_n255), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n571), .A2(new_n575), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n588), .A2(new_n589), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n591), .ZN(new_n651));
  OAI21_X1  g465(.A(G472), .B1(new_n590), .B2(G902), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n647), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n646), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT34), .B(G104), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G6));
  INV_X1    g471(.A(new_n479), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n521), .B(new_n519), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n658), .A2(new_n528), .A3(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n644), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n654), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT35), .B(G107), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G9));
  NAND2_X1  g478(.A1(new_n251), .A2(new_n252), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n189), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n246), .A2(new_n247), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n196), .A2(KEYINPUT36), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n189), .A2(G902), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n536), .A2(new_n672), .A3(new_n651), .A4(new_n652), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT93), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT37), .B(G110), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  AOI21_X1  g490(.A(new_n594), .B1(new_n650), .B2(new_n591), .ZN(new_n677));
  AOI211_X1 g491(.A(KEYINPUT32), .B(new_n592), .C1(new_n648), .C2(new_n649), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n618), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT74), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n603), .A2(new_n537), .A3(new_n618), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(G900), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n531), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n530), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n659), .A2(new_n528), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n479), .ZN(new_n689));
  AOI22_X1  g503(.A1(new_n665), .A2(new_n189), .B1(new_n670), .B2(new_n669), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n690), .A2(new_n351), .A3(new_n418), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n682), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G128), .ZN(G30));
  NOR2_X1   g507(.A1(new_n349), .A2(new_n350), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT38), .ZN(new_n695));
  INV_X1    g509(.A(new_n257), .ZN(new_n696));
  INV_X1    g510(.A(new_n478), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n473), .A2(new_n188), .A3(new_n476), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n642), .A2(new_n699), .ZN(new_n700));
  OR3_X1    g514(.A1(new_n695), .A2(new_n672), .A3(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n604), .A2(new_n188), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n569), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n572), .A2(new_n609), .ZN(new_n705));
  OAI21_X1  g519(.A(G472), .B1(new_n705), .B2(new_n566), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n703), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(new_n707), .B(KEYINPUT94), .Z(new_n708));
  NAND2_X1  g522(.A1(new_n603), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT95), .ZN(new_n711));
  OR3_X1    g525(.A1(new_n701), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n711), .B1(new_n701), .B2(new_n710), .ZN(new_n713));
  INV_X1    g527(.A(new_n418), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n686), .B(KEYINPUT39), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(new_n716), .B(KEYINPUT40), .Z(new_n717));
  NAND3_X1  g531(.A1(new_n712), .A2(new_n713), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G143), .ZN(G45));
  NAND3_X1  g533(.A1(new_n641), .A2(new_n642), .A3(new_n686), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT96), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n641), .A2(KEYINPUT96), .A3(new_n642), .A4(new_n686), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n682), .A2(new_n691), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G146), .ZN(G48));
  INV_X1    g541(.A(KEYINPUT97), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n404), .A2(new_n408), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n728), .B1(new_n729), .B2(G902), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT98), .ZN(new_n731));
  AOI21_X1  g545(.A(G902), .B1(new_n404), .B2(new_n408), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(KEYINPUT97), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n730), .A2(new_n731), .A3(G469), .A4(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n731), .B1(new_n732), .B2(new_n414), .ZN(new_n735));
  OAI21_X1  g549(.A(G469), .B1(new_n732), .B2(KEYINPUT97), .ZN(new_n736));
  AOI211_X1 g550(.A(new_n728), .B(G902), .C1(new_n404), .C2(new_n408), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n360), .B1(new_n734), .B2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n682), .A2(new_n646), .A3(new_n256), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT41), .B(G113), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G15));
  NAND4_X1  g556(.A1(new_n682), .A2(new_n256), .A3(new_n661), .A4(new_n739), .ZN(new_n743));
  XNOR2_X1  g557(.A(KEYINPUT99), .B(G116), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(G18));
  INV_X1    g559(.A(new_n351), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n739), .A2(new_n746), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n747), .A2(new_n535), .A3(new_n690), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n682), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G119), .ZN(G21));
  NAND2_X1  g564(.A1(new_n734), .A2(new_n738), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n700), .A2(new_n694), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n751), .A2(new_n752), .A3(new_n361), .A4(new_n534), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT100), .B(G472), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n754), .B1(new_n590), .B2(G902), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n566), .B1(new_n610), .B2(new_n587), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n591), .B1(new_n597), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n755), .A2(new_n256), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n421), .ZN(G24));
  AND3_X1   g574(.A1(new_n722), .A2(KEYINPUT101), .A3(new_n723), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT101), .B1(new_n722), .B2(new_n723), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n747), .A2(new_n690), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n755), .A2(new_n757), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G125), .ZN(G27));
  INV_X1    g581(.A(KEYINPUT42), .ZN(new_n768));
  INV_X1    g582(.A(new_n694), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(new_n696), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n714), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n256), .B(new_n772), .C1(new_n619), .C2(new_n620), .ZN(new_n773));
  INV_X1    g587(.A(new_n763), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n768), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n603), .A2(KEYINPUT102), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT102), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n593), .A2(new_n777), .A3(new_n602), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n776), .A2(new_n618), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n771), .A2(new_n768), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n779), .A2(new_n763), .A3(new_n256), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n775), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G131), .ZN(G33));
  INV_X1    g597(.A(new_n689), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n773), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(new_n369), .ZN(G36));
  OR2_X1    g600(.A1(new_n521), .A2(new_n519), .ZN(new_n787));
  AOI22_X1  g601(.A1(new_n787), .A2(new_n518), .B1(G475), .B2(new_n527), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT43), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n641), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n789), .B1(new_n641), .B2(new_n788), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(G902), .B1(new_n648), .B2(new_n649), .ZN(new_n793));
  OAI22_X1  g607(.A1(new_n793), .A2(new_n604), .B1(new_n590), .B2(new_n592), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n792), .A2(new_n794), .A3(KEYINPUT44), .A4(new_n672), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT103), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n690), .B1(new_n652), .B2(new_n651), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT103), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n797), .A2(new_n798), .A3(KEYINPUT44), .A4(new_n792), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n796), .A2(new_n770), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT104), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT104), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n796), .A2(new_n802), .A3(new_n770), .A4(new_n799), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT44), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n794), .A2(new_n672), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n790), .A2(new_n791), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT105), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g623(.A(KEYINPUT105), .B(new_n804), .C1(new_n805), .C2(new_n806), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n801), .A2(new_n803), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT106), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n801), .A2(KEYINPUT106), .A3(new_n803), .A4(new_n811), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n411), .B1(new_n412), .B2(new_n403), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT45), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n414), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n411), .B(KEYINPUT45), .C1(new_n412), .C2(new_n403), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n415), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n820), .A2(KEYINPUT46), .ZN(new_n821));
  INV_X1    g635(.A(new_n409), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n822), .B1(new_n820), .B2(KEYINPUT46), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n361), .B(new_n715), .C1(new_n821), .C2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n814), .A2(new_n815), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G137), .ZN(G39));
  INV_X1    g641(.A(new_n256), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(new_n722), .A3(new_n723), .A4(new_n770), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n682), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n361), .B1(new_n821), .B2(new_n823), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n831), .B(KEYINPUT47), .Z(new_n832));
  NAND2_X1  g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(KEYINPUT107), .B(G140), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n833), .B(new_n834), .ZN(G42));
  NOR3_X1   g649(.A1(new_n828), .A2(new_n696), .A3(new_n360), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(new_n788), .A3(new_n641), .A4(new_n695), .ZN(new_n837));
  INV_X1    g651(.A(new_n751), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n837), .B1(KEYINPUT49), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(KEYINPUT49), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n840), .B(KEYINPUT108), .Z(new_n841));
  NAND3_X1  g655(.A1(new_n839), .A2(new_n841), .A3(new_n710), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n739), .A2(new_n770), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n843), .A2(new_n530), .A3(new_n792), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(new_n256), .A3(new_n779), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT48), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n529), .A2(G953), .ZN(new_n847));
  AND4_X1   g661(.A1(new_n256), .A2(new_n710), .A3(new_n530), .A4(new_n843), .ZN(new_n848));
  INV_X1    g662(.A(new_n643), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n806), .A2(new_n758), .A3(new_n685), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(new_n746), .A3(new_n739), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n846), .A2(new_n847), .A3(new_n850), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT112), .ZN(new_n855));
  INV_X1    g669(.A(new_n739), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n855), .B1(new_n856), .B2(new_n257), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n739), .A2(KEYINPUT112), .A3(new_n696), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n695), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT113), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n851), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n859), .A2(new_n860), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n854), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT50), .ZN(new_n865));
  NOR2_X1   g679(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n838), .A2(new_n361), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n770), .B(new_n851), .C1(new_n832), .C2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n641), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n848), .A2(new_n788), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n844), .A2(new_n672), .A3(new_n765), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n868), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n866), .B1(new_n872), .B2(KEYINPUT51), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n853), .B1(new_n865), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n865), .A2(KEYINPUT115), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n872), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n874), .B1(new_n876), .B2(KEYINPUT51), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n654), .A2(new_n645), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT109), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n621), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n881), .B1(new_n621), .B2(new_n880), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n785), .B1(new_n775), .B2(new_n781), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n658), .A2(new_n522), .A3(new_n528), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n644), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n647), .A2(new_n887), .A3(new_n652), .A4(new_n651), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n673), .B(new_n888), .C1(new_n758), .C2(new_n753), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n682), .B2(new_n748), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n740), .A2(new_n890), .A3(new_n743), .ZN(new_n891));
  AOI211_X1 g705(.A(new_n658), .B(new_n688), .C1(new_n680), .C2(new_n681), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n763), .A2(new_n765), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n672), .B(new_n772), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n884), .A2(new_n885), .A3(new_n891), .A4(new_n894), .ZN(new_n895));
  OAI221_X1 g709(.A(new_n691), .B1(new_n725), .B2(new_n689), .C1(new_n619), .C2(new_n620), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n418), .B1(new_n685), .B2(new_n684), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT110), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n897), .A2(new_n898), .A3(new_n690), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n898), .B1(new_n897), .B2(new_n690), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n709), .B(new_n752), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n896), .A2(new_n766), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT52), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n896), .A2(KEYINPUT52), .A3(new_n766), .A4(new_n901), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n879), .B1(new_n895), .B2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n785), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n894), .A2(new_n782), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n740), .A2(new_n890), .A3(new_n743), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n910), .A2(new_n882), .A3(new_n883), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n904), .A2(new_n905), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n909), .A2(new_n911), .A3(KEYINPUT53), .A4(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n878), .B1(new_n907), .B2(new_n913), .ZN(new_n914));
  XOR2_X1   g728(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n915));
  NAND3_X1  g729(.A1(new_n907), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n877), .A2(new_n914), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(G952), .A2(G953), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT116), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n842), .B1(new_n918), .B2(new_n920), .ZN(G75));
  NOR2_X1   g735(.A1(new_n319), .A2(G952), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n188), .B1(new_n907), .B2(new_n913), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT56), .B1(new_n924), .B2(G210), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n304), .A2(new_n323), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(new_n321), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT55), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n923), .B1(new_n925), .B2(new_n929), .ZN(new_n930));
  AOI211_X1 g744(.A(KEYINPUT56), .B(new_n928), .C1(new_n924), .C2(G210), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT117), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n907), .A2(new_n913), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n933), .A2(G210), .A3(G902), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n928), .B1(new_n934), .B2(KEYINPUT56), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT117), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n925), .A2(new_n929), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n935), .A2(new_n936), .A3(new_n937), .A4(new_n923), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n932), .A2(new_n938), .ZN(G51));
  XNOR2_X1  g753(.A(new_n415), .B(KEYINPUT57), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n915), .B1(new_n907), .B2(new_n913), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n940), .B1(new_n917), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n729), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n924), .A2(new_n819), .A3(new_n818), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n922), .B1(new_n944), .B2(new_n945), .ZN(G54));
  AND2_X1   g760(.A1(KEYINPUT58), .A2(G475), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n924), .A2(new_n515), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n515), .B1(new_n924), .B2(new_n947), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n948), .A2(new_n949), .A3(new_n922), .ZN(G60));
  INV_X1    g764(.A(KEYINPUT118), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n627), .A2(new_n633), .ZN(new_n952));
  NAND2_X1  g766(.A1(G478), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT59), .Z(new_n954));
  NOR2_X1   g768(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n915), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n933), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n956), .B1(new_n958), .B2(new_n916), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n951), .B1(new_n959), .B2(new_n922), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n955), .B1(new_n917), .B2(new_n941), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n961), .A2(KEYINPUT118), .A3(new_n923), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n917), .A2(new_n914), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n952), .B1(new_n963), .B2(new_n954), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n960), .A2(new_n962), .A3(new_n964), .ZN(G63));
  XNOR2_X1  g779(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n187), .A2(new_n188), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n907), .B2(new_n913), .ZN(new_n970));
  INV_X1    g784(.A(new_n254), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n923), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT61), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n970), .A2(new_n669), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n973), .A2(KEYINPUT120), .A3(new_n974), .A4(new_n975), .ZN(new_n976));
  OR2_X1    g790(.A1(new_n974), .A2(KEYINPUT120), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n974), .A2(KEYINPUT120), .ZN(new_n978));
  INV_X1    g792(.A(new_n975), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n977), .B(new_n978), .C1(new_n979), .C2(new_n972), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n976), .A2(new_n980), .ZN(G66));
  INV_X1    g795(.A(new_n532), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n319), .B1(new_n982), .B2(G224), .ZN(new_n983));
  INV_X1    g797(.A(new_n911), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n983), .B1(new_n984), .B2(new_n319), .ZN(new_n985));
  INV_X1    g799(.A(G898), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n926), .B1(new_n986), .B2(G953), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n985), .B(new_n987), .ZN(G69));
  INV_X1    g802(.A(KEYINPUT125), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n573), .B(new_n509), .Z(new_n990));
  INV_X1    g804(.A(new_n752), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n824), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n779), .A2(new_n992), .A3(new_n256), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(KEYINPUT122), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT122), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n779), .A2(new_n992), .A3(new_n995), .A4(new_n256), .ZN(new_n996));
  AOI22_X1  g810(.A1(new_n994), .A2(new_n996), .B1(new_n830), .B2(new_n832), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n885), .A2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT121), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n896), .A2(new_n999), .A3(new_n766), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n999), .B1(new_n896), .B2(new_n766), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(G953), .B1(new_n1003), .B2(new_n826), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n319), .A2(G900), .ZN(new_n1005));
  NOR3_X1   g819(.A1(new_n1004), .A2(KEYINPUT123), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT123), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n815), .A2(new_n825), .ZN(new_n1008));
  AOI22_X1  g822(.A1(new_n800), .A2(KEYINPUT104), .B1(new_n809), .B2(new_n810), .ZN(new_n1009));
  AOI21_X1  g823(.A(KEYINPUT106), .B1(new_n1009), .B2(new_n803), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n885), .B(new_n997), .C1(new_n1001), .C2(new_n1000), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n319), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1005), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1007), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n989), .B(new_n990), .C1(new_n1006), .C2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n319), .B1(G227), .B2(G900), .ZN(new_n1017));
  INV_X1    g831(.A(new_n990), .ZN(new_n1018));
  OAI21_X1  g832(.A(KEYINPUT123), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1013), .A2(new_n1007), .A3(new_n1014), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(new_n886), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n715), .B1(new_n849), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n833), .B1(new_n773), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1008), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1024), .B1(new_n1025), .B2(new_n814), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n718), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1027));
  INV_X1    g841(.A(KEYINPUT62), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI211_X1 g843(.A(KEYINPUT62), .B(new_n718), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(G953), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g846(.A(KEYINPUT125), .B1(new_n1032), .B2(new_n990), .ZN(new_n1033));
  OAI211_X1 g847(.A(new_n1016), .B(new_n1017), .C1(new_n1021), .C2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n990), .B1(new_n1006), .B2(new_n1015), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1017), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1036), .B1(new_n1032), .B2(new_n990), .ZN(new_n1037));
  INV_X1    g851(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g852(.A(KEYINPUT124), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g853(.A(KEYINPUT124), .ZN(new_n1040));
  NOR3_X1   g854(.A1(new_n1021), .A2(new_n1040), .A3(new_n1037), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n1034), .B1(new_n1039), .B2(new_n1041), .ZN(G72));
  XNOR2_X1  g856(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1043));
  XNOR2_X1  g857(.A(new_n703), .B(new_n1043), .ZN(new_n1044));
  INV_X1    g858(.A(new_n1044), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n574), .A2(new_n566), .ZN(new_n1046));
  OAI211_X1 g860(.A(new_n933), .B(new_n1045), .C1(new_n1046), .C2(new_n704), .ZN(new_n1047));
  NOR3_X1   g861(.A1(new_n1011), .A2(new_n984), .A3(new_n1012), .ZN(new_n1048));
  OAI211_X1 g862(.A(new_n589), .B(new_n574), .C1(new_n1048), .C2(new_n1044), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n1047), .A2(new_n923), .A3(new_n1049), .ZN(new_n1050));
  NAND3_X1  g864(.A1(new_n1026), .A2(new_n1031), .A3(new_n911), .ZN(new_n1051));
  AOI211_X1 g865(.A(new_n589), .B(new_n574), .C1(new_n1051), .C2(new_n1045), .ZN(new_n1052));
  NOR2_X1   g866(.A1(new_n1050), .A2(new_n1052), .ZN(G57));
endmodule


