//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985;
  INV_X1    g000(.A(KEYINPUT65), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G146), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT64), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n189), .B1(new_n194), .B2(new_n188), .ZN(new_n195));
  AND2_X1   g009(.A1(KEYINPUT0), .A2(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n187), .B1(new_n195), .B2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n191), .A2(new_n193), .A3(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n188), .A2(G146), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(new_n196), .ZN(new_n204));
  INV_X1    g018(.A(new_n189), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT64), .B(G146), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(G143), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT65), .A3(new_n198), .ZN(new_n208));
  AND3_X1   g022(.A1(new_n200), .A2(new_n204), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G137), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT11), .A3(G134), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT67), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(G134), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT11), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI211_X1 g031(.A(KEYINPUT66), .B(KEYINPUT11), .C1(new_n210), .C2(G134), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n213), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G134), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G137), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n212), .B1(new_n211), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(G131), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n216), .B1(new_n220), .B2(G137), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n215), .A2(new_n214), .A3(new_n216), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n211), .A2(new_n221), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT67), .ZN(new_n229));
  INV_X1    g043(.A(G131), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n227), .A2(new_n229), .A3(new_n230), .A4(new_n213), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n223), .A2(KEYINPUT71), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT71), .B1(new_n223), .B2(new_n231), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n209), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G119), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT68), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G119), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n238), .A3(G116), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT69), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT68), .B(G119), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n242), .A3(G116), .ZN(new_n243));
  INV_X1    g057(.A(G116), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G119), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n240), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  XOR2_X1   g060(.A(KEYINPUT2), .B(G113), .Z(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n239), .A2(KEYINPUT69), .B1(new_n244), .B2(G119), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(new_n247), .A3(new_n243), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n249), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n250), .B1(new_n249), .B2(new_n252), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G128), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(KEYINPUT1), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n201), .A2(new_n202), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n256), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(new_n195), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n215), .A2(new_n221), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G131), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n260), .A2(new_n231), .A3(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n234), .A2(new_n255), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(KEYINPUT28), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n263), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n223), .A2(new_n231), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n223), .A2(KEYINPUT71), .A3(new_n231), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n268), .B1(new_n273), .B2(new_n209), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(new_n255), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT28), .B1(new_n275), .B2(new_n265), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n267), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G237), .ZN(new_n278));
  INV_X1    g092(.A(G953), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(new_n279), .A3(G210), .ZN(new_n280));
  XOR2_X1   g094(.A(new_n280), .B(KEYINPUT27), .Z(new_n281));
  XNOR2_X1  g095(.A(new_n281), .B(KEYINPUT26), .ZN(new_n282));
  INV_X1    g096(.A(G101), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n282), .B(new_n283), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n284), .A2(KEYINPUT29), .ZN(new_n285));
  AOI21_X1  g099(.A(G902), .B1(new_n277), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n274), .A2(KEYINPUT30), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n249), .A2(new_n252), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT70), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n249), .A2(new_n250), .A3(new_n252), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n231), .A2(new_n262), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n209), .A2(new_n269), .B1(new_n292), .B2(new_n260), .ZN(new_n293));
  OR2_X1    g107(.A1(new_n293), .A2(KEYINPUT30), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n287), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n264), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n296), .A2(new_n284), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT72), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n298), .B1(new_n255), .B2(new_n293), .ZN(new_n299));
  INV_X1    g113(.A(new_n269), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n200), .A2(new_n204), .A3(new_n208), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n263), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(new_n291), .A3(KEYINPUT72), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n299), .A2(new_n264), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT28), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT73), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n304), .A2(new_n307), .A3(KEYINPUT28), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n306), .A2(new_n267), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n297), .B1(new_n309), .B2(new_n284), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n286), .B1(new_n310), .B2(KEYINPUT29), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G472), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n295), .A2(new_n264), .A3(new_n284), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(KEYINPUT31), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n304), .A2(new_n307), .A3(KEYINPUT28), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n307), .B1(new_n304), .B2(KEYINPUT28), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n315), .A2(new_n316), .A3(new_n266), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT74), .B1(new_n317), .B2(new_n284), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n319));
  INV_X1    g133(.A(new_n284), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n309), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n314), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(G472), .A2(G902), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT32), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n312), .B1(new_n322), .B2(new_n327), .ZN(new_n328));
  XOR2_X1   g142(.A(new_n313), .B(KEYINPUT31), .Z(new_n329));
  AOI21_X1  g143(.A(new_n266), .B1(new_n305), .B2(KEYINPUT73), .ZN(new_n330));
  AOI211_X1 g144(.A(KEYINPUT74), .B(new_n284), .C1(new_n330), .C2(new_n308), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n319), .B1(new_n309), .B2(new_n320), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n329), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT32), .B1(new_n333), .B2(new_n323), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT75), .B1(new_n328), .B2(new_n334), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n333), .A2(new_n326), .B1(new_n311), .B2(G472), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n325), .B1(new_n322), .B2(new_n324), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT23), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n341), .B1(new_n241), .B2(G128), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n235), .A2(new_n256), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n343), .B1(new_n241), .B2(new_n256), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n342), .B1(new_n344), .B2(new_n341), .ZN(new_n345));
  XOR2_X1   g159(.A(KEYINPUT24), .B(G110), .Z(new_n346));
  OAI22_X1  g160(.A1(new_n345), .A2(G110), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT77), .B(G125), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n348), .A2(KEYINPUT16), .A3(G140), .ZN(new_n349));
  NOR2_X1   g163(.A1(G125), .A2(G140), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G140), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n351), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n349), .B1(KEYINPUT16), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G146), .ZN(new_n355));
  XNOR2_X1  g169(.A(G125), .B(G140), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n206), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(KEYINPUT78), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n347), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  OR2_X1    g173(.A1(new_n354), .A2(G146), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n355), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n344), .A2(new_n346), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n345), .A2(G110), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(KEYINPUT76), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n359), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n279), .A2(G221), .A3(G234), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(KEYINPUT22), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(G137), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OR2_X1    g184(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G902), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n366), .A2(new_n370), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  OR2_X1    g188(.A1(new_n374), .A2(KEYINPUT25), .ZN(new_n375));
  INV_X1    g189(.A(G234), .ZN(new_n376));
  OAI21_X1  g190(.A(G217), .B1(new_n376), .B2(G902), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n377), .B1(new_n374), .B2(KEYINPUT25), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n371), .A2(new_n373), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n377), .A2(new_n372), .ZN(new_n381));
  XOR2_X1   g195(.A(new_n381), .B(KEYINPUT79), .Z(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(G210), .B1(G237), .B2(G902), .ZN(new_n386));
  XOR2_X1   g200(.A(new_n386), .B(KEYINPUT92), .Z(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n348), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n301), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT91), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n391), .B1(new_n260), .B2(new_n389), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n390), .A2(KEYINPUT91), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n279), .A2(G224), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n394), .B(new_n395), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n251), .A2(KEYINPUT5), .A3(new_n243), .ZN(new_n397));
  OAI21_X1  g211(.A(G113), .B1(new_n239), .B2(KEYINPUT5), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n252), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G107), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G104), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT3), .ZN(new_n402));
  INV_X1    g216(.A(G104), .ZN(new_n403));
  AOI21_X1  g217(.A(G101), .B1(new_n403), .B2(G107), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT82), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n400), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT81), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT3), .ZN(new_n408));
  NAND2_X1  g222(.A1(KEYINPUT82), .A2(G107), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n406), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT3), .B1(new_n407), .B2(G104), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n402), .B(new_n404), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT83), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT3), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n414), .B1(new_n403), .B2(KEYINPUT81), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n415), .A2(new_n408), .A3(new_n406), .A4(new_n409), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT83), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n416), .A2(new_n417), .A3(new_n402), .A4(new_n404), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n406), .A2(new_n409), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n403), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n283), .B1(new_n421), .B2(new_n401), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n399), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n403), .A2(G107), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n402), .B(new_n426), .C1(new_n410), .C2(new_n411), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT4), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n427), .A2(new_n428), .A3(G101), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n428), .B1(new_n427), .B2(G101), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n429), .B1(new_n419), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n253), .B2(new_n254), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n425), .B1(new_n432), .B2(KEYINPUT88), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT88), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n291), .A2(new_n434), .A3(new_n431), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT89), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT6), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT89), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n433), .A2(new_n439), .A3(new_n435), .ZN(new_n440));
  XNOR2_X1  g254(.A(G110), .B(G122), .ZN(new_n441));
  XOR2_X1   g255(.A(new_n441), .B(KEYINPUT90), .Z(new_n442));
  NAND4_X1  g256(.A1(new_n437), .A2(new_n438), .A3(new_n440), .A4(new_n442), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n433), .A2(new_n439), .A3(new_n435), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n439), .B1(new_n433), .B2(new_n435), .ZN(new_n445));
  INV_X1    g259(.A(new_n442), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n433), .A2(new_n435), .A3(new_n446), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT6), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n396), .B(new_n443), .C1(new_n447), .C2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n394), .A2(KEYINPUT7), .A3(new_n395), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n395), .A2(KEYINPUT7), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(new_n392), .B2(new_n393), .ZN(new_n453));
  XOR2_X1   g267(.A(new_n442), .B(KEYINPUT8), .Z(new_n454));
  AND2_X1   g268(.A1(new_n399), .A2(new_n424), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n454), .B1(new_n455), .B2(new_n425), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n451), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(G902), .B1(new_n457), .B2(new_n448), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n388), .B1(new_n450), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT93), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n450), .A2(new_n458), .A3(new_n386), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n463), .B1(new_n459), .B2(new_n460), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT9), .B(G234), .ZN(new_n466));
  OAI21_X1  g280(.A(G221), .B1(new_n466), .B2(G902), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n279), .A2(G227), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(G140), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT80), .B(G110), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n469), .B(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n422), .B1(new_n413), .B2(new_n418), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n260), .A2(KEYINPUT10), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n431), .A2(new_n209), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n273), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT84), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n256), .B1(new_n205), .B2(KEYINPUT1), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n258), .B1(new_n203), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n419), .A2(new_n423), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT10), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n477), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI211_X1 g296(.A(KEYINPUT84), .B(KEYINPUT10), .C1(new_n473), .C2(new_n479), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n475), .B(new_n476), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n480), .B1(new_n260), .B2(new_n473), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT12), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n300), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT12), .B1(new_n485), .B2(new_n273), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n488), .B1(new_n489), .B2(KEYINPUT85), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT85), .ZN(new_n491));
  AOI211_X1 g305(.A(new_n491), .B(KEYINPUT12), .C1(new_n485), .C2(new_n273), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n472), .B(new_n484), .C1(new_n490), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT87), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n475), .B1(new_n483), .B2(new_n482), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n273), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(KEYINPUT86), .A3(new_n484), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT86), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n495), .A2(new_n498), .A3(new_n273), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n497), .A2(new_n471), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n497), .A2(KEYINPUT87), .A3(new_n471), .A4(new_n499), .ZN(new_n502));
  AOI211_X1 g316(.A(G469), .B(G902), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G469), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n497), .A2(new_n499), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n472), .ZN(new_n506));
  INV_X1    g320(.A(new_n484), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n485), .A2(new_n487), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n419), .A2(new_n423), .A3(new_n479), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n260), .B1(new_n419), .B2(new_n423), .ZN(new_n510));
  OAI22_X1  g324(.A1(new_n509), .A2(new_n510), .B1(new_n232), .B2(new_n233), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n486), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n508), .B1(new_n512), .B2(new_n491), .ZN(new_n513));
  INV_X1    g327(.A(new_n492), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n507), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n506), .B1(new_n472), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n504), .B1(new_n516), .B2(new_n372), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n467), .B1(new_n503), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(G214), .B1(G237), .B2(G902), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(G475), .A2(G902), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n278), .A2(new_n279), .A3(G214), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(G143), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G131), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n230), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT17), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n524), .A2(KEYINPUT17), .A3(G131), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n360), .A2(new_n528), .A3(new_n355), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(KEYINPUT18), .A2(G131), .ZN(new_n531));
  XOR2_X1   g345(.A(new_n523), .B(new_n531), .Z(new_n532));
  OAI21_X1  g346(.A(new_n358), .B1(new_n190), .B2(new_n353), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(G113), .B(G122), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(new_n403), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n525), .A2(new_n526), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT19), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n356), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n541), .B1(new_n353), .B2(new_n540), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n539), .B(new_n355), .C1(new_n194), .C2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n537), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n534), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n538), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n546), .A2(KEYINPUT94), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT94), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(new_n538), .B2(new_n545), .ZN(new_n549));
  OAI211_X1 g363(.A(KEYINPUT20), .B(new_n521), .C1(new_n547), .C2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT20), .ZN(new_n551));
  INV_X1    g365(.A(new_n521), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n551), .B1(new_n546), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n279), .A2(G952), .ZN(new_n555));
  NAND2_X1  g369(.A1(G234), .A2(G237), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(G902), .A3(G953), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT21), .B(G898), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n558), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n535), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n544), .A2(KEYINPUT95), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n372), .B1(new_n564), .B2(new_n565), .ZN(new_n567));
  OAI21_X1  g381(.A(G475), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT97), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n188), .B2(G128), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n256), .A2(KEYINPUT97), .A3(G143), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n572), .B1(new_n256), .B2(G143), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(G134), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n244), .A2(G122), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n244), .A2(G122), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n420), .ZN(new_n578));
  OR2_X1    g392(.A1(new_n577), .A2(new_n420), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n574), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  XOR2_X1   g394(.A(KEYINPUT96), .B(KEYINPUT13), .Z(new_n581));
  NOR2_X1   g395(.A1(new_n256), .A2(G143), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n572), .B1(new_n581), .B2(new_n582), .ZN(new_n584));
  OAI21_X1  g398(.A(G134), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n580), .A2(KEYINPUT98), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT98), .B1(new_n580), .B2(new_n585), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n573), .B(new_n220), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT99), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n579), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT100), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n591), .B1(new_n576), .B2(KEYINPUT14), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT14), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n593), .A2(new_n244), .A3(KEYINPUT100), .A4(G122), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n576), .A2(KEYINPUT14), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n592), .A2(new_n575), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(KEYINPUT101), .A3(G107), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(G107), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT101), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n597), .B(new_n600), .C1(new_n588), .C2(KEYINPUT99), .ZN(new_n601));
  OAI22_X1  g415(.A1(new_n586), .A2(new_n587), .B1(new_n590), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(G217), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n466), .A2(new_n603), .A3(G953), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  OAI221_X1 g420(.A(new_n604), .B1(new_n590), .B2(new_n601), .C1(new_n586), .C2(new_n587), .ZN(new_n607));
  AOI21_X1  g421(.A(G902), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(G478), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(KEYINPUT15), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n608), .B(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n554), .A2(new_n563), .A3(new_n568), .A4(new_n611), .ZN(new_n612));
  NOR4_X1   g426(.A1(new_n465), .A2(new_n518), .A3(new_n520), .A4(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n340), .A2(new_n385), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G101), .ZN(G3));
  OAI21_X1  g429(.A(G472), .B1(new_n322), .B2(G902), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n333), .A2(new_n323), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n617), .A3(new_n385), .ZN(new_n618));
  OR2_X1    g432(.A1(new_n618), .A2(new_n518), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n606), .A2(new_n607), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT33), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n606), .A2(new_n607), .A3(KEYINPUT33), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n609), .A2(G902), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT103), .ZN(new_n626));
  INV_X1    g440(.A(new_n608), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n626), .B1(new_n627), .B2(new_n609), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n608), .A2(KEYINPUT103), .A3(G478), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n550), .A2(new_n553), .A3(new_n568), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n386), .B1(new_n450), .B2(new_n458), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT102), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n463), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AOI211_X1 g449(.A(KEYINPUT102), .B(new_n386), .C1(new_n450), .C2(new_n458), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n519), .B(new_n632), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n619), .A2(new_n562), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT34), .B(G104), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  XNOR2_X1  g454(.A(new_n546), .B(KEYINPUT94), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n521), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n551), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n643), .A2(new_n550), .ZN(new_n644));
  INV_X1    g458(.A(new_n611), .ZN(new_n645));
  AND4_X1   g459(.A1(new_n563), .A2(new_n644), .A3(new_n568), .A4(new_n645), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n646), .B(new_n519), .C1(new_n636), .C2(new_n635), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n619), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT35), .B(G107), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  NOR2_X1   g464(.A1(new_n370), .A2(KEYINPUT36), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n366), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n366), .A2(new_n652), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n653), .A2(new_n382), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n375), .B2(new_n378), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n612), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n616), .A2(new_n617), .A3(new_n657), .ZN(new_n658));
  NOR4_X1   g472(.A1(new_n658), .A2(new_n465), .A3(new_n518), .A4(new_n520), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT37), .B(G110), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT104), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT105), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n659), .B(new_n662), .ZN(G12));
  NAND2_X1  g477(.A1(new_n643), .A2(new_n550), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT106), .B(G900), .Z(new_n665));
  AOI21_X1  g479(.A(new_n558), .B1(new_n560), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n568), .A2(new_n667), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n664), .A2(new_n611), .A3(new_n668), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n669), .B(new_n519), .C1(new_n635), .C2(new_n636), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n518), .A2(new_n656), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n337), .B1(new_n336), .B2(new_n338), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n671), .B(new_n672), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G128), .ZN(G30));
  XOR2_X1   g490(.A(new_n666), .B(KEYINPUT39), .Z(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n518), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n679), .B(KEYINPUT40), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n465), .B(KEYINPUT38), .ZN(new_n681));
  INV_X1    g495(.A(new_n631), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n611), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(G472), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n320), .B1(new_n275), .B2(new_n265), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n688), .A2(new_n313), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n685), .B1(new_n690), .B2(new_n372), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(new_n333), .B2(new_n326), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n684), .B1(new_n338), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n519), .A3(new_n656), .ZN(new_n694));
  OR3_X1    g508(.A1(new_n680), .A2(new_n681), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G143), .ZN(G45));
  NOR2_X1   g510(.A1(new_n637), .A2(new_n666), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n697), .B(new_n672), .C1(new_n673), .C2(new_n674), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  NOR2_X1   g513(.A1(new_n637), .A2(new_n562), .ZN(new_n700));
  AOI21_X1  g514(.A(G902), .B1(new_n501), .B2(new_n502), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n702));
  OAI21_X1  g516(.A(G469), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AOI211_X1 g517(.A(KEYINPUT108), .B(G902), .C1(new_n501), .C2(new_n502), .ZN(new_n704));
  OAI21_X1  g518(.A(KEYINPUT109), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n501), .A2(new_n502), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n372), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT108), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n701), .A2(new_n702), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n708), .A2(new_n709), .A3(G469), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n701), .A2(new_n504), .ZN(new_n712));
  AND4_X1   g526(.A1(new_n467), .A2(new_n705), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n340), .A2(new_n385), .A3(new_n700), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  INV_X1    g530(.A(new_n647), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n340), .A2(new_n717), .A3(new_n385), .A4(new_n713), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G116), .ZN(G18));
  AND3_X1   g533(.A1(new_n450), .A2(new_n458), .A3(new_n386), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n450), .A2(new_n458), .ZN(new_n721));
  INV_X1    g535(.A(new_n386), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n720), .B1(new_n723), .B2(KEYINPUT102), .ZN(new_n724));
  INV_X1    g538(.A(new_n636), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n520), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n340), .A2(new_n726), .A3(new_n657), .A4(new_n713), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  AOI21_X1  g542(.A(new_n284), .B1(new_n277), .B2(KEYINPUT110), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n729), .B1(KEYINPUT110), .B2(new_n277), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n324), .B1(new_n730), .B2(new_n329), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n616), .A2(new_n732), .ZN(new_n733));
  OAI211_X1 g547(.A(KEYINPUT111), .B(G472), .C1(new_n322), .C2(G902), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n731), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n519), .B1(new_n635), .B2(new_n636), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n736), .A2(new_n562), .A3(new_n684), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n713), .A2(new_n735), .A3(new_n737), .A4(new_n385), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT112), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G122), .ZN(G24));
  INV_X1    g554(.A(new_n656), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n713), .A2(new_n735), .A3(new_n741), .A4(new_n697), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G125), .ZN(G27));
  OAI211_X1 g557(.A(KEYINPUT42), .B(new_n385), .C1(new_n328), .C2(new_n334), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT113), .B1(new_n515), .B2(new_n472), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n484), .B1(new_n490), .B2(new_n492), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n747), .A3(new_n471), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n745), .A2(new_n506), .A3(G469), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(G469), .A2(G902), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n467), .B1(new_n503), .B2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n632), .A2(new_n667), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n465), .A2(new_n753), .A3(new_n755), .A4(new_n519), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n744), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n721), .A2(new_n387), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT93), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n759), .A2(new_n519), .A3(new_n461), .A4(new_n463), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n760), .A2(new_n754), .A3(new_n752), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n761), .B(new_n385), .C1(new_n673), .C2(new_n674), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n757), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT114), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G131), .ZN(G33));
  AOI21_X1  g580(.A(new_n384), .B1(new_n335), .B2(new_n339), .ZN(new_n767));
  INV_X1    g581(.A(new_n760), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n768), .A2(new_n669), .A3(new_n753), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(KEYINPUT115), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n220), .ZN(G36));
  INV_X1    g586(.A(new_n630), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n631), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(KEYINPUT116), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(KEYINPUT43), .Z(new_n776));
  NAND2_X1  g590(.A1(new_n616), .A2(new_n617), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n777), .A3(new_n741), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT44), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n467), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n516), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n745), .A2(new_n506), .A3(KEYINPUT45), .A4(new_n748), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(G469), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n750), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT46), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n503), .B1(new_n786), .B2(new_n787), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n781), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n791), .A2(new_n677), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n778), .A2(new_n779), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n780), .A2(new_n768), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G137), .ZN(G39));
  INV_X1    g609(.A(KEYINPUT47), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n791), .B(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n340), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(new_n384), .A3(new_n755), .A4(new_n768), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(new_n352), .ZN(G42));
  NAND4_X1  g615(.A1(new_n776), .A2(new_n385), .A3(new_n558), .A4(new_n735), .ZN(new_n802));
  OR2_X1    g616(.A1(KEYINPUT121), .A2(KEYINPUT50), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n681), .A2(new_n520), .A3(new_n713), .A4(new_n803), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(KEYINPUT121), .A2(KEYINPUT50), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  AOI211_X1 g622(.A(new_n656), .B(new_n731), .C1(new_n733), .C2(new_n734), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n705), .A2(new_n711), .A3(new_n712), .ZN(new_n810));
  NOR4_X1   g624(.A1(new_n810), .A2(new_n781), .A3(new_n557), .A4(new_n760), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n776), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n808), .B1(new_n809), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n338), .A2(new_n692), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n384), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n811), .A2(new_n682), .A3(new_n773), .A4(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n797), .B1(new_n467), .B2(new_n810), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n802), .A2(new_n760), .ZN(new_n819));
  AOI22_X1  g633(.A1(new_n818), .A2(new_n819), .B1(new_n807), .B2(new_n805), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n814), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n811), .A2(new_n632), .A3(new_n816), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n713), .A2(new_n726), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n825), .B(new_n555), .C1(new_n802), .C2(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n384), .B1(new_n336), .B2(new_n338), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n813), .A2(new_n828), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n829), .A2(KEYINPUT48), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(KEYINPUT48), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n827), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n823), .A2(new_n824), .A3(new_n832), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n518), .A2(new_n656), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n335), .B2(new_n339), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n655), .B(new_n666), .C1(new_n375), .C2(new_n378), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n467), .B(new_n836), .C1(new_n503), .C2(new_n751), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT120), .ZN(new_n838));
  AND4_X1   g652(.A1(new_n726), .A2(new_n815), .A3(new_n838), .A4(new_n683), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n837), .A2(KEYINPUT120), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n835), .A2(new_n697), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(KEYINPUT52), .A3(new_n675), .A4(new_n742), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n840), .A2(new_n693), .A3(new_n726), .A4(new_n838), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n742), .A2(new_n698), .A3(new_n675), .A4(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT52), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n631), .A2(new_n611), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n849));
  AOI22_X1  g663(.A1(new_n848), .A2(new_n849), .B1(new_n630), .B2(new_n631), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n849), .B2(new_n848), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n563), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n658), .B1(new_n852), .B2(new_n618), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n465), .A2(new_n518), .A3(new_n520), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n714), .A2(new_n614), .A3(new_n738), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n718), .A2(new_n727), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n856), .A2(new_n857), .A3(new_n764), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n847), .A2(new_n858), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n767), .A2(new_n769), .B1(new_n809), .B2(new_n761), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n644), .A2(new_n568), .A3(new_n611), .A4(new_n667), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n760), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n672), .B(new_n862), .C1(new_n673), .C2(new_n674), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT118), .B1(new_n835), .B2(new_n862), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n860), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n863), .A2(new_n864), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n835), .A2(KEYINPUT118), .A3(new_n862), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n872), .A2(KEYINPUT119), .A3(new_n860), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT53), .B1(new_n859), .B2(new_n874), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n872), .A2(KEYINPUT119), .A3(new_n860), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT119), .B1(new_n872), .B2(new_n860), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n847), .B(new_n858), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT54), .B1(new_n875), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n878), .A2(new_n879), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n874), .A2(KEYINPUT53), .A3(new_n847), .A4(new_n858), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n833), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(G952), .A2(G953), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT122), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n810), .A2(KEYINPUT49), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n810), .A2(KEYINPUT49), .ZN(new_n891));
  NOR4_X1   g705(.A1(new_n773), .A2(new_n781), .A3(new_n520), .A4(new_n631), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n681), .A2(new_n891), .A3(new_n816), .A4(new_n892), .ZN(new_n893));
  OAI22_X1  g707(.A1(new_n887), .A2(new_n889), .B1(new_n890), .B2(new_n893), .ZN(G75));
  NOR2_X1   g708(.A1(new_n279), .A2(G952), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n443), .B1(new_n447), .B2(new_n449), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(new_n396), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT55), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n372), .B1(new_n882), .B2(new_n884), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(G210), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT56), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n899), .A2(new_n387), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n898), .A2(new_n901), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n895), .B(new_n902), .C1(new_n903), .C2(new_n904), .ZN(G51));
  AOI211_X1 g719(.A(new_n372), .B(new_n785), .C1(new_n882), .C2(new_n884), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n750), .B(KEYINPUT57), .Z(new_n907));
  AND3_X1   g721(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n883), .B1(new_n882), .B2(new_n884), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n906), .B1(new_n910), .B2(new_n706), .ZN(new_n911));
  OAI21_X1  g725(.A(KEYINPUT123), .B1(new_n911), .B2(new_n895), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n913));
  INV_X1    g727(.A(new_n895), .ZN(new_n914));
  INV_X1    g728(.A(new_n706), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n886), .B2(new_n907), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n913), .B(new_n914), .C1(new_n916), .C2(new_n906), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n912), .A2(new_n917), .ZN(G54));
  AND2_X1   g732(.A1(KEYINPUT58), .A2(G475), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n899), .A2(new_n641), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n641), .B1(new_n899), .B2(new_n919), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n920), .A2(new_n921), .A3(new_n895), .ZN(G60));
  NAND2_X1  g736(.A1(G478), .A2(G902), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT59), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n923), .A2(KEYINPUT59), .ZN(new_n925));
  AOI22_X1  g739(.A1(new_n881), .A2(new_n885), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n622), .A2(new_n623), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n914), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(KEYINPUT124), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n926), .A2(new_n931), .A3(new_n927), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n928), .B1(new_n930), .B2(new_n932), .ZN(G63));
  NAND2_X1  g747(.A1(new_n882), .A2(new_n884), .ZN(new_n934));
  NAND2_X1  g748(.A1(G217), .A2(G902), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT60), .Z(new_n936));
  NAND4_X1  g750(.A1(new_n934), .A2(new_n653), .A3(new_n654), .A4(new_n936), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n934), .A2(new_n936), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n380), .B(KEYINPUT125), .Z(new_n939));
  OAI211_X1 g753(.A(new_n914), .B(new_n937), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(G66));
  INV_X1    g756(.A(G224), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n561), .A2(new_n943), .A3(new_n279), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n856), .A2(new_n857), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n944), .B1(new_n945), .B2(new_n279), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n896), .B1(G898), .B2(new_n279), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(G69));
  AOI21_X1  g762(.A(new_n279), .B1(G227), .B2(G900), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n287), .A2(new_n294), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n542), .B(KEYINPUT126), .Z(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n767), .A2(new_n679), .A3(new_n768), .A4(new_n851), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n794), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n954), .A2(new_n800), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n742), .A2(new_n675), .A3(new_n698), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n695), .A2(new_n956), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n955), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n952), .B1(new_n960), .B2(new_n279), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(KEYINPUT127), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(G900), .A2(G953), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n794), .A2(new_n770), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n792), .A2(new_n726), .A3(new_n683), .A4(new_n828), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n800), .A2(new_n764), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n965), .A2(new_n956), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n952), .B(new_n964), .C1(new_n968), .C2(G953), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n969), .B1(new_n961), .B2(KEYINPUT127), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n949), .B1(new_n963), .B2(new_n970), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n961), .A2(KEYINPUT127), .ZN(new_n972));
  INV_X1    g786(.A(new_n949), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n972), .A2(new_n973), .A3(new_n962), .A4(new_n969), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n971), .A2(new_n974), .ZN(G72));
  NAND2_X1  g789(.A1(G472), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT63), .Z(new_n977));
  INV_X1    g791(.A(new_n945), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n977), .B1(new_n960), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n979), .A2(new_n296), .A3(new_n284), .ZN(new_n980));
  INV_X1    g794(.A(new_n297), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n296), .A2(new_n284), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n934), .A2(new_n981), .A3(new_n982), .A4(new_n977), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n977), .B1(new_n968), .B2(new_n978), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n895), .B1(new_n984), .B2(new_n297), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n980), .A2(new_n983), .A3(new_n985), .ZN(G57));
endmodule


