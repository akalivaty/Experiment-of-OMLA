

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U558 ( .A1(n534), .A2(G2105), .ZN(n531) );
  XOR2_X2 U559 ( .A(n544), .B(n543), .Z(n527) );
  AND2_X1 U560 ( .A1(n685), .A2(n822), .ZN(n686) );
  INV_X1 U561 ( .A(KEYINPUT64), .ZN(n760) );
  XOR2_X1 U562 ( .A(KEYINPUT27), .B(n706), .Z(n528) );
  XOR2_X1 U563 ( .A(n541), .B(KEYINPUT23), .Z(n529) );
  NOR2_X1 U564 ( .A1(n703), .A2(n933), .ZN(n698) );
  NOR2_X1 U565 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U566 ( .A1(G164), .A2(G1384), .ZN(n822) );
  AND2_X1 U567 ( .A1(n835), .A2(n834), .ZN(n836) );
  NOR2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n530) );
  XOR2_X2 U569 ( .A(KEYINPUT17), .B(n530), .Z(n904) );
  NAND2_X1 U570 ( .A1(n904), .A2(G138), .ZN(n533) );
  INV_X1 U571 ( .A(G2104), .ZN(n534) );
  XNOR2_X2 U572 ( .A(n531), .B(KEYINPUT66), .ZN(n901) );
  NAND2_X1 U573 ( .A1(G102), .A2(n901), .ZN(n532) );
  NAND2_X1 U574 ( .A1(n533), .A2(n532), .ZN(n538) );
  AND2_X1 U575 ( .A1(n534), .A2(G2105), .ZN(n896) );
  NAND2_X1 U576 ( .A1(G126), .A2(n896), .ZN(n536) );
  AND2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n897) );
  NAND2_X1 U578 ( .A1(G114), .A2(n897), .ZN(n535) );
  NAND2_X1 U579 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U580 ( .A1(n538), .A2(n537), .ZN(G164) );
  NAND2_X1 U581 ( .A1(n897), .A2(G113), .ZN(n540) );
  NAND2_X1 U582 ( .A1(n904), .A2(G137), .ZN(n539) );
  AND2_X1 U583 ( .A1(n540), .A2(n539), .ZN(n684) );
  INV_X1 U584 ( .A(KEYINPUT67), .ZN(n544) );
  NAND2_X1 U585 ( .A1(G101), .A2(n901), .ZN(n541) );
  NAND2_X1 U586 ( .A1(n896), .A2(G125), .ZN(n542) );
  NAND2_X1 U587 ( .A1(n529), .A2(n542), .ZN(n543) );
  AND2_X1 U588 ( .A1(n684), .A2(n527), .ZN(G160) );
  XOR2_X1 U589 ( .A(G543), .B(KEYINPUT0), .Z(n632) );
  NOR2_X1 U590 ( .A1(G651), .A2(n632), .ZN(n545) );
  XOR2_X1 U591 ( .A(KEYINPUT65), .B(n545), .Z(n648) );
  NAND2_X1 U592 ( .A1(G47), .A2(n648), .ZN(n548) );
  INV_X1 U593 ( .A(G651), .ZN(n549) );
  NOR2_X1 U594 ( .A1(G543), .A2(n549), .ZN(n546) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n546), .Z(n653) );
  NAND2_X1 U596 ( .A1(G60), .A2(n653), .ZN(n547) );
  NAND2_X1 U597 ( .A1(n548), .A2(n547), .ZN(n553) );
  NOR2_X1 U598 ( .A1(n632), .A2(n549), .ZN(n649) );
  NAND2_X1 U599 ( .A1(G72), .A2(n649), .ZN(n551) );
  NOR2_X1 U600 ( .A1(G651), .A2(G543), .ZN(n650) );
  NAND2_X1 U601 ( .A1(G85), .A2(n650), .ZN(n550) );
  NAND2_X1 U602 ( .A1(n551), .A2(n550), .ZN(n552) );
  OR2_X1 U603 ( .A1(n553), .A2(n552), .ZN(G290) );
  NAND2_X1 U604 ( .A1(G52), .A2(n648), .ZN(n555) );
  NAND2_X1 U605 ( .A1(G64), .A2(n653), .ZN(n554) );
  NAND2_X1 U606 ( .A1(n555), .A2(n554), .ZN(n560) );
  NAND2_X1 U607 ( .A1(G77), .A2(n649), .ZN(n557) );
  NAND2_X1 U608 ( .A1(G90), .A2(n650), .ZN(n556) );
  NAND2_X1 U609 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U610 ( .A(KEYINPUT9), .B(n558), .Z(n559) );
  NOR2_X1 U611 ( .A1(n560), .A2(n559), .ZN(G171) );
  AND2_X1 U612 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U613 ( .A(G132), .ZN(G219) );
  INV_X1 U614 ( .A(G82), .ZN(G220) );
  INV_X1 U615 ( .A(G120), .ZN(G236) );
  NAND2_X1 U616 ( .A1(n650), .A2(G89), .ZN(n561) );
  XNOR2_X1 U617 ( .A(n561), .B(KEYINPUT4), .ZN(n563) );
  NAND2_X1 U618 ( .A1(G76), .A2(n649), .ZN(n562) );
  NAND2_X1 U619 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U620 ( .A(n564), .B(KEYINPUT5), .ZN(n570) );
  NAND2_X1 U621 ( .A1(n653), .A2(G63), .ZN(n565) );
  XNOR2_X1 U622 ( .A(n565), .B(KEYINPUT72), .ZN(n567) );
  NAND2_X1 U623 ( .A1(G51), .A2(n648), .ZN(n566) );
  NAND2_X1 U624 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U625 ( .A(KEYINPUT6), .B(n568), .Z(n569) );
  NAND2_X1 U626 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U627 ( .A(n571), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U628 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U629 ( .A1(G7), .A2(G661), .ZN(n572) );
  XNOR2_X1 U630 ( .A(n572), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U631 ( .A(G223), .ZN(n837) );
  NAND2_X1 U632 ( .A1(n837), .A2(G567), .ZN(n573) );
  XOR2_X1 U633 ( .A(KEYINPUT11), .B(n573), .Z(G234) );
  XOR2_X1 U634 ( .A(G860), .B(KEYINPUT70), .Z(n604) );
  NAND2_X1 U635 ( .A1(n653), .A2(G56), .ZN(n574) );
  XNOR2_X1 U636 ( .A(n574), .B(KEYINPUT14), .ZN(n576) );
  NAND2_X1 U637 ( .A1(G43), .A2(n648), .ZN(n575) );
  NAND2_X1 U638 ( .A1(n576), .A2(n575), .ZN(n583) );
  NAND2_X1 U639 ( .A1(n650), .A2(G81), .ZN(n577) );
  XNOR2_X1 U640 ( .A(n577), .B(KEYINPUT12), .ZN(n579) );
  NAND2_X1 U641 ( .A1(G68), .A2(n649), .ZN(n578) );
  NAND2_X1 U642 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT69), .B(n580), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT13), .B(n581), .ZN(n582) );
  NOR2_X1 U645 ( .A1(n583), .A2(n582), .ZN(n954) );
  INV_X1 U646 ( .A(n954), .ZN(n610) );
  OR2_X1 U647 ( .A1(n604), .A2(n610), .ZN(G153) );
  INV_X1 U648 ( .A(G171), .ZN(G301) );
  NAND2_X1 U649 ( .A1(G868), .A2(G301), .ZN(n593) );
  NAND2_X1 U650 ( .A1(G79), .A2(n649), .ZN(n585) );
  NAND2_X1 U651 ( .A1(G54), .A2(n648), .ZN(n584) );
  NAND2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n590) );
  NAND2_X1 U653 ( .A1(G66), .A2(n653), .ZN(n587) );
  NAND2_X1 U654 ( .A1(G92), .A2(n650), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U656 ( .A(KEYINPUT71), .B(n588), .Z(n589) );
  NOR2_X1 U657 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U658 ( .A(KEYINPUT15), .B(n591), .ZN(n933) );
  INV_X1 U659 ( .A(G868), .ZN(n667) );
  NAND2_X1 U660 ( .A1(n933), .A2(n667), .ZN(n592) );
  NAND2_X1 U661 ( .A1(n593), .A2(n592), .ZN(G284) );
  NAND2_X1 U662 ( .A1(G78), .A2(n649), .ZN(n595) );
  NAND2_X1 U663 ( .A1(G91), .A2(n650), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U665 ( .A1(n648), .A2(G53), .ZN(n596) );
  XOR2_X1 U666 ( .A(KEYINPUT68), .B(n596), .Z(n597) );
  NOR2_X1 U667 ( .A1(n598), .A2(n597), .ZN(n600) );
  NAND2_X1 U668 ( .A1(n653), .A2(G65), .ZN(n599) );
  NAND2_X1 U669 ( .A1(n600), .A2(n599), .ZN(G299) );
  INV_X1 U670 ( .A(G299), .ZN(n712) );
  NAND2_X1 U671 ( .A1(n712), .A2(n667), .ZN(n601) );
  XNOR2_X1 U672 ( .A(n601), .B(KEYINPUT73), .ZN(n603) );
  NOR2_X1 U673 ( .A1(n667), .A2(G286), .ZN(n602) );
  NOR2_X1 U674 ( .A1(n603), .A2(n602), .ZN(G297) );
  NAND2_X1 U675 ( .A1(n604), .A2(G559), .ZN(n605) );
  INV_X1 U676 ( .A(n933), .ZN(n647) );
  NAND2_X1 U677 ( .A1(n605), .A2(n647), .ZN(n606) );
  XNOR2_X1 U678 ( .A(n606), .B(KEYINPUT74), .ZN(n607) );
  XNOR2_X1 U679 ( .A(KEYINPUT16), .B(n607), .ZN(G148) );
  NOR2_X1 U680 ( .A1(G559), .A2(n667), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n647), .A2(n608), .ZN(n609) );
  XNOR2_X1 U682 ( .A(n609), .B(KEYINPUT75), .ZN(n612) );
  NOR2_X1 U683 ( .A1(n610), .A2(G868), .ZN(n611) );
  NOR2_X1 U684 ( .A1(n612), .A2(n611), .ZN(G282) );
  NAND2_X1 U685 ( .A1(G123), .A2(n896), .ZN(n613) );
  XNOR2_X1 U686 ( .A(n613), .B(KEYINPUT18), .ZN(n614) );
  XNOR2_X1 U687 ( .A(n614), .B(KEYINPUT76), .ZN(n616) );
  NAND2_X1 U688 ( .A1(G111), .A2(n897), .ZN(n615) );
  NAND2_X1 U689 ( .A1(n616), .A2(n615), .ZN(n620) );
  NAND2_X1 U690 ( .A1(n904), .A2(G135), .ZN(n618) );
  NAND2_X1 U691 ( .A1(G99), .A2(n901), .ZN(n617) );
  NAND2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n1012) );
  XNOR2_X1 U694 ( .A(n1012), .B(G2096), .ZN(n622) );
  INV_X1 U695 ( .A(G2100), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n622), .A2(n621), .ZN(G156) );
  NAND2_X1 U697 ( .A1(G73), .A2(n649), .ZN(n623) );
  XNOR2_X1 U698 ( .A(n623), .B(KEYINPUT2), .ZN(n625) );
  NAND2_X1 U699 ( .A1(n653), .A2(G61), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U701 ( .A1(G48), .A2(n648), .ZN(n626) );
  XNOR2_X1 U702 ( .A(KEYINPUT81), .B(n626), .ZN(n627) );
  NOR2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U704 ( .A1(n650), .A2(G86), .ZN(n629) );
  NAND2_X1 U705 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U706 ( .A(KEYINPUT82), .B(n631), .ZN(G305) );
  NAND2_X1 U707 ( .A1(G74), .A2(G651), .ZN(n637) );
  NAND2_X1 U708 ( .A1(G49), .A2(n648), .ZN(n634) );
  NAND2_X1 U709 ( .A1(G87), .A2(n632), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U711 ( .A1(n653), .A2(n635), .ZN(n636) );
  NAND2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U713 ( .A(n638), .B(KEYINPUT80), .ZN(G288) );
  NAND2_X1 U714 ( .A1(G75), .A2(n649), .ZN(n640) );
  NAND2_X1 U715 ( .A1(G88), .A2(n650), .ZN(n639) );
  NAND2_X1 U716 ( .A1(n640), .A2(n639), .ZN(n645) );
  NAND2_X1 U717 ( .A1(G50), .A2(n648), .ZN(n642) );
  NAND2_X1 U718 ( .A1(G62), .A2(n653), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U720 ( .A(KEYINPUT83), .B(n643), .Z(n644) );
  NOR2_X1 U721 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U722 ( .A(KEYINPUT84), .B(n646), .ZN(G166) );
  INV_X1 U723 ( .A(G166), .ZN(G303) );
  NAND2_X1 U724 ( .A1(n647), .A2(G559), .ZN(n844) );
  NAND2_X1 U725 ( .A1(n648), .A2(G55), .ZN(n658) );
  NAND2_X1 U726 ( .A1(G80), .A2(n649), .ZN(n652) );
  NAND2_X1 U727 ( .A1(G93), .A2(n650), .ZN(n651) );
  NAND2_X1 U728 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U729 ( .A1(n653), .A2(G67), .ZN(n654) );
  XOR2_X1 U730 ( .A(KEYINPUT78), .B(n654), .Z(n655) );
  NOR2_X1 U731 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U732 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U733 ( .A(KEYINPUT79), .B(n659), .Z(n848) );
  XOR2_X1 U734 ( .A(n848), .B(G299), .Z(n661) );
  XNOR2_X1 U735 ( .A(G305), .B(n954), .ZN(n660) );
  XNOR2_X1 U736 ( .A(n661), .B(n660), .ZN(n665) );
  XNOR2_X1 U737 ( .A(G290), .B(KEYINPUT19), .ZN(n663) );
  XNOR2_X1 U738 ( .A(G288), .B(G303), .ZN(n662) );
  XNOR2_X1 U739 ( .A(n663), .B(n662), .ZN(n664) );
  XOR2_X1 U740 ( .A(n665), .B(n664), .Z(n911) );
  XNOR2_X1 U741 ( .A(n844), .B(n911), .ZN(n666) );
  NAND2_X1 U742 ( .A1(n666), .A2(G868), .ZN(n669) );
  NAND2_X1 U743 ( .A1(n667), .A2(n848), .ZN(n668) );
  NAND2_X1 U744 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U745 ( .A1(G2078), .A2(G2084), .ZN(n670) );
  XOR2_X1 U746 ( .A(KEYINPUT20), .B(n670), .Z(n671) );
  NAND2_X1 U747 ( .A1(G2090), .A2(n671), .ZN(n672) );
  XNOR2_X1 U748 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U749 ( .A1(n673), .A2(G2072), .ZN(n674) );
  XOR2_X1 U750 ( .A(KEYINPUT85), .B(n674), .Z(G158) );
  XNOR2_X1 U751 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U752 ( .A1(G69), .A2(G57), .ZN(n675) );
  NOR2_X1 U753 ( .A1(G236), .A2(n675), .ZN(n676) );
  XNOR2_X1 U754 ( .A(KEYINPUT86), .B(n676), .ZN(n677) );
  NAND2_X1 U755 ( .A1(n677), .A2(G108), .ZN(n842) );
  NAND2_X1 U756 ( .A1(n842), .A2(G567), .ZN(n682) );
  NOR2_X1 U757 ( .A1(G220), .A2(G219), .ZN(n678) );
  XOR2_X1 U758 ( .A(KEYINPUT22), .B(n678), .Z(n679) );
  NOR2_X1 U759 ( .A1(G218), .A2(n679), .ZN(n680) );
  NAND2_X1 U760 ( .A1(G96), .A2(n680), .ZN(n843) );
  NAND2_X1 U761 ( .A1(n843), .A2(G2106), .ZN(n681) );
  NAND2_X1 U762 ( .A1(n682), .A2(n681), .ZN(n849) );
  NAND2_X1 U763 ( .A1(G483), .A2(G661), .ZN(n683) );
  NOR2_X1 U764 ( .A1(n849), .A2(n683), .ZN(n839) );
  NAND2_X1 U765 ( .A1(n839), .A2(G36), .ZN(G176) );
  AND2_X1 U766 ( .A1(n684), .A2(G40), .ZN(n685) );
  NAND2_X2 U767 ( .A1(n527), .A2(n686), .ZN(n732) );
  NAND2_X1 U768 ( .A1(G8), .A2(n732), .ZN(n780) );
  NOR2_X1 U769 ( .A1(G1981), .A2(G305), .ZN(n687) );
  XOR2_X1 U770 ( .A(n687), .B(KEYINPUT24), .Z(n688) );
  NOR2_X1 U771 ( .A1(n780), .A2(n688), .ZN(n773) );
  INV_X1 U772 ( .A(KEYINPUT95), .ZN(n690) );
  AND2_X1 U773 ( .A1(G1341), .A2(n732), .ZN(n689) );
  XNOR2_X1 U774 ( .A(n690), .B(n689), .ZN(n696) );
  INV_X1 U775 ( .A(n732), .ZN(n691) );
  NAND2_X1 U776 ( .A1(n691), .A2(G1996), .ZN(n693) );
  XNOR2_X1 U777 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n692) );
  XNOR2_X1 U778 ( .A(n693), .B(n692), .ZN(n694) );
  INV_X1 U779 ( .A(n694), .ZN(n695) );
  NOR2_X1 U780 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U781 ( .A1(n697), .A2(n954), .ZN(n703) );
  XOR2_X1 U782 ( .A(n698), .B(KEYINPUT96), .Z(n702) );
  NOR2_X1 U783 ( .A1(G2067), .A2(n732), .ZN(n700) );
  INV_X1 U784 ( .A(n732), .ZN(n717) );
  NOR2_X1 U785 ( .A1(n717), .A2(G1348), .ZN(n699) );
  NOR2_X1 U786 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U787 ( .A1(n702), .A2(n701), .ZN(n705) );
  NAND2_X1 U788 ( .A1(n933), .A2(n703), .ZN(n704) );
  NAND2_X1 U789 ( .A1(n705), .A2(n704), .ZN(n710) );
  NAND2_X1 U790 ( .A1(n732), .A2(G1956), .ZN(n707) );
  NAND2_X1 U791 ( .A1(n717), .A2(G2072), .ZN(n706) );
  NAND2_X1 U792 ( .A1(n707), .A2(n528), .ZN(n708) );
  XNOR2_X1 U793 ( .A(n708), .B(KEYINPUT93), .ZN(n711) );
  NAND2_X1 U794 ( .A1(n712), .A2(n711), .ZN(n709) );
  NAND2_X1 U795 ( .A1(n710), .A2(n709), .ZN(n715) );
  NOR2_X1 U796 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U797 ( .A(n713), .B(KEYINPUT28), .Z(n714) );
  NAND2_X1 U798 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U799 ( .A(n716), .B(KEYINPUT29), .ZN(n721) );
  XNOR2_X1 U800 ( .A(G2078), .B(KEYINPUT25), .ZN(n960) );
  NOR2_X1 U801 ( .A1(n732), .A2(n960), .ZN(n719) );
  INV_X1 U802 ( .A(G1961), .ZN(n934) );
  NOR2_X1 U803 ( .A1(n717), .A2(n934), .ZN(n718) );
  NOR2_X1 U804 ( .A1(n719), .A2(n718), .ZN(n728) );
  AND2_X1 U805 ( .A1(G171), .A2(n728), .ZN(n720) );
  NOR2_X1 U806 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U807 ( .A(n722), .B(KEYINPUT97), .ZN(n747) );
  NOR2_X1 U808 ( .A1(G1966), .A2(n780), .ZN(n750) );
  NOR2_X1 U809 ( .A1(G2084), .A2(n732), .ZN(n746) );
  NOR2_X1 U810 ( .A1(n750), .A2(n746), .ZN(n723) );
  NAND2_X1 U811 ( .A1(G8), .A2(n723), .ZN(n724) );
  XNOR2_X1 U812 ( .A(KEYINPUT99), .B(n724), .ZN(n726) );
  XOR2_X1 U813 ( .A(KEYINPUT30), .B(KEYINPUT98), .Z(n725) );
  XNOR2_X1 U814 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U815 ( .A1(G168), .A2(n727), .ZN(n730) );
  NOR2_X1 U816 ( .A1(G171), .A2(n728), .ZN(n729) );
  NOR2_X1 U817 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U818 ( .A(KEYINPUT31), .B(n731), .Z(n748) );
  INV_X1 U819 ( .A(G8), .ZN(n739) );
  NOR2_X1 U820 ( .A1(G1971), .A2(n780), .ZN(n734) );
  NOR2_X1 U821 ( .A1(G2090), .A2(n732), .ZN(n733) );
  NOR2_X1 U822 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U823 ( .A(KEYINPUT100), .B(n735), .Z(n736) );
  NOR2_X1 U824 ( .A1(G166), .A2(n736), .ZN(n737) );
  XNOR2_X1 U825 ( .A(n737), .B(KEYINPUT101), .ZN(n738) );
  OR2_X1 U826 ( .A1(n739), .A2(n738), .ZN(n741) );
  AND2_X1 U827 ( .A1(n748), .A2(n741), .ZN(n740) );
  NAND2_X1 U828 ( .A1(n747), .A2(n740), .ZN(n744) );
  INV_X1 U829 ( .A(n741), .ZN(n742) );
  OR2_X1 U830 ( .A1(n742), .A2(G286), .ZN(n743) );
  NAND2_X1 U831 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U832 ( .A(n745), .B(KEYINPUT32), .ZN(n774) );
  INV_X1 U833 ( .A(n780), .ZN(n764) );
  AND2_X1 U834 ( .A1(n774), .A2(n764), .ZN(n754) );
  NAND2_X1 U835 ( .A1(G8), .A2(n746), .ZN(n752) );
  AND2_X1 U836 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U837 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U838 ( .A1(n752), .A2(n751), .ZN(n775) );
  NAND2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n938) );
  AND2_X1 U840 ( .A1(n775), .A2(n938), .ZN(n753) );
  NAND2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n759) );
  INV_X1 U842 ( .A(n938), .ZN(n756) );
  NOR2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n763) );
  NOR2_X1 U844 ( .A1(G1971), .A2(G303), .ZN(n755) );
  NOR2_X1 U845 ( .A1(n763), .A2(n755), .ZN(n947) );
  OR2_X1 U846 ( .A1(n756), .A2(n947), .ZN(n757) );
  OR2_X1 U847 ( .A1(n780), .A2(n757), .ZN(n758) );
  NAND2_X1 U848 ( .A1(n759), .A2(n758), .ZN(n761) );
  XNOR2_X1 U849 ( .A(n761), .B(n760), .ZN(n762) );
  INV_X1 U850 ( .A(KEYINPUT33), .ZN(n766) );
  NAND2_X1 U851 ( .A1(n762), .A2(n766), .ZN(n771) );
  XNOR2_X1 U852 ( .A(G1981), .B(G305), .ZN(n950) );
  INV_X1 U853 ( .A(n950), .ZN(n769) );
  NAND2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n767) );
  XOR2_X1 U856 ( .A(n767), .B(KEYINPUT102), .Z(n768) );
  AND2_X1 U857 ( .A1(n769), .A2(n768), .ZN(n770) );
  AND2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U859 ( .A1(n773), .A2(n772), .ZN(n826) );
  AND2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n778) );
  NAND2_X1 U861 ( .A1(G166), .A2(G8), .ZN(n776) );
  NOR2_X1 U862 ( .A1(G2090), .A2(n776), .ZN(n777) );
  XNOR2_X1 U863 ( .A(n779), .B(KEYINPUT103), .ZN(n781) );
  NAND2_X1 U864 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U865 ( .A(n782), .B(KEYINPUT104), .ZN(n824) );
  XNOR2_X1 U866 ( .A(G2067), .B(KEYINPUT37), .ZN(n819) );
  XNOR2_X1 U867 ( .A(KEYINPUT36), .B(KEYINPUT88), .ZN(n793) );
  NAND2_X1 U868 ( .A1(G128), .A2(n896), .ZN(n784) );
  NAND2_X1 U869 ( .A1(G116), .A2(n897), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U871 ( .A(n785), .B(KEYINPUT35), .ZN(n791) );
  XNOR2_X1 U872 ( .A(KEYINPUT34), .B(KEYINPUT87), .ZN(n789) );
  NAND2_X1 U873 ( .A1(n904), .A2(G140), .ZN(n787) );
  NAND2_X1 U874 ( .A1(G104), .A2(n901), .ZN(n786) );
  NAND2_X1 U875 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U876 ( .A(n789), .B(n788), .ZN(n790) );
  NAND2_X1 U877 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U878 ( .A(n793), .B(n792), .Z(n879) );
  NOR2_X1 U879 ( .A1(n819), .A2(n879), .ZN(n1017) );
  NAND2_X1 U880 ( .A1(G129), .A2(n896), .ZN(n795) );
  NAND2_X1 U881 ( .A1(G117), .A2(n897), .ZN(n794) );
  NAND2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n800) );
  XOR2_X1 U883 ( .A(KEYINPUT91), .B(KEYINPUT38), .Z(n797) );
  NAND2_X1 U884 ( .A1(G105), .A2(n901), .ZN(n796) );
  XNOR2_X1 U885 ( .A(n797), .B(n796), .ZN(n798) );
  XOR2_X1 U886 ( .A(KEYINPUT90), .B(n798), .Z(n799) );
  NOR2_X1 U887 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U888 ( .A(n801), .B(KEYINPUT92), .ZN(n803) );
  NAND2_X1 U889 ( .A1(G141), .A2(n904), .ZN(n802) );
  NAND2_X1 U890 ( .A1(n803), .A2(n802), .ZN(n886) );
  NOR2_X1 U891 ( .A1(G1996), .A2(n886), .ZN(n1028) );
  NAND2_X1 U892 ( .A1(G119), .A2(n896), .ZN(n805) );
  NAND2_X1 U893 ( .A1(G131), .A2(n904), .ZN(n804) );
  NAND2_X1 U894 ( .A1(n805), .A2(n804), .ZN(n809) );
  NAND2_X1 U895 ( .A1(n897), .A2(G107), .ZN(n807) );
  NAND2_X1 U896 ( .A1(G95), .A2(n901), .ZN(n806) );
  NAND2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n808) );
  OR2_X1 U898 ( .A1(n809), .A2(n808), .ZN(n878) );
  NAND2_X1 U899 ( .A1(G1991), .A2(n878), .ZN(n810) );
  XOR2_X1 U900 ( .A(KEYINPUT89), .B(n810), .Z(n812) );
  NAND2_X1 U901 ( .A1(G1996), .A2(n886), .ZN(n811) );
  NAND2_X1 U902 ( .A1(n812), .A2(n811), .ZN(n1011) );
  NOR2_X1 U903 ( .A1(G1986), .A2(G290), .ZN(n813) );
  NOR2_X1 U904 ( .A1(G1991), .A2(n878), .ZN(n1013) );
  NOR2_X1 U905 ( .A1(n813), .A2(n1013), .ZN(n814) );
  NOR2_X1 U906 ( .A1(n1011), .A2(n814), .ZN(n815) );
  NOR2_X1 U907 ( .A1(n1028), .A2(n815), .ZN(n816) );
  XOR2_X1 U908 ( .A(KEYINPUT39), .B(n816), .Z(n817) );
  NOR2_X1 U909 ( .A1(n1017), .A2(n817), .ZN(n818) );
  XNOR2_X1 U910 ( .A(n818), .B(KEYINPUT105), .ZN(n820) );
  NAND2_X1 U911 ( .A1(n879), .A2(n819), .ZN(n1014) );
  NAND2_X1 U912 ( .A1(n820), .A2(n1014), .ZN(n823) );
  NAND2_X1 U913 ( .A1(G160), .A2(G40), .ZN(n821) );
  NOR2_X1 U914 ( .A1(n822), .A2(n821), .ZN(n830) );
  NAND2_X1 U915 ( .A1(n823), .A2(n830), .ZN(n827) );
  AND2_X1 U916 ( .A1(n824), .A2(n827), .ZN(n825) );
  NAND2_X1 U917 ( .A1(n826), .A2(n825), .ZN(n835) );
  INV_X1 U918 ( .A(n827), .ZN(n833) );
  XNOR2_X1 U919 ( .A(G1986), .B(G290), .ZN(n941) );
  NOR2_X1 U920 ( .A1(n1011), .A2(n941), .ZN(n829) );
  INV_X1 U921 ( .A(n1017), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n829), .A2(n828), .ZN(n831) );
  NAND2_X1 U923 ( .A1(n831), .A2(n830), .ZN(n832) );
  OR2_X1 U924 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U925 ( .A(n836), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U928 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G1), .A2(G3), .ZN(n840) );
  NAND2_X1 U930 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U931 ( .A(n841), .B(KEYINPUT108), .ZN(G188) );
  XNOR2_X1 U932 ( .A(G69), .B(KEYINPUT109), .ZN(G235) );
  INV_X1 U934 ( .A(G108), .ZN(G238) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  INV_X1 U936 ( .A(G57), .ZN(G237) );
  NOR2_X1 U937 ( .A1(n843), .A2(n842), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U939 ( .A(n954), .B(KEYINPUT77), .ZN(n845) );
  XNOR2_X1 U940 ( .A(n845), .B(n844), .ZN(n846) );
  NOR2_X1 U941 ( .A1(G860), .A2(n846), .ZN(n847) );
  XOR2_X1 U942 ( .A(n848), .B(n847), .Z(G145) );
  INV_X1 U943 ( .A(n849), .ZN(G319) );
  XNOR2_X1 U944 ( .A(G1976), .B(KEYINPUT41), .ZN(n859) );
  XOR2_X1 U945 ( .A(G1986), .B(G1961), .Z(n851) );
  XNOR2_X1 U946 ( .A(G1981), .B(G1971), .ZN(n850) );
  XNOR2_X1 U947 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U948 ( .A(G1991), .B(G1956), .Z(n853) );
  XNOR2_X1 U949 ( .A(G1966), .B(G1996), .ZN(n852) );
  XNOR2_X1 U950 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U951 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U952 ( .A(KEYINPUT112), .B(G2474), .ZN(n856) );
  XNOR2_X1 U953 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U954 ( .A(n859), .B(n858), .ZN(G229) );
  XOR2_X1 U955 ( .A(KEYINPUT43), .B(KEYINPUT111), .Z(n861) );
  XNOR2_X1 U956 ( .A(KEYINPUT110), .B(G2678), .ZN(n860) );
  XNOR2_X1 U957 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U958 ( .A(KEYINPUT42), .B(G2090), .Z(n863) );
  XNOR2_X1 U959 ( .A(G2067), .B(G2072), .ZN(n862) );
  XNOR2_X1 U960 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U961 ( .A(n865), .B(n864), .Z(n867) );
  XNOR2_X1 U962 ( .A(G2096), .B(G2100), .ZN(n866) );
  XNOR2_X1 U963 ( .A(n867), .B(n866), .ZN(n869) );
  XOR2_X1 U964 ( .A(G2078), .B(G2084), .Z(n868) );
  XNOR2_X1 U965 ( .A(n869), .B(n868), .ZN(G227) );
  NAND2_X1 U966 ( .A1(G124), .A2(n896), .ZN(n870) );
  XOR2_X1 U967 ( .A(KEYINPUT113), .B(n870), .Z(n871) );
  XNOR2_X1 U968 ( .A(n871), .B(KEYINPUT44), .ZN(n873) );
  NAND2_X1 U969 ( .A1(G112), .A2(n897), .ZN(n872) );
  NAND2_X1 U970 ( .A1(n873), .A2(n872), .ZN(n877) );
  NAND2_X1 U971 ( .A1(n904), .A2(G136), .ZN(n875) );
  NAND2_X1 U972 ( .A1(G100), .A2(n901), .ZN(n874) );
  NAND2_X1 U973 ( .A1(n875), .A2(n874), .ZN(n876) );
  NOR2_X1 U974 ( .A1(n877), .A2(n876), .ZN(G162) );
  XNOR2_X1 U975 ( .A(G162), .B(n878), .ZN(n880) );
  XOR2_X1 U976 ( .A(n880), .B(n879), .Z(n881) );
  XOR2_X1 U977 ( .A(n881), .B(KEYINPUT48), .Z(n883) );
  XNOR2_X1 U978 ( .A(G164), .B(KEYINPUT46), .ZN(n882) );
  XNOR2_X1 U979 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U980 ( .A(G160), .B(n884), .Z(n885) );
  XNOR2_X1 U981 ( .A(n886), .B(n885), .ZN(n895) );
  NAND2_X1 U982 ( .A1(G130), .A2(n896), .ZN(n888) );
  NAND2_X1 U983 ( .A1(G118), .A2(n897), .ZN(n887) );
  NAND2_X1 U984 ( .A1(n888), .A2(n887), .ZN(n893) );
  NAND2_X1 U985 ( .A1(n904), .A2(G142), .ZN(n890) );
  NAND2_X1 U986 ( .A1(G106), .A2(n901), .ZN(n889) );
  NAND2_X1 U987 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U988 ( .A(KEYINPUT45), .B(n891), .Z(n892) );
  NOR2_X1 U989 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U990 ( .A(n895), .B(n894), .Z(n909) );
  NAND2_X1 U991 ( .A1(G127), .A2(n896), .ZN(n899) );
  NAND2_X1 U992 ( .A1(G115), .A2(n897), .ZN(n898) );
  NAND2_X1 U993 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U994 ( .A(n900), .B(KEYINPUT47), .ZN(n903) );
  NAND2_X1 U995 ( .A1(G103), .A2(n901), .ZN(n902) );
  NAND2_X1 U996 ( .A1(n903), .A2(n902), .ZN(n907) );
  NAND2_X1 U997 ( .A1(n904), .A2(G139), .ZN(n905) );
  XOR2_X1 U998 ( .A(KEYINPUT114), .B(n905), .Z(n906) );
  NOR2_X1 U999 ( .A1(n907), .A2(n906), .ZN(n1020) );
  XNOR2_X1 U1000 ( .A(n1020), .B(n1012), .ZN(n908) );
  XNOR2_X1 U1001 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n910), .ZN(G395) );
  XOR2_X1 U1003 ( .A(KEYINPUT115), .B(n911), .Z(n913) );
  XNOR2_X1 U1004 ( .A(G171), .B(G286), .ZN(n912) );
  XNOR2_X1 U1005 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1006 ( .A(n914), .B(n933), .ZN(n915) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n915), .ZN(G397) );
  XNOR2_X1 U1008 ( .A(G2451), .B(G2446), .ZN(n925) );
  XOR2_X1 U1009 ( .A(G2430), .B(G2443), .Z(n917) );
  XNOR2_X1 U1010 ( .A(G2454), .B(G2435), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(n917), .B(n916), .ZN(n921) );
  XOR2_X1 U1012 ( .A(G2438), .B(KEYINPUT106), .Z(n919) );
  XNOR2_X1 U1013 ( .A(G1348), .B(G1341), .ZN(n918) );
  XNOR2_X1 U1014 ( .A(n919), .B(n918), .ZN(n920) );
  XOR2_X1 U1015 ( .A(n921), .B(n920), .Z(n923) );
  XNOR2_X1 U1016 ( .A(KEYINPUT107), .B(G2427), .ZN(n922) );
  XNOR2_X1 U1017 ( .A(n923), .B(n922), .ZN(n924) );
  XNOR2_X1 U1018 ( .A(n925), .B(n924), .ZN(n926) );
  NAND2_X1 U1019 ( .A1(n926), .A2(G14), .ZN(n932) );
  NAND2_X1 U1020 ( .A1(G319), .A2(n932), .ZN(n929) );
  NOR2_X1 U1021 ( .A1(G229), .A2(G227), .ZN(n927) );
  XNOR2_X1 U1022 ( .A(KEYINPUT49), .B(n927), .ZN(n928) );
  NOR2_X1 U1023 ( .A1(n929), .A2(n928), .ZN(n931) );
  NOR2_X1 U1024 ( .A1(G395), .A2(G397), .ZN(n930) );
  NAND2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(G225) );
  INV_X1 U1026 ( .A(G225), .ZN(G308) );
  INV_X1 U1027 ( .A(n932), .ZN(G401) );
  XNOR2_X1 U1028 ( .A(G1348), .B(n933), .ZN(n945) );
  XNOR2_X1 U1029 ( .A(G171), .B(KEYINPUT122), .ZN(n935) );
  XNOR2_X1 U1030 ( .A(n935), .B(n934), .ZN(n937) );
  XNOR2_X1 U1031 ( .A(G1956), .B(G299), .ZN(n936) );
  NOR2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n939) );
  NAND2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n943) );
  NAND2_X1 U1035 ( .A1(G1971), .A2(G303), .ZN(n942) );
  NAND2_X1 U1036 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1037 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1038 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1039 ( .A(KEYINPUT123), .B(n948), .ZN(n953) );
  XOR2_X1 U1040 ( .A(G1966), .B(G168), .Z(n949) );
  NOR2_X1 U1041 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1042 ( .A(KEYINPUT57), .B(n951), .Z(n952) );
  NAND2_X1 U1043 ( .A1(n953), .A2(n952), .ZN(n956) );
  XOR2_X1 U1044 ( .A(n954), .B(G1341), .Z(n955) );
  NOR2_X1 U1045 ( .A1(n956), .A2(n955), .ZN(n958) );
  XOR2_X1 U1046 ( .A(G16), .B(KEYINPUT56), .Z(n957) );
  NOR2_X1 U1047 ( .A1(n958), .A2(n957), .ZN(n1040) );
  XNOR2_X1 U1048 ( .A(G2067), .B(KEYINPUT118), .ZN(n959) );
  XNOR2_X1 U1049 ( .A(n959), .B(G26), .ZN(n965) );
  XOR2_X1 U1050 ( .A(n960), .B(G27), .Z(n962) );
  XNOR2_X1 U1051 ( .A(G32), .B(G1996), .ZN(n961) );
  NOR2_X1 U1052 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1053 ( .A(KEYINPUT119), .B(n963), .ZN(n964) );
  NOR2_X1 U1054 ( .A1(n965), .A2(n964), .ZN(n970) );
  XOR2_X1 U1055 ( .A(G2072), .B(G33), .Z(n966) );
  NAND2_X1 U1056 ( .A1(n966), .A2(G28), .ZN(n968) );
  XNOR2_X1 U1057 ( .A(G25), .B(G1991), .ZN(n967) );
  NOR2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1059 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1060 ( .A(n971), .B(KEYINPUT120), .ZN(n972) );
  XNOR2_X1 U1061 ( .A(KEYINPUT53), .B(n972), .ZN(n978) );
  XOR2_X1 U1062 ( .A(KEYINPUT121), .B(G34), .Z(n974) );
  XNOR2_X1 U1063 ( .A(G2084), .B(KEYINPUT54), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(n974), .B(n973), .ZN(n976) );
  XNOR2_X1 U1065 ( .A(G35), .B(G2090), .ZN(n975) );
  NOR2_X1 U1066 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1067 ( .A1(n978), .A2(n977), .ZN(n1005) );
  NOR2_X1 U1068 ( .A1(G29), .A2(KEYINPUT55), .ZN(n979) );
  NAND2_X1 U1069 ( .A1(n1005), .A2(n979), .ZN(n980) );
  NAND2_X1 U1070 ( .A1(G11), .A2(n980), .ZN(n1009) );
  XOR2_X1 U1071 ( .A(G16), .B(KEYINPUT124), .Z(n1004) );
  XOR2_X1 U1072 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n987) );
  XNOR2_X1 U1073 ( .A(G1976), .B(G23), .ZN(n982) );
  XNOR2_X1 U1074 ( .A(G1971), .B(G22), .ZN(n981) );
  NOR2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n985) );
  XNOR2_X1 U1076 ( .A(G1986), .B(KEYINPUT125), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(n983), .B(G24), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(n987), .B(n986), .ZN(n991) );
  XNOR2_X1 U1080 ( .A(G1966), .B(G21), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(G1961), .B(G5), .ZN(n988) );
  NOR2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n1001) );
  XOR2_X1 U1084 ( .A(G1348), .B(KEYINPUT59), .Z(n992) );
  XNOR2_X1 U1085 ( .A(G4), .B(n992), .ZN(n994) );
  XNOR2_X1 U1086 ( .A(G20), .B(G1956), .ZN(n993) );
  NOR2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(G1981), .B(G6), .ZN(n996) );
  XNOR2_X1 U1089 ( .A(G1341), .B(G19), .ZN(n995) );
  NOR2_X1 U1090 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1092 ( .A(KEYINPUT60), .B(n999), .ZN(n1000) );
  NOR2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1094 ( .A(n1002), .B(KEYINPUT61), .ZN(n1003) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1007) );
  INV_X1 U1096 ( .A(KEYINPUT55), .ZN(n1034) );
  OR2_X1 U1097 ( .A1(n1034), .A2(n1005), .ZN(n1006) );
  NAND2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1038) );
  XOR2_X1 U1100 ( .A(G160), .B(G2084), .Z(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1019) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1026) );
  XOR2_X1 U1106 ( .A(G2072), .B(n1020), .Z(n1022) );
  XOR2_X1 U1107 ( .A(G164), .B(G2078), .Z(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1109 ( .A(KEYINPUT116), .B(n1023), .Z(n1024) );
  XNOR2_X1 U1110 ( .A(KEYINPUT50), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1031) );
  XOR2_X1 U1112 ( .A(G2090), .B(G162), .Z(n1027) );
  NOR2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1114 ( .A(KEYINPUT51), .B(n1029), .Z(n1030) );
  NAND2_X1 U1115 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1116 ( .A(n1032), .B(KEYINPUT52), .ZN(n1033) );
  XNOR2_X1 U1117 ( .A(KEYINPUT117), .B(n1033), .ZN(n1035) );
  NAND2_X1 U1118 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1119 ( .A1(n1036), .A2(G29), .ZN(n1037) );
  NAND2_X1 U1120 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NOR2_X1 U1121 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XOR2_X1 U1122 ( .A(KEYINPUT127), .B(n1041), .Z(n1042) );
  XNOR2_X1 U1123 ( .A(KEYINPUT62), .B(n1042), .ZN(G311) );
  INV_X1 U1124 ( .A(G311), .ZN(G150) );
endmodule

