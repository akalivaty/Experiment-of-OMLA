

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U325 ( .A(n396), .B(KEYINPUT48), .ZN(n541) );
  XNOR2_X1 U326 ( .A(n379), .B(n378), .ZN(n381) );
  XNOR2_X1 U327 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U328 ( .A(n441), .B(KEYINPUT55), .ZN(n456) );
  XNOR2_X1 U329 ( .A(n457), .B(G190GAT), .ZN(n458) );
  XNOR2_X1 U330 ( .A(n459), .B(n458), .ZN(G1351GAT) );
  XNOR2_X1 U331 ( .A(G36GAT), .B(G190GAT), .ZN(n293) );
  XNOR2_X1 U332 ( .A(n293), .B(G218GAT), .ZN(n323) );
  XNOR2_X1 U333 ( .A(G50GAT), .B(KEYINPUT80), .ZN(n294) );
  XOR2_X1 U334 ( .A(n294), .B(G162GAT), .Z(n436) );
  INV_X1 U335 ( .A(n436), .ZN(n295) );
  XOR2_X1 U336 ( .A(n323), .B(n295), .Z(n312) );
  XOR2_X1 U337 ( .A(KEYINPUT10), .B(G106GAT), .Z(n297) );
  XNOR2_X1 U338 ( .A(KEYINPUT81), .B(KEYINPUT66), .ZN(n296) );
  XNOR2_X1 U339 ( .A(n297), .B(n296), .ZN(n299) );
  INV_X1 U340 ( .A(KEYINPUT68), .ZN(n298) );
  XNOR2_X1 U341 ( .A(n299), .B(n298), .ZN(n301) );
  XOR2_X1 U342 ( .A(G99GAT), .B(G85GAT), .Z(n329) );
  XNOR2_X1 U343 ( .A(n329), .B(G92GAT), .ZN(n300) );
  XNOR2_X1 U344 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U345 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n303) );
  NAND2_X1 U346 ( .A1(G232GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U347 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U348 ( .A(n305), .B(n304), .Z(n310) );
  XOR2_X1 U349 ( .A(KEYINPUT71), .B(KEYINPUT7), .Z(n307) );
  XNOR2_X1 U350 ( .A(G43GAT), .B(G29GAT), .ZN(n306) );
  XNOR2_X1 U351 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U352 ( .A(KEYINPUT8), .B(n308), .Z(n359) );
  XNOR2_X1 U353 ( .A(n359), .B(G134GAT), .ZN(n309) );
  XNOR2_X1 U354 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U355 ( .A(n312), .B(n311), .Z(n535) );
  XOR2_X1 U356 ( .A(KEYINPUT90), .B(KEYINPUT17), .Z(n314) );
  XNOR2_X1 U357 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n313) );
  XNOR2_X1 U358 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U359 ( .A(G169GAT), .B(n315), .Z(n453) );
  XOR2_X1 U360 ( .A(G204GAT), .B(KEYINPUT78), .Z(n317) );
  XNOR2_X1 U361 ( .A(G176GAT), .B(G92GAT), .ZN(n316) );
  XNOR2_X1 U362 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U363 ( .A(G64GAT), .B(n318), .Z(n340) );
  XNOR2_X1 U364 ( .A(n453), .B(n340), .ZN(n327) );
  XOR2_X1 U365 ( .A(G197GAT), .B(KEYINPUT21), .Z(n428) );
  XNOR2_X1 U366 ( .A(G8GAT), .B(G183GAT), .ZN(n319) );
  XNOR2_X1 U367 ( .A(n319), .B(G211GAT), .ZN(n362) );
  XOR2_X1 U368 ( .A(n428), .B(n362), .Z(n321) );
  NAND2_X1 U369 ( .A1(G226GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U370 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U371 ( .A(n322), .B(KEYINPUT98), .Z(n325) );
  XNOR2_X1 U372 ( .A(n323), .B(KEYINPUT99), .ZN(n324) );
  XNOR2_X1 U373 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U374 ( .A(n327), .B(n326), .ZN(n513) );
  XNOR2_X1 U375 ( .A(KEYINPUT120), .B(n513), .ZN(n397) );
  XNOR2_X1 U376 ( .A(G106GAT), .B(KEYINPUT76), .ZN(n328) );
  XNOR2_X1 U377 ( .A(n328), .B(G148GAT), .ZN(n424) );
  XOR2_X1 U378 ( .A(KEYINPUT32), .B(n424), .Z(n331) );
  XNOR2_X1 U379 ( .A(n329), .B(G78GAT), .ZN(n330) );
  XNOR2_X1 U380 ( .A(n331), .B(n330), .ZN(n336) );
  XNOR2_X1 U381 ( .A(G71GAT), .B(G57GAT), .ZN(n332) );
  XNOR2_X1 U382 ( .A(n332), .B(KEYINPUT13), .ZN(n376) );
  XOR2_X1 U383 ( .A(n376), .B(KEYINPUT31), .Z(n334) );
  NAND2_X1 U384 ( .A1(G230GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U385 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U386 ( .A(n336), .B(n335), .Z(n342) );
  XOR2_X1 U387 ( .A(KEYINPUT77), .B(KEYINPUT79), .Z(n338) );
  XNOR2_X1 U388 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n337) );
  XNOR2_X1 U389 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U390 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U391 ( .A(n342), .B(n341), .ZN(n572) );
  XNOR2_X1 U392 ( .A(G113GAT), .B(G15GAT), .ZN(n344) );
  XNOR2_X1 U393 ( .A(G197GAT), .B(G22GAT), .ZN(n343) );
  XNOR2_X1 U394 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U395 ( .A(KEYINPUT75), .B(KEYINPUT70), .Z(n346) );
  XNOR2_X1 U396 ( .A(G141GAT), .B(KEYINPUT74), .ZN(n345) );
  XNOR2_X1 U397 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U398 ( .A(n348), .B(n347), .ZN(n353) );
  XOR2_X1 U399 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n350) );
  NAND2_X1 U400 ( .A1(G229GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U401 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U402 ( .A(KEYINPUT69), .B(n351), .ZN(n352) );
  XNOR2_X1 U403 ( .A(n353), .B(n352), .ZN(n358) );
  XOR2_X1 U404 ( .A(G50GAT), .B(G36GAT), .Z(n356) );
  XNOR2_X1 U405 ( .A(G1GAT), .B(KEYINPUT72), .ZN(n354) );
  XNOR2_X1 U406 ( .A(n354), .B(KEYINPUT73), .ZN(n365) );
  XNOR2_X1 U407 ( .A(G8GAT), .B(n365), .ZN(n355) );
  XNOR2_X1 U408 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U409 ( .A(n358), .B(n357), .Z(n361) );
  XNOR2_X1 U410 ( .A(G169GAT), .B(n359), .ZN(n360) );
  XOR2_X1 U411 ( .A(n361), .B(n360), .Z(n544) );
  INV_X1 U412 ( .A(n544), .ZN(n567) );
  XNOR2_X1 U413 ( .A(n362), .B(KEYINPUT84), .ZN(n364) );
  AND2_X1 U414 ( .A1(G231GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U415 ( .A(n364), .B(n363), .ZN(n369) );
  XOR2_X1 U416 ( .A(KEYINPUT88), .B(G64GAT), .Z(n367) );
  XOR2_X1 U417 ( .A(G15GAT), .B(G127GAT), .Z(n442) );
  XNOR2_X1 U418 ( .A(n365), .B(n442), .ZN(n366) );
  XNOR2_X1 U419 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U420 ( .A(n369), .B(n368), .ZN(n379) );
  XOR2_X1 U421 ( .A(KEYINPUT86), .B(KEYINPUT83), .Z(n371) );
  XNOR2_X1 U422 ( .A(KEYINPUT82), .B(KEYINPUT14), .ZN(n370) );
  XNOR2_X1 U423 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U424 ( .A(KEYINPUT12), .B(KEYINPUT87), .Z(n373) );
  XNOR2_X1 U425 ( .A(KEYINPUT85), .B(KEYINPUT15), .ZN(n372) );
  XNOR2_X1 U426 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U427 ( .A(n375), .B(n374), .Z(n377) );
  XNOR2_X1 U428 ( .A(G22GAT), .B(G155GAT), .ZN(n380) );
  XNOR2_X1 U429 ( .A(n380), .B(G78GAT), .ZN(n435) );
  XOR2_X1 U430 ( .A(n381), .B(n435), .Z(n550) );
  XOR2_X1 U431 ( .A(KEYINPUT36), .B(n535), .Z(n581) );
  NAND2_X1 U432 ( .A1(n550), .A2(n581), .ZN(n384) );
  XOR2_X1 U433 ( .A(KEYINPUT113), .B(KEYINPUT45), .Z(n382) );
  XNOR2_X1 U434 ( .A(KEYINPUT67), .B(n382), .ZN(n383) );
  XNOR2_X1 U435 ( .A(n384), .B(n383), .ZN(n385) );
  AND2_X1 U436 ( .A1(n567), .A2(n385), .ZN(n386) );
  NAND2_X1 U437 ( .A1(n572), .A2(n386), .ZN(n395) );
  XOR2_X1 U438 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n387) );
  XNOR2_X1 U439 ( .A(n572), .B(n387), .ZN(n559) );
  NOR2_X1 U440 ( .A1(n567), .A2(n559), .ZN(n388) );
  XNOR2_X1 U441 ( .A(n388), .B(KEYINPUT111), .ZN(n389) );
  XNOR2_X1 U442 ( .A(n389), .B(KEYINPUT46), .ZN(n390) );
  XOR2_X1 U443 ( .A(n550), .B(KEYINPUT110), .Z(n562) );
  NAND2_X1 U444 ( .A1(n390), .A2(n562), .ZN(n391) );
  INV_X1 U445 ( .A(n535), .ZN(n554) );
  NOR2_X1 U446 ( .A1(n391), .A2(n554), .ZN(n393) );
  XNOR2_X1 U447 ( .A(KEYINPUT47), .B(KEYINPUT112), .ZN(n392) );
  XNOR2_X1 U448 ( .A(n393), .B(n392), .ZN(n394) );
  NAND2_X1 U449 ( .A1(n395), .A2(n394), .ZN(n396) );
  NAND2_X1 U450 ( .A1(n397), .A2(n541), .ZN(n398) );
  XNOR2_X1 U451 ( .A(n398), .B(KEYINPUT54), .ZN(n399) );
  XNOR2_X1 U452 ( .A(n399), .B(KEYINPUT121), .ZN(n421) );
  XOR2_X1 U453 ( .A(G57GAT), .B(G85GAT), .Z(n401) );
  XNOR2_X1 U454 ( .A(G29GAT), .B(G162GAT), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U456 ( .A(G148GAT), .B(G155GAT), .Z(n403) );
  XNOR2_X1 U457 ( .A(G1GAT), .B(G127GAT), .ZN(n402) );
  XNOR2_X1 U458 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U459 ( .A(n405), .B(n404), .Z(n410) );
  XOR2_X1 U460 ( .A(KEYINPUT95), .B(KEYINPUT1), .Z(n407) );
  NAND2_X1 U461 ( .A1(G225GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U463 ( .A(KEYINPUT6), .B(n408), .ZN(n409) );
  XNOR2_X1 U464 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U465 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n412) );
  XNOR2_X1 U466 ( .A(KEYINPUT97), .B(KEYINPUT96), .ZN(n411) );
  XNOR2_X1 U467 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U468 ( .A(n414), .B(n413), .Z(n420) );
  XOR2_X1 U469 ( .A(KEYINPUT0), .B(G120GAT), .Z(n416) );
  XNOR2_X1 U470 ( .A(G113GAT), .B(G134GAT), .ZN(n415) );
  XNOR2_X1 U471 ( .A(n416), .B(n415), .ZN(n443) );
  XOR2_X1 U472 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n418) );
  XNOR2_X1 U473 ( .A(G141GAT), .B(KEYINPUT92), .ZN(n417) );
  XNOR2_X1 U474 ( .A(n418), .B(n417), .ZN(n423) );
  XNOR2_X1 U475 ( .A(n443), .B(n423), .ZN(n419) );
  XOR2_X1 U476 ( .A(n420), .B(n419), .Z(n469) );
  AND2_X1 U477 ( .A1(n421), .A2(n469), .ZN(n422) );
  XOR2_X1 U478 ( .A(KEYINPUT65), .B(n422), .Z(n566) );
  XNOR2_X1 U479 ( .A(n424), .B(n423), .ZN(n440) );
  XOR2_X1 U480 ( .A(KEYINPUT23), .B(G204GAT), .Z(n426) );
  XNOR2_X1 U481 ( .A(G218GAT), .B(G211GAT), .ZN(n425) );
  XNOR2_X1 U482 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U483 ( .A(n428), .B(n427), .Z(n430) );
  NAND2_X1 U484 ( .A1(G228GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U486 ( .A(KEYINPUT22), .B(KEYINPUT94), .Z(n432) );
  XNOR2_X1 U487 ( .A(KEYINPUT24), .B(KEYINPUT93), .ZN(n431) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U489 ( .A(n434), .B(n433), .Z(n438) );
  XOR2_X1 U490 ( .A(n436), .B(n435), .Z(n437) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n465) );
  NAND2_X1 U493 ( .A1(n566), .A2(n465), .ZN(n441) );
  XOR2_X1 U494 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U495 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U496 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U497 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n447) );
  XNOR2_X1 U498 ( .A(G183GAT), .B(G71GAT), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U500 ( .A(n449), .B(n448), .Z(n455) );
  XOR2_X1 U501 ( .A(G176GAT), .B(G99GAT), .Z(n451) );
  XNOR2_X1 U502 ( .A(G43GAT), .B(G190GAT), .ZN(n450) );
  XNOR2_X1 U503 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U504 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U505 ( .A(n455), .B(n454), .Z(n525) );
  INV_X1 U506 ( .A(n525), .ZN(n516) );
  NAND2_X1 U507 ( .A1(n456), .A2(n516), .ZN(n563) );
  NOR2_X1 U508 ( .A1(n535), .A2(n563), .ZN(n459) );
  INV_X1 U509 ( .A(KEYINPUT58), .ZN(n457) );
  NAND2_X1 U510 ( .A1(n572), .A2(n544), .ZN(n485) );
  NAND2_X1 U511 ( .A1(n550), .A2(n535), .ZN(n460) );
  XNOR2_X1 U512 ( .A(n460), .B(KEYINPUT89), .ZN(n461) );
  XNOR2_X1 U513 ( .A(n461), .B(KEYINPUT16), .ZN(n473) );
  XOR2_X1 U514 ( .A(n465), .B(KEYINPUT28), .Z(n518) );
  INV_X1 U515 ( .A(n469), .ZN(n511) );
  XNOR2_X1 U516 ( .A(n513), .B(KEYINPUT27), .ZN(n463) );
  NAND2_X1 U517 ( .A1(n511), .A2(n463), .ZN(n543) );
  NOR2_X1 U518 ( .A1(n518), .A2(n543), .ZN(n523) );
  NAND2_X1 U519 ( .A1(n523), .A2(n525), .ZN(n472) );
  NOR2_X1 U520 ( .A1(n465), .A2(n516), .ZN(n462) );
  XNOR2_X1 U521 ( .A(n462), .B(KEYINPUT26), .ZN(n565) );
  NAND2_X1 U522 ( .A1(n463), .A2(n565), .ZN(n468) );
  NAND2_X1 U523 ( .A1(n516), .A2(n513), .ZN(n464) );
  NAND2_X1 U524 ( .A1(n465), .A2(n464), .ZN(n466) );
  XOR2_X1 U525 ( .A(KEYINPUT25), .B(n466), .Z(n467) );
  NAND2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n470) );
  NAND2_X1 U527 ( .A1(n470), .A2(n469), .ZN(n471) );
  NAND2_X1 U528 ( .A1(n472), .A2(n471), .ZN(n481) );
  NAND2_X1 U529 ( .A1(n473), .A2(n481), .ZN(n500) );
  NOR2_X1 U530 ( .A1(n485), .A2(n500), .ZN(n479) );
  NAND2_X1 U531 ( .A1(n479), .A2(n511), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n474), .B(KEYINPUT34), .ZN(n475) );
  XNOR2_X1 U533 ( .A(G1GAT), .B(n475), .ZN(G1324GAT) );
  NAND2_X1 U534 ( .A1(n479), .A2(n513), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n476), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(G15GAT), .B(KEYINPUT35), .Z(n478) );
  NAND2_X1 U537 ( .A1(n479), .A2(n516), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  NAND2_X1 U539 ( .A1(n479), .A2(n518), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n480), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U541 ( .A(KEYINPUT39), .B(KEYINPUT101), .Z(n488) );
  INV_X1 U542 ( .A(n550), .ZN(n576) );
  NAND2_X1 U543 ( .A1(n576), .A2(n481), .ZN(n482) );
  XOR2_X1 U544 ( .A(KEYINPUT100), .B(n482), .Z(n483) );
  NAND2_X1 U545 ( .A1(n483), .A2(n581), .ZN(n484) );
  XOR2_X1 U546 ( .A(KEYINPUT37), .B(n484), .Z(n509) );
  NOR2_X1 U547 ( .A1(n485), .A2(n509), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n486), .B(KEYINPUT38), .ZN(n495) );
  NAND2_X1 U549 ( .A1(n511), .A2(n495), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U551 ( .A(G29GAT), .B(n489), .Z(G1328GAT) );
  NAND2_X1 U552 ( .A1(n495), .A2(n513), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n490), .B(KEYINPUT102), .ZN(n491) );
  XNOR2_X1 U554 ( .A(G36GAT), .B(n491), .ZN(G1329GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n493) );
  NAND2_X1 U556 ( .A1(n516), .A2(n495), .ZN(n492) );
  XNOR2_X1 U557 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U558 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT105), .B(KEYINPUT104), .Z(n497) );
  NAND2_X1 U560 ( .A1(n518), .A2(n495), .ZN(n496) );
  XNOR2_X1 U561 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U562 ( .A(G50GAT), .B(n498), .ZN(G1331GAT) );
  XNOR2_X1 U563 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n502) );
  NOR2_X1 U564 ( .A1(n544), .A2(n559), .ZN(n499) );
  XOR2_X1 U565 ( .A(KEYINPUT106), .B(n499), .Z(n510) );
  NOR2_X1 U566 ( .A1(n510), .A2(n500), .ZN(n505) );
  NAND2_X1 U567 ( .A1(n511), .A2(n505), .ZN(n501) );
  XNOR2_X1 U568 ( .A(n502), .B(n501), .ZN(G1332GAT) );
  NAND2_X1 U569 ( .A1(n505), .A2(n513), .ZN(n503) );
  XNOR2_X1 U570 ( .A(n503), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U571 ( .A1(n505), .A2(n516), .ZN(n504) );
  XNOR2_X1 U572 ( .A(n504), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n507) );
  NAND2_X1 U574 ( .A1(n505), .A2(n518), .ZN(n506) );
  XNOR2_X1 U575 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U576 ( .A(G78GAT), .B(n508), .Z(G1335GAT) );
  NOR2_X1 U577 ( .A1(n510), .A2(n509), .ZN(n519) );
  NAND2_X1 U578 ( .A1(n511), .A2(n519), .ZN(n512) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(n512), .ZN(G1336GAT) );
  NAND2_X1 U580 ( .A1(n519), .A2(n513), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n514), .B(KEYINPUT108), .ZN(n515) );
  XNOR2_X1 U582 ( .A(G92GAT), .B(n515), .ZN(G1337GAT) );
  NAND2_X1 U583 ( .A1(n519), .A2(n516), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n517), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT109), .B(KEYINPUT44), .Z(n521) );
  NAND2_X1 U586 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n522), .ZN(G1339GAT) );
  NAND2_X1 U589 ( .A1(n541), .A2(n523), .ZN(n524) );
  NOR2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n531) );
  NAND2_X1 U591 ( .A1(n544), .A2(n531), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n526), .B(KEYINPUT114), .ZN(n527) );
  XNOR2_X1 U593 ( .A(G113GAT), .B(n527), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n529) );
  INV_X1 U595 ( .A(n559), .ZN(n546) );
  NAND2_X1 U596 ( .A1(n531), .A2(n546), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U598 ( .A(G120GAT), .B(n530), .Z(G1341GAT) );
  INV_X1 U599 ( .A(n531), .ZN(n536) );
  NOR2_X1 U600 ( .A1(n562), .A2(n536), .ZN(n533) );
  XNOR2_X1 U601 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n532) );
  XNOR2_X1 U602 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U603 ( .A(G127GAT), .B(n534), .Z(G1342GAT) );
  NOR2_X1 U604 ( .A1(n536), .A2(n535), .ZN(n540) );
  XOR2_X1 U605 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n538) );
  XNOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT117), .ZN(n537) );
  XNOR2_X1 U607 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  NAND2_X1 U609 ( .A1(n541), .A2(n565), .ZN(n542) );
  NOR2_X1 U610 ( .A1(n543), .A2(n542), .ZN(n553) );
  NAND2_X1 U611 ( .A1(n544), .A2(n553), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n545), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n548) );
  NAND2_X1 U614 ( .A1(n553), .A2(n546), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(n549), .ZN(G1345GAT) );
  XOR2_X1 U617 ( .A(G155GAT), .B(KEYINPUT119), .Z(n552) );
  NAND2_X1 U618 ( .A1(n553), .A2(n550), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(G1346GAT) );
  NAND2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U622 ( .A1(n567), .A2(n563), .ZN(n556) );
  XOR2_X1 U623 ( .A(G169GAT), .B(n556), .Z(G1348GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n558) );
  XNOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(n561) );
  NOR2_X1 U627 ( .A1(n563), .A2(n559), .ZN(n560) );
  XOR2_X1 U628 ( .A(n561), .B(n560), .Z(G1349GAT) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U630 ( .A(G183GAT), .B(n564), .Z(G1350GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n580) );
  NOR2_X1 U632 ( .A1(n580), .A2(n567), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n580), .ZN(n574) );
  XNOR2_X1 U638 ( .A(KEYINPUT61), .B(KEYINPUT124), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(n575), .ZN(G1353GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n580), .ZN(n578) );
  XNOR2_X1 U642 ( .A(KEYINPUT125), .B(KEYINPUT126), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(n579), .ZN(G1354GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n584) );
  INV_X1 U646 ( .A(n580), .ZN(n582) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

