

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760;

  XNOR2_X1 U377 ( .A(n693), .B(n370), .ZN(n602) );
  AND2_X1 U378 ( .A1(n624), .A2(n623), .ZN(n747) );
  INV_X2 U379 ( .A(G953), .ZN(n748) );
  NOR2_X2 U380 ( .A1(n759), .A2(n563), .ZN(n450) );
  NOR2_X2 U381 ( .A1(n688), .A2(n550), .ZN(n547) );
  XNOR2_X2 U382 ( .A(n412), .B(n545), .ZN(n688) );
  NAND2_X1 U383 ( .A1(n757), .A2(n758), .ZN(n388) );
  NOR2_X2 U384 ( .A1(n550), .A2(n359), .ZN(n429) );
  NOR2_X2 U385 ( .A1(n583), .A2(n577), .ZN(n578) );
  INV_X1 U386 ( .A(n418), .ZN(n696) );
  XNOR2_X1 U387 ( .A(n518), .B(n517), .ZN(n746) );
  XNOR2_X1 U388 ( .A(n388), .B(n458), .ZN(n387) );
  XNOR2_X1 U389 ( .A(n582), .B(KEYINPUT40), .ZN(n757) );
  NAND2_X1 U390 ( .A1(n621), .A2(n655), .ZN(n582) );
  XNOR2_X1 U391 ( .A(n456), .B(n363), .ZN(n621) );
  XNOR2_X2 U392 ( .A(n423), .B(n477), .ZN(n379) );
  OR2_X1 U393 ( .A1(n730), .A2(G902), .ZN(n460) );
  NAND2_X1 U394 ( .A1(n453), .A2(n486), .ZN(n518) );
  INV_X1 U395 ( .A(KEYINPUT0), .ZN(n420) );
  NAND2_X1 U396 ( .A1(n360), .A2(n387), .ZN(n386) );
  AND2_X1 U397 ( .A1(n579), .A2(n580), .ZN(n592) );
  BUF_X1 U398 ( .A(n695), .Z(n385) );
  XNOR2_X1 U399 ( .A(n417), .B(n413), .ZN(n537) );
  XNOR2_X1 U400 ( .A(n415), .B(n414), .ZN(n413) );
  XNOR2_X1 U401 ( .A(n416), .B(G128), .ZN(n415) );
  INV_X1 U402 ( .A(KEYINPUT23), .ZN(n416) );
  XNOR2_X1 U403 ( .A(KEYINPUT96), .B(KEYINPUT95), .ZN(n414) );
  AND2_X1 U404 ( .A1(n399), .A2(n423), .ZN(n398) );
  OR2_X1 U405 ( .A1(n602), .A2(n402), .ZN(n399) );
  XNOR2_X1 U406 ( .A(n586), .B(n524), .ZN(n695) );
  XNOR2_X1 U407 ( .A(n358), .B(n465), .ZN(n525) );
  XNOR2_X1 U408 ( .A(G119), .B(KEYINPUT3), .ZN(n465) );
  XNOR2_X1 U409 ( .A(n443), .B(G140), .ZN(n538) );
  INV_X1 U410 ( .A(G137), .ZN(n443) );
  OR2_X1 U411 ( .A1(n725), .A2(G902), .ZN(n454) );
  INV_X1 U412 ( .A(KEYINPUT6), .ZN(n370) );
  XNOR2_X1 U413 ( .A(n746), .B(n519), .ZN(n409) );
  OR2_X1 U414 ( .A1(n602), .A2(n378), .ZN(n377) );
  NAND2_X1 U415 ( .A1(n695), .A2(n690), .ZN(n378) );
  XNOR2_X1 U416 ( .A(n429), .B(KEYINPUT22), .ZN(n422) );
  OR2_X1 U417 ( .A1(n756), .A2(n649), .ZN(n375) );
  XNOR2_X1 U418 ( .A(G122), .B(G140), .ZN(n504) );
  XNOR2_X1 U419 ( .A(n406), .B(G146), .ZN(n497) );
  INV_X1 U420 ( .A(G125), .ZN(n406) );
  INV_X1 U421 ( .A(G134), .ZN(n485) );
  NAND2_X1 U422 ( .A1(n418), .A2(KEYINPUT110), .ZN(n436) );
  AND2_X1 U423 ( .A1(n410), .A2(n437), .ZN(n384) );
  NAND2_X1 U424 ( .A1(n444), .A2(n401), .ZN(n400) );
  AND2_X1 U425 ( .A1(n602), .A2(n402), .ZN(n401) );
  INV_X1 U426 ( .A(KEYINPUT112), .ZN(n402) );
  XNOR2_X1 U427 ( .A(n604), .B(KEYINPUT89), .ZN(n605) );
  AND2_X1 U428 ( .A1(n655), .A2(n445), .ZN(n444) );
  INV_X1 U429 ( .A(n603), .ZN(n445) );
  INV_X1 U430 ( .A(KEYINPUT90), .ZN(n451) );
  XNOR2_X1 U431 ( .A(n508), .B(n507), .ZN(n557) );
  XNOR2_X1 U432 ( .A(KEYINPUT13), .B(G475), .ZN(n507) );
  XNOR2_X1 U433 ( .A(n409), .B(n446), .ZN(n637) );
  XNOR2_X1 U434 ( .A(n529), .B(n447), .ZN(n446) );
  INV_X1 U435 ( .A(n525), .ZN(n447) );
  XNOR2_X1 U436 ( .A(n386), .B(n457), .ZN(n624) );
  XNOR2_X1 U437 ( .A(n424), .B(n525), .ZN(n733) );
  XNOR2_X1 U438 ( .A(n421), .B(n461), .ZN(n424) );
  XNOR2_X1 U439 ( .A(n382), .B(KEYINPUT16), .ZN(n461) );
  XNOR2_X1 U440 ( .A(KEYINPUT67), .B(G122), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n407), .B(n403), .ZN(n726) );
  XNOR2_X1 U442 ( .A(n539), .B(n404), .ZN(n403) );
  XNOR2_X1 U443 ( .A(n506), .B(n408), .ZN(n407) );
  XNOR2_X1 U444 ( .A(n498), .B(n501), .ZN(n404) );
  NOR2_X1 U445 ( .A1(n385), .A2(n602), .ZN(n380) );
  XNOR2_X1 U446 ( .A(n542), .B(n543), .ZN(n459) );
  XNOR2_X1 U447 ( .A(n442), .B(n441), .ZN(n523) );
  XNOR2_X1 U448 ( .A(n521), .B(KEYINPUT75), .ZN(n441) );
  XNOR2_X1 U449 ( .A(KEYINPUT46), .B(KEYINPUT85), .ZN(n458) );
  NOR2_X1 U450 ( .A1(n418), .A2(KEYINPUT110), .ZN(n438) );
  INV_X1 U451 ( .A(KEYINPUT48), .ZN(n457) );
  XNOR2_X1 U452 ( .A(n505), .B(n502), .ZN(n408) );
  XNOR2_X1 U453 ( .A(G113), .B(G104), .ZN(n499) );
  XNOR2_X1 U454 ( .A(n497), .B(n405), .ZN(n539) );
  INV_X1 U455 ( .A(KEYINPUT10), .ZN(n405) );
  XNOR2_X1 U456 ( .A(n516), .B(n515), .ZN(n517) );
  INV_X1 U457 ( .A(KEYINPUT4), .ZN(n515) );
  XNOR2_X1 U458 ( .A(G131), .B(KEYINPUT66), .ZN(n516) );
  XNOR2_X1 U459 ( .A(n533), .B(n534), .ZN(n417) );
  XNOR2_X1 U460 ( .A(G116), .B(G107), .ZN(n487) );
  XOR2_X1 U461 ( .A(KEYINPUT9), .B(G122), .Z(n488) );
  NOR2_X1 U462 ( .A1(KEYINPUT69), .A2(n626), .ZN(n625) );
  XOR2_X1 U463 ( .A(G902), .B(KEYINPUT15), .Z(n628) );
  INV_X1 U464 ( .A(KEYINPUT74), .ZN(n520) );
  XNOR2_X1 U465 ( .A(n522), .B(n538), .ZN(n442) );
  XNOR2_X1 U466 ( .A(n470), .B(n471), .ZN(n426) );
  INV_X1 U467 ( .A(KEYINPUT33), .ZN(n545) );
  NOR2_X1 U468 ( .A1(n673), .A2(n672), .ZN(n674) );
  INV_X1 U469 ( .A(n591), .ZN(n619) );
  NAND2_X1 U470 ( .A1(n444), .A2(n602), .ZN(n616) );
  NAND2_X1 U471 ( .A1(n398), .A2(n396), .ZN(n395) );
  INV_X1 U472 ( .A(n400), .ZN(n394) );
  OR2_X1 U473 ( .A1(n444), .A2(n402), .ZN(n397) );
  OR2_X1 U474 ( .A1(n444), .A2(n364), .ZN(n389) );
  NAND2_X1 U475 ( .A1(n392), .A2(n605), .ZN(n391) );
  XNOR2_X1 U476 ( .A(n440), .B(n367), .ZN(n372) );
  NOR2_X1 U477 ( .A1(n553), .A2(n371), .ZN(n701) );
  NOR2_X1 U478 ( .A1(n371), .A2(n603), .ZN(n585) );
  XNOR2_X1 U479 ( .A(n557), .B(KEYINPUT106), .ZN(n559) );
  XNOR2_X1 U480 ( .A(n637), .B(n636), .ZN(n638) );
  INV_X1 U481 ( .A(KEYINPUT79), .ZN(n376) );
  AND2_X1 U482 ( .A1(n559), .A2(n558), .ZN(n655) );
  AND2_X1 U483 ( .A1(n422), .A2(n368), .ZN(n649) );
  NOR2_X1 U484 ( .A1(n385), .A2(n369), .ZN(n368) );
  NAND2_X1 U485 ( .A1(n371), .A2(n690), .ZN(n369) );
  NAND2_X1 U486 ( .A1(n554), .A2(n371), .ZN(n551) );
  XNOR2_X1 U487 ( .A(n434), .B(KEYINPUT109), .ZN(n759) );
  XNOR2_X1 U488 ( .A(n381), .B(KEYINPUT87), .ZN(n544) );
  INV_X1 U489 ( .A(KEYINPUT60), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n725), .B(n724), .ZN(n463) );
  XOR2_X1 U491 ( .A(KEYINPUT100), .B(G472), .Z(n357) );
  XOR2_X1 U492 ( .A(G113), .B(G116), .Z(n358) );
  NAND2_X1 U493 ( .A1(n588), .A2(n513), .ZN(n359) );
  AND2_X1 U494 ( .A1(n614), .A2(n615), .ZN(n360) );
  AND2_X1 U495 ( .A1(n391), .A2(n389), .ZN(n361) );
  INV_X1 U496 ( .A(n690), .ZN(n564) );
  OR2_X2 U497 ( .A1(n690), .A2(n689), .ZN(n418) );
  XOR2_X1 U498 ( .A(n377), .B(n376), .Z(n362) );
  XOR2_X1 U499 ( .A(n581), .B(KEYINPUT39), .Z(n363) );
  INV_X1 U500 ( .A(KEYINPUT110), .ZN(n452) );
  OR2_X1 U501 ( .A1(n396), .A2(n402), .ZN(n364) );
  XOR2_X1 U502 ( .A(n721), .B(n720), .Z(n365) );
  XNOR2_X1 U503 ( .A(n726), .B(KEYINPUT59), .ZN(n366) );
  XNOR2_X1 U504 ( .A(KEYINPUT76), .B(KEYINPUT35), .ZN(n367) );
  NOR2_X1 U505 ( .A1(G952), .A2(n748), .ZN(n732) );
  INV_X1 U506 ( .A(n732), .ZN(n432) );
  AND2_X1 U507 ( .A1(n436), .A2(n602), .ZN(n411) );
  INV_X1 U508 ( .A(n693), .ZN(n371) );
  XNOR2_X2 U509 ( .A(n530), .B(n357), .ZN(n693) );
  INV_X1 U510 ( .A(n372), .ZN(n373) );
  NAND2_X1 U511 ( .A1(n372), .A2(KEYINPUT44), .ZN(n439) );
  NAND2_X1 U512 ( .A1(n374), .A2(n372), .ZN(n566) );
  XNOR2_X1 U513 ( .A(n373), .B(G122), .ZN(G24) );
  INV_X1 U514 ( .A(n375), .ZN(n374) );
  XNOR2_X1 U515 ( .A(n375), .B(KEYINPUT44), .ZN(n567) );
  NOR2_X2 U516 ( .A1(n379), .A2(n482), .ZN(n419) );
  NOR2_X1 U517 ( .A1(n595), .A2(n379), .ZN(n656) );
  NAND2_X1 U518 ( .A1(n422), .A2(n380), .ZN(n381) );
  XNOR2_X1 U519 ( .A(n383), .B(n428), .ZN(n427) );
  XNOR2_X1 U520 ( .A(n497), .B(n514), .ZN(n383) );
  INV_X2 U521 ( .A(n466), .ZN(n468) );
  XNOR2_X2 U522 ( .A(n468), .B(n467), .ZN(n421) );
  NAND2_X1 U523 ( .A1(n384), .A2(n411), .ZN(n412) );
  XNOR2_X1 U524 ( .A(n427), .B(n426), .ZN(n425) );
  XNOR2_X1 U525 ( .A(n733), .B(n425), .ZN(n719) );
  NAND2_X1 U526 ( .A1(n390), .A2(n361), .ZN(n606) );
  NAND2_X1 U527 ( .A1(n393), .A2(n397), .ZN(n390) );
  NAND2_X1 U528 ( .A1(n400), .A2(n398), .ZN(n392) );
  NOR2_X1 U529 ( .A1(n395), .A2(n394), .ZN(n393) );
  INV_X1 U530 ( .A(n605), .ZN(n396) );
  XNOR2_X1 U531 ( .A(n409), .B(n455), .ZN(n725) );
  OR2_X1 U532 ( .A1(n695), .A2(n452), .ZN(n410) );
  XNOR2_X2 U533 ( .A(n460), .B(n459), .ZN(n690) );
  XNOR2_X2 U534 ( .A(n419), .B(n420), .ZN(n550) );
  XNOR2_X2 U535 ( .A(n475), .B(n451), .ZN(n423) );
  XNOR2_X1 U536 ( .A(n421), .B(n523), .ZN(n455) );
  AND2_X1 U537 ( .A1(n422), .A2(n362), .ZN(n565) );
  XNOR2_X1 U538 ( .A(n484), .B(n469), .ZN(n428) );
  XNOR2_X1 U539 ( .A(n722), .B(n365), .ZN(n723) );
  NAND2_X1 U540 ( .A1(n728), .A2(G210), .ZN(n722) );
  XNOR2_X1 U541 ( .A(n431), .B(n430), .ZN(G60) );
  NAND2_X1 U542 ( .A1(n433), .A2(n432), .ZN(n431) );
  XNOR2_X1 U543 ( .A(n727), .B(n366), .ZN(n433) );
  NAND2_X1 U544 ( .A1(n544), .A2(n564), .ZN(n434) );
  XNOR2_X1 U545 ( .A(n448), .B(KEYINPUT45), .ZN(n670) );
  XNOR2_X2 U546 ( .A(n675), .B(n625), .ZN(n630) );
  XNOR2_X2 U547 ( .A(G110), .B(KEYINPUT68), .ZN(n467) );
  NOR2_X2 U548 ( .A1(n640), .A2(n732), .ZN(n642) );
  XNOR2_X1 U549 ( .A(n435), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U550 ( .A1(n723), .A2(n732), .ZN(n435) );
  NAND2_X1 U551 ( .A1(n385), .A2(n696), .ZN(n553) );
  NAND2_X1 U552 ( .A1(n695), .A2(n438), .ZN(n437) );
  NAND2_X1 U553 ( .A1(n439), .A2(n562), .ZN(n563) );
  NAND2_X1 U554 ( .A1(n549), .A2(n548), .ZN(n440) );
  INV_X1 U555 ( .A(n483), .ZN(n484) );
  XNOR2_X2 U556 ( .A(G128), .B(G143), .ZN(n483) );
  NAND2_X1 U557 ( .A1(n484), .A2(n485), .ZN(n453) );
  NAND2_X1 U558 ( .A1(n449), .A2(n568), .ZN(n448) );
  XNOR2_X1 U559 ( .A(n450), .B(KEYINPUT88), .ZN(n449) );
  XNOR2_X2 U560 ( .A(n454), .B(G469), .ZN(n586) );
  NAND2_X1 U561 ( .A1(n592), .A2(n680), .ZN(n456) );
  NOR2_X1 U562 ( .A1(n462), .A2(n732), .ZN(G54) );
  XNOR2_X1 U563 ( .A(n464), .B(n463), .ZN(n462) );
  NAND2_X1 U564 ( .A1(n728), .A2(G469), .ZN(n464) );
  XNOR2_X1 U565 ( .A(n473), .B(n472), .ZN(n569) );
  NOR2_X1 U566 ( .A1(n719), .A2(n628), .ZN(n473) );
  INV_X1 U567 ( .A(KEYINPUT104), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(n505) );
  INV_X1 U569 ( .A(n667), .ZN(n622) );
  INV_X1 U570 ( .A(n689), .ZN(n513) );
  AND2_X1 U571 ( .A1(n669), .A2(n622), .ZN(n623) );
  XNOR2_X1 U572 ( .A(n520), .B(KEYINPUT94), .ZN(n521) );
  INV_X1 U573 ( .A(KEYINPUT86), .ZN(n581) );
  XNOR2_X1 U574 ( .A(n476), .B(KEYINPUT19), .ZN(n477) );
  XNOR2_X1 U575 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X2 U576 ( .A(G104), .B(G107), .ZN(n466) );
  XOR2_X2 U577 ( .A(G101), .B(KEYINPUT65), .Z(n514) );
  XOR2_X1 U578 ( .A(KEYINPUT4), .B(KEYINPUT17), .Z(n470) );
  XNOR2_X1 U579 ( .A(KEYINPUT92), .B(KEYINPUT18), .ZN(n469) );
  NAND2_X1 U580 ( .A1(G224), .A2(n748), .ZN(n471) );
  OR2_X1 U581 ( .A1(G902), .A2(G237), .ZN(n474) );
  NAND2_X1 U582 ( .A1(G210), .A2(n474), .ZN(n472) );
  NAND2_X1 U583 ( .A1(G214), .A2(n474), .ZN(n679) );
  NAND2_X1 U584 ( .A1(n569), .A2(n679), .ZN(n475) );
  INV_X1 U585 ( .A(KEYINPUT71), .ZN(n476) );
  NOR2_X1 U586 ( .A1(G898), .A2(n748), .ZN(n478) );
  XOR2_X1 U587 ( .A(KEYINPUT93), .B(n478), .Z(n735) );
  NAND2_X1 U588 ( .A1(n735), .A2(G902), .ZN(n479) );
  NAND2_X1 U589 ( .A1(G952), .A2(n748), .ZN(n574) );
  NAND2_X1 U590 ( .A1(n479), .A2(n574), .ZN(n481) );
  NAND2_X1 U591 ( .A1(G234), .A2(G237), .ZN(n480) );
  XOR2_X1 U592 ( .A(KEYINPUT14), .B(n480), .Z(n710) );
  INV_X1 U593 ( .A(n710), .ZN(n576) );
  NAND2_X1 U594 ( .A1(n481), .A2(n576), .ZN(n482) );
  NAND2_X1 U595 ( .A1(G134), .A2(n483), .ZN(n486) );
  XNOR2_X1 U596 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U597 ( .A(n518), .B(n489), .Z(n492) );
  NAND2_X1 U598 ( .A1(G234), .A2(n748), .ZN(n490) );
  XOR2_X1 U599 ( .A(KEYINPUT8), .B(n490), .Z(n535) );
  NAND2_X1 U600 ( .A1(G217), .A2(n535), .ZN(n491) );
  XNOR2_X1 U601 ( .A(n492), .B(n491), .ZN(n494) );
  XOR2_X1 U602 ( .A(KEYINPUT107), .B(KEYINPUT7), .Z(n493) );
  XNOR2_X1 U603 ( .A(n494), .B(n493), .ZN(n631) );
  NOR2_X1 U604 ( .A1(G902), .A2(n631), .ZN(n496) );
  XNOR2_X1 U605 ( .A(KEYINPUT108), .B(G478), .ZN(n495) );
  XNOR2_X1 U606 ( .A(n496), .B(n495), .ZN(n558) );
  INV_X1 U607 ( .A(n558), .ZN(n560) );
  NOR2_X1 U608 ( .A1(G953), .A2(G237), .ZN(n526) );
  NAND2_X1 U609 ( .A1(n526), .A2(G214), .ZN(n498) );
  XOR2_X1 U610 ( .A(KEYINPUT11), .B(G143), .Z(n500) );
  XNOR2_X1 U611 ( .A(n500), .B(n499), .ZN(n506) );
  XOR2_X1 U612 ( .A(KEYINPUT12), .B(KEYINPUT103), .Z(n502) );
  XNOR2_X1 U613 ( .A(G131), .B(KEYINPUT105), .ZN(n501) );
  NOR2_X1 U614 ( .A1(G902), .A2(n726), .ZN(n508) );
  NOR2_X1 U615 ( .A1(n560), .A2(n557), .ZN(n588) );
  INV_X1 U616 ( .A(n628), .ZN(n509) );
  NAND2_X1 U617 ( .A1(G234), .A2(n509), .ZN(n510) );
  XNOR2_X1 U618 ( .A(KEYINPUT20), .B(n510), .ZN(n541) );
  NAND2_X1 U619 ( .A1(n541), .A2(G221), .ZN(n511) );
  XNOR2_X1 U620 ( .A(n511), .B(KEYINPUT21), .ZN(n512) );
  XOR2_X1 U621 ( .A(KEYINPUT99), .B(n512), .Z(n689) );
  XNOR2_X1 U622 ( .A(G146), .B(n514), .ZN(n519) );
  NAND2_X1 U623 ( .A1(G227), .A2(n748), .ZN(n522) );
  XNOR2_X1 U624 ( .A(KEYINPUT64), .B(KEYINPUT1), .ZN(n524) );
  XOR2_X1 U625 ( .A(G137), .B(KEYINPUT5), .Z(n528) );
  NAND2_X1 U626 ( .A1(n526), .A2(G210), .ZN(n527) );
  XNOR2_X1 U627 ( .A(n528), .B(n527), .ZN(n529) );
  NOR2_X1 U628 ( .A1(G902), .A2(n637), .ZN(n530) );
  XOR2_X1 U629 ( .A(KEYINPUT72), .B(KEYINPUT98), .Z(n532) );
  XNOR2_X1 U630 ( .A(KEYINPUT25), .B(KEYINPUT97), .ZN(n531) );
  XNOR2_X1 U631 ( .A(n532), .B(n531), .ZN(n543) );
  XNOR2_X1 U632 ( .A(G119), .B(G110), .ZN(n533) );
  XNOR2_X1 U633 ( .A(KEYINPUT24), .B(KEYINPUT73), .ZN(n534) );
  NAND2_X1 U634 ( .A1(G221), .A2(n535), .ZN(n536) );
  XNOR2_X1 U635 ( .A(n537), .B(n536), .ZN(n540) );
  XNOR2_X1 U636 ( .A(n539), .B(n538), .ZN(n745) );
  XNOR2_X1 U637 ( .A(n540), .B(n745), .ZN(n730) );
  NAND2_X1 U638 ( .A1(G217), .A2(n541), .ZN(n542) );
  XNOR2_X1 U639 ( .A(KEYINPUT34), .B(KEYINPUT78), .ZN(n546) );
  XNOR2_X1 U640 ( .A(n547), .B(n546), .ZN(n549) );
  NAND2_X1 U641 ( .A1(n557), .A2(n560), .ZN(n594) );
  XNOR2_X1 U642 ( .A(n594), .B(KEYINPUT77), .ZN(n548) );
  INV_X1 U643 ( .A(n550), .ZN(n554) );
  NAND2_X1 U644 ( .A1(n586), .A2(n696), .ZN(n577) );
  NOR2_X1 U645 ( .A1(n551), .A2(n577), .ZN(n552) );
  XNOR2_X1 U646 ( .A(n552), .B(KEYINPUT101), .ZN(n644) );
  AND2_X1 U647 ( .A1(n554), .A2(n701), .ZN(n556) );
  XNOR2_X1 U648 ( .A(KEYINPUT102), .B(KEYINPUT31), .ZN(n555) );
  XNOR2_X1 U649 ( .A(n556), .B(n555), .ZN(n661) );
  NAND2_X1 U650 ( .A1(n644), .A2(n661), .ZN(n561) );
  NOR2_X1 U651 ( .A1(n558), .A2(n559), .ZN(n651) );
  NOR2_X1 U652 ( .A1(n651), .A2(n655), .ZN(n684) );
  INV_X1 U653 ( .A(n684), .ZN(n598) );
  NAND2_X1 U654 ( .A1(n561), .A2(n598), .ZN(n562) );
  XNOR2_X1 U655 ( .A(KEYINPUT32), .B(n565), .ZN(n756) );
  NAND2_X1 U656 ( .A1(n567), .A2(n566), .ZN(n568) );
  BUF_X1 U657 ( .A(n569), .Z(n591) );
  XNOR2_X1 U658 ( .A(KEYINPUT38), .B(n619), .ZN(n680) );
  NAND2_X1 U659 ( .A1(n693), .A2(n679), .ZN(n570) );
  XNOR2_X1 U660 ( .A(n570), .B(KEYINPUT111), .ZN(n571) );
  XNOR2_X1 U661 ( .A(KEYINPUT30), .B(n571), .ZN(n580) );
  NOR2_X1 U662 ( .A1(G900), .A2(n748), .ZN(n572) );
  NAND2_X1 U663 ( .A1(G902), .A2(n572), .ZN(n573) );
  NAND2_X1 U664 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U665 ( .A1(n576), .A2(n575), .ZN(n583) );
  XNOR2_X1 U666 ( .A(KEYINPUT70), .B(n578), .ZN(n579) );
  NOR2_X1 U667 ( .A1(n689), .A2(n583), .ZN(n584) );
  NAND2_X1 U668 ( .A1(n690), .A2(n584), .ZN(n603) );
  XNOR2_X1 U669 ( .A(KEYINPUT28), .B(n585), .ZN(n587) );
  NAND2_X1 U670 ( .A1(n587), .A2(n586), .ZN(n595) );
  INV_X1 U671 ( .A(n588), .ZN(n682) );
  NAND2_X1 U672 ( .A1(n680), .A2(n679), .ZN(n683) );
  NOR2_X1 U673 ( .A1(n682), .A2(n683), .ZN(n589) );
  XNOR2_X1 U674 ( .A(KEYINPUT41), .B(n589), .ZN(n704) );
  OR2_X1 U675 ( .A1(n595), .A2(n704), .ZN(n590) );
  XNOR2_X1 U676 ( .A(n590), .B(KEYINPUT42), .ZN(n758) );
  NAND2_X1 U677 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U678 ( .A1(n594), .A2(n593), .ZN(n654) );
  XNOR2_X1 U679 ( .A(KEYINPUT83), .B(n654), .ZN(n601) );
  INV_X1 U680 ( .A(KEYINPUT47), .ZN(n596) );
  NAND2_X1 U681 ( .A1(n596), .A2(n656), .ZN(n597) );
  NAND2_X1 U682 ( .A1(n597), .A2(KEYINPUT82), .ZN(n599) );
  NAND2_X1 U683 ( .A1(n599), .A2(n598), .ZN(n600) );
  AND2_X1 U684 ( .A1(n601), .A2(n600), .ZN(n615) );
  INV_X1 U685 ( .A(n385), .ZN(n607) );
  INV_X1 U686 ( .A(KEYINPUT36), .ZN(n604) );
  NOR2_X1 U687 ( .A1(n607), .A2(n606), .ZN(n665) );
  INV_X1 U688 ( .A(n665), .ZN(n613) );
  NAND2_X1 U689 ( .A1(KEYINPUT82), .A2(n684), .ZN(n608) );
  NAND2_X1 U690 ( .A1(n608), .A2(n656), .ZN(n609) );
  AND2_X1 U691 ( .A1(n609), .A2(KEYINPUT47), .ZN(n611) );
  NOR2_X1 U692 ( .A1(KEYINPUT82), .A2(KEYINPUT47), .ZN(n610) );
  NOR2_X1 U693 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U694 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U695 ( .A1(n385), .A2(n616), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n617), .A2(n679), .ZN(n618) );
  XNOR2_X1 U697 ( .A(n618), .B(KEYINPUT43), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n620), .A2(n619), .ZN(n669) );
  AND2_X1 U699 ( .A1(n621), .A2(n651), .ZN(n667) );
  AND2_X2 U700 ( .A1(n670), .A2(n747), .ZN(n675) );
  INV_X1 U701 ( .A(KEYINPUT2), .ZN(n626) );
  NAND2_X1 U702 ( .A1(KEYINPUT69), .A2(n626), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X4 U704 ( .A1(n630), .A2(n629), .ZN(n728) );
  NAND2_X1 U705 ( .A1(G478), .A2(n728), .ZN(n633) );
  INV_X1 U706 ( .A(n631), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n634), .A2(n432), .ZN(n635) );
  XNOR2_X1 U708 ( .A(n635), .B(KEYINPUT123), .ZN(G63) );
  NAND2_X1 U709 ( .A1(n728), .A2(G472), .ZN(n639) );
  XOR2_X1 U710 ( .A(KEYINPUT62), .B(KEYINPUT91), .Z(n636) );
  XNOR2_X1 U711 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U712 ( .A(KEYINPUT63), .B(KEYINPUT113), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n642), .B(n641), .ZN(G57) );
  INV_X1 U714 ( .A(n655), .ZN(n658) );
  NOR2_X1 U715 ( .A1(n658), .A2(n644), .ZN(n643) );
  XOR2_X1 U716 ( .A(G104), .B(n643), .Z(G6) );
  INV_X1 U717 ( .A(n651), .ZN(n660) );
  NOR2_X1 U718 ( .A1(n644), .A2(n660), .ZN(n648) );
  XOR2_X1 U719 ( .A(KEYINPUT26), .B(KEYINPUT115), .Z(n646) );
  XNOR2_X1 U720 ( .A(G107), .B(KEYINPUT27), .ZN(n645) );
  XNOR2_X1 U721 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U722 ( .A(n648), .B(n647), .ZN(G9) );
  XOR2_X1 U723 ( .A(G110), .B(n649), .Z(n650) );
  XNOR2_X1 U724 ( .A(KEYINPUT116), .B(n650), .ZN(G12) );
  XOR2_X1 U725 ( .A(G128), .B(KEYINPUT29), .Z(n653) );
  NAND2_X1 U726 ( .A1(n656), .A2(n651), .ZN(n652) );
  XNOR2_X1 U727 ( .A(n653), .B(n652), .ZN(G30) );
  XOR2_X1 U728 ( .A(G143), .B(n654), .Z(G45) );
  NAND2_X1 U729 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U730 ( .A(n657), .B(G146), .ZN(G48) );
  NOR2_X1 U731 ( .A1(n661), .A2(n658), .ZN(n659) );
  XOR2_X1 U732 ( .A(G113), .B(n659), .Z(G15) );
  NOR2_X1 U733 ( .A1(n661), .A2(n660), .ZN(n663) );
  XNOR2_X1 U734 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n662) );
  XNOR2_X1 U735 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U736 ( .A(G116), .B(n664), .ZN(G18) );
  XNOR2_X1 U737 ( .A(G125), .B(n665), .ZN(n666) );
  XNOR2_X1 U738 ( .A(n666), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U739 ( .A(G134), .B(n667), .ZN(n668) );
  XNOR2_X1 U740 ( .A(n668), .B(KEYINPUT119), .ZN(G36) );
  XNOR2_X1 U741 ( .A(G140), .B(n669), .ZN(G42) );
  BUF_X1 U742 ( .A(n670), .Z(n740) );
  NOR2_X1 U743 ( .A1(KEYINPUT2), .A2(n740), .ZN(n671) );
  XNOR2_X1 U744 ( .A(n671), .B(KEYINPUT84), .ZN(n673) );
  NOR2_X1 U745 ( .A1(KEYINPUT2), .A2(n747), .ZN(n672) );
  XNOR2_X1 U746 ( .A(n674), .B(KEYINPUT80), .ZN(n678) );
  NAND2_X1 U747 ( .A1(n675), .A2(KEYINPUT2), .ZN(n676) );
  XOR2_X1 U748 ( .A(KEYINPUT69), .B(n676), .Z(n677) );
  NAND2_X1 U749 ( .A1(n678), .A2(n677), .ZN(n716) );
  OR2_X1 U750 ( .A1(n688), .A2(n704), .ZN(n713) );
  NOR2_X1 U751 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U752 ( .A1(n682), .A2(n681), .ZN(n686) );
  NOR2_X1 U753 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U754 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U755 ( .A1(n688), .A2(n687), .ZN(n706) );
  AND2_X1 U756 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U757 ( .A(KEYINPUT49), .B(n691), .Z(n692) );
  NOR2_X1 U758 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U759 ( .A(KEYINPUT120), .B(n694), .Z(n699) );
  NOR2_X1 U760 ( .A1(n696), .A2(n385), .ZN(n697) );
  XNOR2_X1 U761 ( .A(KEYINPUT50), .B(n697), .ZN(n698) );
  NOR2_X1 U762 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U763 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U764 ( .A(KEYINPUT51), .B(n702), .Z(n703) );
  NOR2_X1 U765 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U766 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U767 ( .A(KEYINPUT121), .B(n707), .Z(n708) );
  XNOR2_X1 U768 ( .A(n708), .B(KEYINPUT52), .ZN(n709) );
  NOR2_X1 U769 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U770 ( .A1(n711), .A2(G952), .ZN(n712) );
  NAND2_X1 U771 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U772 ( .A1(G953), .A2(n714), .ZN(n715) );
  NAND2_X1 U773 ( .A1(n716), .A2(n715), .ZN(n718) );
  XOR2_X1 U774 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n717) );
  XNOR2_X1 U775 ( .A(n718), .B(n717), .ZN(G75) );
  XOR2_X1 U776 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n721) );
  XNOR2_X1 U777 ( .A(n719), .B(KEYINPUT81), .ZN(n720) );
  XOR2_X1 U778 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n724) );
  NAND2_X1 U779 ( .A1(n728), .A2(G475), .ZN(n727) );
  NAND2_X1 U780 ( .A1(G217), .A2(n728), .ZN(n729) );
  XNOR2_X1 U781 ( .A(n730), .B(n729), .ZN(n731) );
  NOR2_X1 U782 ( .A1(n732), .A2(n731), .ZN(G66) );
  XOR2_X1 U783 ( .A(n733), .B(G101), .Z(n734) );
  NOR2_X1 U784 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U785 ( .A(KEYINPUT125), .B(n736), .Z(n744) );
  NAND2_X1 U786 ( .A1(G224), .A2(G953), .ZN(n737) );
  XNOR2_X1 U787 ( .A(n737), .B(KEYINPUT61), .ZN(n738) );
  XNOR2_X1 U788 ( .A(KEYINPUT124), .B(n738), .ZN(n739) );
  NAND2_X1 U789 ( .A1(G898), .A2(n739), .ZN(n742) );
  NAND2_X1 U790 ( .A1(n740), .A2(n748), .ZN(n741) );
  NAND2_X1 U791 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U792 ( .A(n744), .B(n743), .ZN(G69) );
  XOR2_X1 U793 ( .A(n746), .B(n745), .Z(n750) );
  XOR2_X1 U794 ( .A(n747), .B(n750), .Z(n749) );
  NAND2_X1 U795 ( .A1(n749), .A2(n748), .ZN(n754) );
  XNOR2_X1 U796 ( .A(G227), .B(n750), .ZN(n751) );
  NAND2_X1 U797 ( .A1(n751), .A2(G900), .ZN(n752) );
  NAND2_X1 U798 ( .A1(G953), .A2(n752), .ZN(n753) );
  NAND2_X1 U799 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U800 ( .A(KEYINPUT126), .B(n755), .ZN(G72) );
  XOR2_X1 U801 ( .A(G119), .B(n756), .Z(G21) );
  XNOR2_X1 U802 ( .A(G131), .B(n757), .ZN(G33) );
  XNOR2_X1 U803 ( .A(G137), .B(n758), .ZN(G39) );
  XOR2_X1 U804 ( .A(n759), .B(G101), .Z(n760) );
  XNOR2_X1 U805 ( .A(KEYINPUT114), .B(n760), .ZN(G3) );
endmodule

