//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995,
    new_n996;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n202));
  AND2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT2), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n207), .B1(G155gat), .B2(G162gat), .ZN(new_n208));
  INV_X1    g007(.A(G148gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G141gat), .ZN(new_n210));
  INV_X1    g009(.A(G141gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G148gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT80), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n208), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n210), .A2(new_n212), .A3(KEYINPUT80), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n206), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n203), .B1(new_n207), .B2(new_n204), .ZN(new_n218));
  OR2_X1    g017(.A1(KEYINPUT81), .A2(G141gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(KEYINPUT81), .A2(G141gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(G148gat), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n218), .B1(new_n210), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n202), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G155gat), .ZN(new_n224));
  INV_X1    g023(.A(G162gat), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT2), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G141gat), .B(G148gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n226), .B1(new_n227), .B2(KEYINPUT80), .ZN(new_n228));
  INV_X1    g027(.A(new_n216), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n205), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n221), .A2(new_n210), .ZN(new_n231));
  INV_X1    g030(.A(new_n218), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(KEYINPUT82), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G134gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G127gat), .ZN(new_n236));
  INV_X1    g035(.A(G127gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G134gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(G113gat), .B2(G120gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT68), .B(G120gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G113gat), .ZN(new_n244));
  INV_X1    g043(.A(G113gat), .ZN(new_n245));
  INV_X1    g044(.A(G120gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n247), .A2(new_n241), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n242), .A2(new_n244), .B1(new_n248), .B2(new_n239), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n223), .A2(new_n234), .A3(KEYINPUT4), .A4(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT3), .B1(new_n217), .B2(new_n222), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n242), .A2(new_n244), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n248), .A2(new_n239), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n230), .A2(new_n255), .A3(new_n233), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n251), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G225gat), .A2(G233gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n249), .A2(new_n230), .A3(new_n233), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n250), .A2(new_n257), .A3(new_n258), .A4(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT5), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n254), .B1(new_n217), .B2(new_n222), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(new_n259), .ZN(new_n265));
  INV_X1    g064(.A(new_n258), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n263), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n223), .A2(new_n234), .A3(new_n260), .A4(new_n249), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n259), .A2(KEYINPUT4), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n230), .A2(new_n233), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n249), .B1(new_n272), .B2(KEYINPUT3), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n266), .B1(new_n273), .B2(new_n256), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n271), .A2(new_n274), .A3(new_n263), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n276));
  XOR2_X1   g075(.A(G1gat), .B(G29gat), .Z(new_n277));
  XNOR2_X1  g076(.A(G57gat), .B(G85gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n268), .A2(new_n275), .A3(new_n276), .A4(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G204gat), .ZN(new_n284));
  AND2_X1   g083(.A1(KEYINPUT75), .A2(G197gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(KEYINPUT75), .A2(G197gat), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT75), .ZN(new_n288));
  INV_X1    g087(.A(G197gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(KEYINPUT75), .A2(G197gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(G204gat), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(G211gat), .A2(G218gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(G211gat), .A2(G218gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n294), .A2(KEYINPUT22), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n293), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n297), .B1(new_n293), .B2(new_n298), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G226gat), .A2(G233gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT24), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n306));
  INV_X1    g105(.A(G183gat), .ZN(new_n307));
  INV_X1    g106(.A(G190gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n305), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT23), .ZN(new_n312));
  INV_X1    g111(.A(G169gat), .ZN(new_n313));
  INV_X1    g112(.A(G176gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT23), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(KEYINPUT64), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT64), .ZN(new_n319));
  NOR2_X1   g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n319), .B1(new_n320), .B2(KEYINPUT23), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n310), .B(new_n316), .C1(new_n318), .C2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT25), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT65), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n303), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT24), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n303), .A2(new_n324), .A3(new_n304), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT66), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n328), .B1(G183gat), .B2(G190gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n307), .A2(new_n308), .A3(KEYINPUT66), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n326), .A2(new_n327), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n320), .B1(KEYINPUT23), .B2(new_n311), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT25), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n322), .A2(new_n323), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT26), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n315), .A2(new_n336), .A3(new_n311), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n320), .A2(KEYINPUT26), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n303), .A3(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT27), .B(G183gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(new_n308), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT67), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n342), .A2(KEYINPUT28), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n343), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n340), .A2(new_n345), .A3(new_n308), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n339), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT77), .B1(new_n335), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n337), .A2(new_n303), .A3(new_n338), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n340), .A2(new_n345), .A3(new_n308), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n345), .B1(new_n340), .B2(new_n308), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354));
  AND2_X1   g153(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n354), .B1(new_n355), .B2(G190gat), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n356), .A2(new_n305), .B1(new_n315), .B2(new_n312), .ZN(new_n357));
  INV_X1    g156(.A(new_n321), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n320), .A2(new_n319), .A3(KEYINPUT23), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT25), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n323), .B1(new_n320), .B2(KEYINPUT23), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n316), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n330), .A2(new_n329), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n304), .B1(new_n303), .B2(new_n324), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n363), .B1(new_n366), .B2(new_n327), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n349), .B(new_n353), .C1(new_n361), .C2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n302), .B1(new_n348), .B2(new_n368), .ZN(new_n369));
  XOR2_X1   g168(.A(new_n302), .B(KEYINPUT76), .Z(new_n370));
  NAND2_X1  g169(.A1(new_n322), .A2(new_n323), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n331), .A2(new_n334), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n353), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n370), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n301), .B1(new_n369), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n301), .B1(new_n374), .B2(new_n370), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT29), .B1(new_n348), .B2(new_n368), .ZN(new_n379));
  INV_X1    g178(.A(new_n302), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  XOR2_X1   g180(.A(G8gat), .B(G36gat), .Z(new_n382));
  XOR2_X1   g181(.A(G64gat), .B(G92gat), .Z(new_n383));
  XOR2_X1   g182(.A(new_n382), .B(new_n383), .Z(new_n384));
  NAND3_X1  g183(.A1(new_n377), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT79), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n268), .A2(new_n275), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n282), .A2(new_n276), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n281), .A2(KEYINPUT6), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n387), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT79), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n377), .A2(new_n381), .A3(new_n393), .A4(new_n384), .ZN(new_n394));
  AND4_X1   g193(.A1(new_n283), .A2(new_n386), .A3(new_n392), .A4(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT37), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n377), .A2(new_n381), .A3(new_n396), .ZN(new_n397));
  XOR2_X1   g196(.A(new_n384), .B(KEYINPUT78), .Z(new_n398));
  NOR2_X1   g197(.A1(new_n398), .A2(KEYINPUT38), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n348), .A2(new_n368), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n380), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n285), .A2(new_n286), .A3(new_n284), .ZN(new_n403));
  AOI21_X1  g202(.A(G204gat), .B1(new_n290), .B2(new_n291), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n298), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n296), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n293), .A2(new_n297), .A3(new_n298), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n370), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n335), .A2(new_n347), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n409), .B1(new_n410), .B2(KEYINPUT29), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n402), .A2(new_n408), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT90), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT90), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n402), .A2(new_n414), .A3(new_n408), .A4(new_n411), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n380), .B1(new_n401), .B2(new_n375), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n410), .A2(new_n409), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n301), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n413), .A2(new_n415), .A3(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n400), .B1(new_n419), .B2(new_n396), .ZN(new_n420));
  INV_X1    g219(.A(new_n384), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n397), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n396), .B1(new_n377), .B2(new_n381), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT38), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n395), .A2(new_n420), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n271), .A2(new_n257), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT88), .B(KEYINPUT39), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n266), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n264), .A2(new_n259), .A3(new_n258), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n429), .A2(KEYINPUT39), .ZN(new_n430));
  AOI22_X1  g229(.A1(new_n269), .A2(new_n270), .B1(new_n273), .B2(new_n256), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n430), .B1(new_n431), .B2(new_n258), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT40), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n282), .B1(KEYINPUT89), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n428), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n433), .A2(KEYINPUT89), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n436), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n428), .A2(new_n432), .A3(new_n434), .A4(new_n438), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n437), .A2(new_n439), .B1(new_n387), .B2(new_n282), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT30), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n386), .A2(new_n441), .A3(new_n394), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n398), .B1(new_n377), .B2(new_n381), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n377), .A2(new_n381), .A3(new_n384), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n443), .B1(new_n444), .B2(KEYINPUT30), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G228gat), .ZN(new_n448));
  INV_X1    g247(.A(G233gat), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n211), .A2(G148gat), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n209), .A2(G141gat), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n214), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(new_n216), .A3(new_n226), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n454), .A2(new_n205), .B1(new_n231), .B2(new_n232), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT29), .B1(new_n455), .B2(new_n255), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n450), .B1(new_n456), .B2(new_n408), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n375), .B1(new_n299), .B2(new_n300), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT84), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n408), .A2(KEYINPUT84), .A3(new_n375), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n461), .A3(new_n255), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n457), .B1(new_n462), .B2(new_n272), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT29), .B1(new_n406), .B2(new_n407), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n217), .A2(new_n202), .A3(new_n222), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT82), .B1(new_n230), .B2(new_n233), .ZN(new_n466));
  OAI22_X1  g265(.A1(KEYINPUT3), .A2(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n217), .A2(KEYINPUT3), .A3(new_n222), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n301), .B1(new_n468), .B2(KEYINPUT29), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n450), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(G22gat), .B1(new_n463), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n450), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n255), .A2(new_n458), .B1(new_n223), .B2(new_n234), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n408), .B1(new_n375), .B2(new_n256), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(G22gat), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT3), .B1(new_n458), .B2(new_n459), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n455), .B1(new_n477), .B2(new_n461), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n475), .B(new_n476), .C1(new_n478), .C2(new_n457), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n255), .B1(new_n464), .B2(KEYINPUT84), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n458), .A2(new_n459), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n272), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n457), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n465), .A2(new_n466), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT3), .B1(new_n408), .B2(new_n375), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n469), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n483), .A2(new_n484), .B1(new_n487), .B2(new_n472), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT85), .B1(new_n488), .B2(new_n476), .ZN(new_n489));
  XNOR2_X1  g288(.A(G78gat), .B(G106gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(KEYINPUT31), .B(G50gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n480), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n471), .A2(new_n479), .A3(KEYINPUT85), .A4(new_n492), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n425), .A2(new_n447), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT86), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT85), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n479), .A2(new_n499), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n500), .A2(new_n492), .B1(new_n479), .B2(new_n471), .ZN(new_n501));
  AND4_X1   g300(.A1(KEYINPUT85), .A2(new_n471), .A3(new_n479), .A4(new_n492), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n494), .A2(KEYINPUT86), .A3(new_n495), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n392), .A2(new_n283), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n442), .A2(new_n445), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G227gat), .A2(G233gat), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n254), .B1(new_n373), .B2(new_n353), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n335), .A2(new_n249), .A3(new_n347), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT34), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT72), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n514), .B1(new_n510), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  OAI221_X1 g316(.A(new_n510), .B1(new_n515), .B2(new_n514), .C1(new_n511), .C2(new_n512), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n249), .B1(new_n335), .B2(new_n347), .ZN(new_n519));
  INV_X1    g318(.A(new_n510), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n254), .B(new_n353), .C1(new_n361), .C2(new_n367), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT69), .B(KEYINPUT33), .ZN(new_n523));
  XNOR2_X1  g322(.A(G15gat), .B(G43gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(G71gat), .B(G99gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n523), .B1(new_n527), .B2(KEYINPUT71), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(KEYINPUT71), .B2(new_n527), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n522), .A2(KEYINPUT32), .A3(new_n529), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n517), .A2(new_n518), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n526), .B1(new_n522), .B2(new_n523), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT70), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n522), .A2(KEYINPUT32), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n533), .B1(new_n532), .B2(new_n534), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n531), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT74), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT74), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n531), .B(new_n539), .C1(new_n535), .C2(new_n536), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n530), .B1(new_n535), .B2(new_n536), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n517), .A2(new_n518), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n509), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(KEYINPUT36), .A3(new_n537), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n507), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT87), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n497), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n538), .A2(new_n540), .B1(new_n543), .B2(new_n542), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n546), .B1(new_n551), .B2(new_n509), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(KEYINPUT87), .A3(new_n507), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n496), .A2(new_n544), .A3(new_n537), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT35), .B1(new_n554), .B2(new_n506), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT91), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n442), .A2(new_n445), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT35), .B1(new_n392), .B2(new_n283), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(new_n496), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n541), .A2(new_n544), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n556), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT35), .ZN(new_n562));
  AOI211_X1 g361(.A(new_n388), .B(new_n390), .C1(new_n268), .C2(new_n275), .ZN(new_n563));
  AND4_X1   g362(.A1(new_n276), .A2(new_n268), .A3(new_n275), .A4(new_n282), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n565), .B1(new_n494), .B2(new_n495), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n566), .A2(new_n551), .A3(KEYINPUT91), .A4(new_n557), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n550), .A2(new_n553), .B1(new_n555), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G57gat), .B(G64gat), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g371(.A1(KEYINPUT97), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(G71gat), .B2(G78gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n572), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT21), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(new_n237), .ZN(new_n580));
  XNOR2_X1  g379(.A(G183gat), .B(G211gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G15gat), .B(G22gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT16), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n584), .B1(new_n585), .B2(G1gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(KEYINPUT93), .A2(G8gat), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n586), .B(new_n587), .C1(G1gat), .C2(new_n584), .ZN(new_n588));
  NOR2_X1   g387(.A1(KEYINPUT93), .A2(G8gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n590), .B1(new_n576), .B2(new_n575), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT98), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(new_n224), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n592), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n583), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n595), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n582), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT99), .B(KEYINPUT7), .ZN(new_n600));
  INV_X1    g399(.A(G85gat), .ZN(new_n601));
  INV_X1    g400(.A(G92gat), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n600), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  AOI22_X1  g405(.A1(KEYINPUT8), .A2(new_n606), .B1(new_n601), .B2(new_n602), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G99gat), .B(G106gat), .Z(new_n609));
  OR2_X1    g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(G36gat), .ZN(new_n614));
  AND2_X1   g413(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n615));
  NOR2_X1   g414(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(G29gat), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n618), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n620), .A2(KEYINPUT15), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(KEYINPUT15), .ZN(new_n622));
  XNOR2_X1  g421(.A(G43gat), .B(G50gat), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g425(.A1(G232gat), .A2(G233gat), .ZN(new_n627));
  AOI22_X1  g426(.A1(new_n613), .A2(new_n626), .B1(KEYINPUT41), .B2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n612), .B(KEYINPUT100), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT17), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n626), .B(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n628), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G190gat), .B(G218gat), .ZN(new_n633));
  OAI21_X1  g432(.A(KEYINPUT101), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G134gat), .B(G162gat), .ZN(new_n635));
  OR3_X1    g434(.A1(new_n635), .A2(KEYINPUT41), .A3(new_n627), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n635), .B1(KEYINPUT41), .B2(new_n627), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n632), .B(new_n633), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n638), .A2(new_n639), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT102), .B1(new_n599), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n626), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(new_n590), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(G229gat), .A2(G233gat), .ZN(new_n648));
  INV_X1    g447(.A(new_n590), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n647), .B(new_n648), .C1(new_n631), .C2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT18), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n626), .B(KEYINPUT17), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n646), .B1(new_n653), .B2(new_n590), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n654), .A2(KEYINPUT18), .A3(new_n648), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT95), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n656), .B1(new_n645), .B2(new_n590), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n647), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT94), .B(KEYINPUT13), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(new_n648), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n649), .A2(new_n656), .A3(new_n626), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n652), .A2(new_n655), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G113gat), .B(G141gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(G197gat), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT11), .B(G169gat), .Z(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT12), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT92), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT96), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n652), .A2(new_n655), .A3(new_n662), .A4(new_n668), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT96), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n663), .A2(new_n673), .A3(new_n669), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n671), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n642), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n640), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n596), .A2(new_n598), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(G230gat), .A2(G233gat), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(KEYINPUT106), .Z(new_n682));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n608), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n608), .A2(new_n683), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(new_n609), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(KEYINPUT105), .ZN(new_n687));
  INV_X1    g486(.A(new_n575), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n684), .A2(new_n689), .A3(new_n609), .A4(new_n685), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n687), .A2(new_n610), .A3(new_n688), .A4(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT103), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n612), .A2(new_n692), .A3(new_n575), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT10), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT103), .B1(new_n613), .B2(new_n688), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n691), .A2(new_n693), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n613), .A2(KEYINPUT10), .A3(new_n688), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n682), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n682), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n695), .A2(new_n693), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n699), .B1(new_n700), .B2(new_n691), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(G120gat), .B(G148gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(G176gat), .B(G204gat), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n703), .B(new_n704), .Z(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  OR3_X1    g505(.A1(new_n702), .A2(KEYINPUT107), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n706), .B1(new_n702), .B2(KEYINPUT107), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n644), .A2(new_n675), .A3(new_n680), .A4(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n569), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n505), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT108), .B(G1gat), .Z(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1324gat));
  XOR2_X1   g514(.A(KEYINPUT16), .B(G8gat), .Z(new_n716));
  NAND3_X1  g515(.A1(new_n711), .A2(new_n446), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT42), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n720), .A2(KEYINPUT109), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n711), .A2(new_n446), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n718), .B1(new_n722), .B2(G8gat), .ZN(new_n723));
  INV_X1    g522(.A(new_n717), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n720), .B(KEYINPUT109), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT110), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n721), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(new_n721), .B2(new_n725), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(G1325gat));
  INV_X1    g528(.A(G15gat), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n711), .A2(new_n730), .A3(new_n551), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n569), .A2(new_n552), .A3(new_n710), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n731), .B1(new_n732), .B2(new_n730), .ZN(G1326gat));
  NAND2_X1  g532(.A1(new_n503), .A2(new_n504), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n711), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(KEYINPUT43), .B(G22gat), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1327gat));
  NOR2_X1   g537(.A1(new_n569), .A2(new_n677), .ZN(new_n739));
  INV_X1    g538(.A(new_n709), .ZN(new_n740));
  INV_X1    g539(.A(new_n675), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n740), .A2(new_n741), .A3(new_n679), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(new_n618), .A3(new_n712), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n745), .A2(KEYINPUT111), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(KEYINPUT111), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n677), .A2(KEYINPUT44), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n558), .B1(new_n501), .B2(new_n502), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n446), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT91), .B1(new_n753), .B2(new_n551), .ZN(new_n754));
  AND4_X1   g553(.A1(KEYINPUT91), .A2(new_n566), .A3(new_n551), .A4(new_n557), .ZN(new_n755));
  OAI211_X1 g554(.A(KEYINPUT112), .B(new_n555), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n548), .A2(new_n497), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT112), .B1(new_n568), .B2(new_n555), .ZN(new_n759));
  OAI211_X1 g558(.A(KEYINPUT113), .B(new_n751), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT44), .B1(new_n569), .B2(new_n677), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n555), .B1(new_n754), .B2(new_n755), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n765), .A2(new_n756), .A3(new_n757), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT113), .B1(new_n766), .B2(new_n751), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n742), .ZN(new_n769));
  OAI21_X1  g568(.A(G29gat), .B1(new_n769), .B2(new_n505), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n746), .A2(KEYINPUT45), .A3(new_n747), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n750), .A2(new_n770), .A3(new_n771), .ZN(G1328gat));
  OAI21_X1  g571(.A(G36gat), .B1(new_n769), .B2(new_n557), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n743), .A2(G36gat), .A3(new_n557), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT46), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(G1329gat));
  INV_X1    g575(.A(G43gat), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(new_n743), .B2(new_n560), .ZN(new_n778));
  INV_X1    g577(.A(new_n552), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G43gat), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n778), .B1(new_n769), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g581(.A(G50gat), .B1(new_n769), .B2(new_n496), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT48), .ZN(new_n784));
  AOI211_X1 g583(.A(G50gat), .B(new_n734), .C1(new_n744), .C2(KEYINPUT114), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n744), .A2(KEYINPUT114), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n768), .A2(new_n735), .A3(new_n742), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n789), .A2(G50gat), .B1(new_n785), .B2(new_n786), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n790), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g590(.A1(new_n709), .A2(new_n675), .ZN(new_n792));
  AND4_X1   g591(.A1(new_n644), .A2(new_n766), .A3(new_n680), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n712), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n446), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n797));
  XOR2_X1   g596(.A(KEYINPUT49), .B(G64gat), .Z(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n796), .B2(new_n798), .ZN(G1333gat));
  XNOR2_X1  g598(.A(new_n551), .B(KEYINPUT115), .ZN(new_n800));
  AOI21_X1  g599(.A(G71gat), .B1(new_n793), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n779), .A2(G71gat), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n801), .B1(new_n793), .B2(new_n803), .ZN(new_n804));
  XOR2_X1   g603(.A(new_n804), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g604(.A1(new_n793), .A2(new_n735), .ZN(new_n806));
  XNOR2_X1  g605(.A(KEYINPUT116), .B(G78gat), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n806), .B(new_n807), .ZN(G1335gat));
  NAND2_X1  g607(.A1(new_n741), .A2(new_n599), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(new_n677), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n810), .B1(new_n758), .B2(new_n759), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n766), .A2(KEYINPUT51), .A3(new_n810), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n815), .A2(new_n601), .A3(new_n712), .A4(new_n740), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n809), .A2(new_n709), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n768), .A2(new_n712), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n816), .B1(new_n819), .B2(new_n601), .ZN(G1336gat));
  NOR3_X1   g619(.A1(new_n709), .A2(G92gat), .A3(new_n557), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT52), .B1(new_n815), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n768), .A2(new_n446), .A3(new_n817), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n824), .B2(new_n602), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n811), .A2(new_n826), .A3(KEYINPUT51), .ZN(new_n827));
  AOI21_X1  g626(.A(KEYINPUT51), .B1(new_n811), .B2(new_n826), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI22_X1  g628(.A1(new_n823), .A2(G92gat), .B1(new_n829), .B2(new_n821), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n825), .B1(new_n830), .B2(new_n831), .ZN(G1337gat));
  NOR3_X1   g631(.A1(new_n709), .A2(G99gat), .A3(new_n560), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(KEYINPUT119), .Z(new_n834));
  NAND2_X1  g633(.A1(new_n815), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n768), .A2(new_n817), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT118), .B1(new_n836), .B2(new_n552), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(G99gat), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n836), .A2(KEYINPUT118), .A3(new_n552), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(G1338gat));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n735), .B(new_n817), .C1(new_n762), .C2(new_n767), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(G106gat), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n709), .A2(G106gat), .A3(new_n496), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  OR3_X1    g644(.A1(new_n827), .A2(new_n828), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n841), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n845), .B1(new_n813), .B2(new_n814), .ZN(new_n848));
  INV_X1    g647(.A(new_n496), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n849), .B(new_n817), .C1(new_n762), .C2(new_n767), .ZN(new_n850));
  AOI211_X1 g649(.A(KEYINPUT53), .B(new_n848), .C1(new_n850), .C2(G106gat), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT120), .B1(new_n847), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(G106gat), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n848), .A2(KEYINPUT53), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856));
  AOI22_X1  g655(.A1(G106gat), .A2(new_n842), .B1(new_n829), .B2(new_n844), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n855), .B(new_n856), .C1(new_n857), .C2(new_n841), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n852), .A2(new_n858), .ZN(G1339gat));
  NAND2_X1  g658(.A1(new_n696), .A2(new_n697), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n699), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n696), .A2(new_n682), .A3(new_n697), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(KEYINPUT54), .A3(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n705), .B1(new_n698), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT55), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n702), .A2(new_n705), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n863), .A2(KEYINPUT55), .A3(new_n865), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n675), .A2(new_n868), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n654), .A2(new_n648), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n660), .B1(new_n658), .B2(new_n661), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n667), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n672), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n707), .A2(new_n708), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n643), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n643), .A2(new_n875), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n599), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n644), .A2(new_n741), .A3(new_n680), .A4(new_n709), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(new_n735), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n446), .A2(new_n505), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n551), .A3(new_n886), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n887), .A2(new_n245), .A3(new_n741), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n884), .A2(new_n505), .A3(new_n554), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n889), .A2(new_n557), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n675), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n888), .B1(new_n891), .B2(new_n245), .ZN(G1340gat));
  NOR2_X1   g691(.A1(new_n709), .A2(new_n243), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(G120gat), .B1(new_n887), .B2(new_n709), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1341gat));
  NAND3_X1  g695(.A1(new_n890), .A2(new_n237), .A3(new_n679), .ZN(new_n897));
  OAI21_X1  g696(.A(G127gat), .B1(new_n887), .B2(new_n599), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1342gat));
  NOR2_X1   g698(.A1(new_n677), .A2(new_n446), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n889), .A2(new_n235), .A3(new_n900), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n901), .A2(KEYINPUT56), .ZN(new_n902));
  OAI21_X1  g701(.A(G134gat), .B1(new_n887), .B2(new_n677), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(KEYINPUT56), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(G1343gat));
  NOR2_X1   g704(.A1(new_n779), .A2(new_n496), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n883), .A2(new_n712), .A3(new_n557), .A4(new_n906), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n907), .A2(G141gat), .A3(new_n741), .ZN(new_n908));
  INV_X1    g707(.A(new_n886), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n779), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT57), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n734), .A2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT121), .ZN(new_n914));
  OAI22_X1  g713(.A1(new_n877), .A2(new_n914), .B1(new_n879), .B2(new_n878), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n877), .A2(new_n914), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n599), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n913), .B1(new_n917), .B2(new_n882), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n496), .B1(new_n881), .B2(new_n882), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n919), .A2(KEYINPUT57), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n675), .B(new_n910), .C1(new_n918), .C2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n219), .A2(new_n220), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n908), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g722(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n923), .B(new_n925), .ZN(G1344gat));
  NOR3_X1   g725(.A1(new_n907), .A2(G148gat), .A3(new_n709), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT123), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n910), .B1(new_n918), .B2(new_n920), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(new_n709), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n930), .A2(KEYINPUT59), .A3(new_n209), .ZN(new_n931));
  XNOR2_X1  g730(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n911), .B1(new_n883), .B2(new_n849), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n734), .A2(KEYINPUT57), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n935), .B1(new_n881), .B2(new_n882), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n910), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n709), .B1(new_n938), .B2(KEYINPUT125), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n937), .B(new_n939), .C1(KEYINPUT125), .C2(new_n938), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n932), .B1(new_n940), .B2(G148gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n928), .B1(new_n931), .B2(new_n941), .ZN(G1345gat));
  OAI21_X1  g741(.A(G155gat), .B1(new_n929), .B2(new_n599), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n679), .A2(new_n224), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n907), .B2(new_n944), .ZN(G1346gat));
  OAI21_X1  g744(.A(G162gat), .B1(new_n929), .B2(new_n677), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n884), .A2(new_n505), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n947), .A2(new_n225), .A3(new_n900), .A4(new_n906), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(G1347gat));
  NOR2_X1   g748(.A1(new_n557), .A2(new_n712), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n800), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n885), .A2(new_n951), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n952), .A2(new_n313), .A3(new_n741), .ZN(new_n953));
  NOR4_X1   g752(.A1(new_n884), .A2(new_n712), .A3(new_n557), .A4(new_n554), .ZN(new_n954));
  AOI21_X1  g753(.A(G169gat), .B1(new_n954), .B2(new_n675), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n953), .A2(new_n955), .ZN(G1348gat));
  OAI21_X1  g755(.A(G176gat), .B1(new_n952), .B2(new_n709), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n954), .A2(new_n314), .A3(new_n740), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1349gat));
  OAI21_X1  g758(.A(G183gat), .B1(new_n952), .B2(new_n599), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n954), .A2(new_n340), .A3(new_n679), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g762(.A1(new_n954), .A2(new_n308), .A3(new_n643), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n883), .A2(new_n734), .A3(new_n643), .A4(new_n951), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n965), .B1(new_n966), .B2(G190gat), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n966), .A2(new_n965), .A3(G190gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT126), .ZN(G1351gat));
  AND2_X1   g769(.A1(new_n883), .A2(new_n950), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n971), .A2(new_n906), .ZN(new_n972));
  AOI21_X1  g771(.A(G197gat), .B1(new_n972), .B2(new_n675), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n883), .A2(new_n934), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n552), .A2(new_n950), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  OAI211_X1 g775(.A(new_n974), .B(new_n976), .C1(new_n911), .C2(new_n919), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n977), .A2(new_n289), .A3(new_n741), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n973), .A2(new_n978), .ZN(G1352gat));
  NAND4_X1  g778(.A1(new_n971), .A2(new_n284), .A3(new_n740), .A4(new_n906), .ZN(new_n980));
  XOR2_X1   g779(.A(new_n980), .B(KEYINPUT62), .Z(new_n981));
  OAI21_X1  g780(.A(G204gat), .B1(new_n977), .B2(new_n709), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1353gat));
  INV_X1    g782(.A(G211gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n972), .A2(new_n984), .A3(new_n679), .ZN(new_n985));
  NOR4_X1   g784(.A1(new_n933), .A2(new_n599), .A3(new_n936), .A4(new_n975), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n984), .B1(new_n986), .B2(KEYINPUT127), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n988), .B1(new_n977), .B2(new_n599), .ZN(new_n989));
  AOI21_X1  g788(.A(KEYINPUT63), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NAND4_X1  g789(.A1(new_n937), .A2(KEYINPUT127), .A3(new_n679), .A4(new_n976), .ZN(new_n991));
  AND4_X1   g790(.A1(KEYINPUT63), .A2(new_n991), .A3(new_n989), .A4(G211gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n985), .B1(new_n990), .B2(new_n992), .ZN(G1354gat));
  INV_X1    g792(.A(G218gat), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n972), .A2(new_n994), .A3(new_n643), .ZN(new_n995));
  OAI21_X1  g794(.A(G218gat), .B1(new_n977), .B2(new_n677), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(G1355gat));
endmodule


