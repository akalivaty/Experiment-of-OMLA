//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n446, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n544,
    new_n546, new_n547, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n608, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NAND4_X1  g032(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT67), .Z(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  AOI22_X1  g036(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n465), .A2(new_n467), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(G137), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n464), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n471), .A2(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n468), .A2(new_n473), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n468), .A2(G2105), .ZN(new_n480));
  AOI22_X1  g055(.A1(G124), .A2(new_n479), .B1(new_n480), .B2(G136), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT68), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n481), .A2(new_n485), .ZN(G162));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G114), .C2(new_n473), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n465), .A2(new_n467), .A3(G126), .A4(G2105), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n472), .A2(G138), .A3(new_n473), .A4(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n473), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n491), .B2(new_n492), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n490), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  AND2_X1   g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(KEYINPUT70), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT6), .A3(G651), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n501), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n501), .B2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n507), .A2(G88), .B1(new_n510), .B2(G651), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n512), .B1(new_n504), .B2(new_n506), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n511), .A2(new_n514), .ZN(G166));
  XNOR2_X1  g090(.A(KEYINPUT71), .B(G51), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT5), .B(G543), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT72), .B(G89), .ZN(new_n519));
  AND3_X1   g094(.A1(new_n505), .A2(KEYINPUT6), .A3(G651), .ZN(new_n520));
  AOI21_X1  g095(.A(KEYINPUT6), .B1(new_n505), .B2(G651), .ZN(new_n521));
  OAI211_X1 g096(.A(new_n518), .B(new_n519), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(G63), .A2(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT7), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n526), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n518), .A2(new_n523), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n517), .A2(new_n522), .A3(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  NAND2_X1  g105(.A1(new_n513), .A2(G52), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n518), .B(G90), .C1(new_n520), .C2(new_n521), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n531), .B(new_n532), .C1(new_n533), .C2(new_n503), .ZN(G301));
  INV_X1    g109(.A(G301), .ZN(G171));
  AOI22_X1  g110(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(new_n503), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n513), .A2(G43), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT73), .B(G81), .Z(new_n539));
  NAND2_X1  g114(.A1(new_n507), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  AND3_X1   g118(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G36), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n544), .A2(new_n547), .ZN(G188));
  INV_X1    g123(.A(KEYINPUT75), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n507), .A2(G91), .ZN(new_n550));
  OAI21_X1  g125(.A(G65), .B1(new_n499), .B2(new_n500), .ZN(new_n551));
  NAND2_X1  g126(.A1(G78), .A2(G543), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n551), .A2(KEYINPUT74), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  AOI21_X1  g129(.A(KEYINPUT74), .B1(new_n551), .B2(new_n552), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n550), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  AND3_X1   g132(.A1(new_n513), .A2(new_n557), .A3(G53), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n557), .B1(new_n513), .B2(G53), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n549), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g136(.A(G543), .B1(new_n520), .B2(new_n521), .ZN(new_n562));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT9), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n513), .A2(new_n557), .A3(G53), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n551), .A2(new_n552), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n569), .A2(G651), .A3(new_n553), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n566), .A2(new_n570), .A3(KEYINPUT75), .A4(new_n550), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n561), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G299));
  NAND2_X1  g148(.A1(new_n511), .A2(new_n514), .ZN(G303));
  NAND2_X1  g149(.A1(new_n513), .A2(G49), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n518), .B(G87), .C1(new_n520), .C2(new_n521), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G288));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n501), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n513), .A2(G48), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n518), .B(G86), .C1(new_n520), .C2(new_n521), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(G72), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G60), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n501), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(G47), .B2(new_n513), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n507), .A2(G85), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT76), .Z(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n501), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(G54), .B2(new_n513), .ZN(new_n597));
  AND3_X1   g172(.A1(new_n507), .A2(KEYINPUT10), .A3(G92), .ZN(new_n598));
  AOI21_X1  g173(.A(KEYINPUT10), .B1(new_n507), .B2(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT77), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n593), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n593), .B1(new_n602), .B2(G868), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n572), .B2(G868), .ZN(G297));
  OAI21_X1  g181(.A(new_n605), .B1(new_n572), .B2(G868), .ZN(G280));
  NOR2_X1   g182(.A1(new_n601), .A2(G559), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(G860), .B2(new_n602), .ZN(G148));
  OAI21_X1  g184(.A(G868), .B1(new_n601), .B2(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G2100), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n480), .A2(G2104), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT12), .Z(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT13), .Z(new_n617));
  NOR2_X1   g192(.A1(new_n613), .A2(G2100), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n479), .A2(G123), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n473), .A2(G111), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n480), .A2(G135), .ZN(new_n623));
  AND2_X1   g198(.A1(new_n623), .A2(KEYINPUT79), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n623), .A2(KEYINPUT79), .ZN(new_n625));
  OAI221_X1 g200(.A(new_n620), .B1(new_n621), .B2(new_n622), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2096), .Z(new_n627));
  OAI211_X1 g202(.A(new_n619), .B(new_n627), .C1(new_n617), .C2(new_n614), .ZN(G156));
  XOR2_X1   g203(.A(KEYINPUT80), .B(KEYINPUT14), .Z(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2427), .B(G2430), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n631), .B2(new_n632), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n634), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  AND3_X1   g217(.A1(new_n641), .A2(G14), .A3(new_n642), .ZN(G401));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT81), .Z(new_n645));
  NOR2_X1   g220(.A1(G2072), .A2(G2078), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n444), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(KEYINPUT17), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n648), .B(new_n650), .C1(new_n645), .C2(new_n651), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n649), .B(new_n644), .C1(new_n444), .C2(new_n646), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT18), .Z(new_n654));
  NAND3_X1  g229(.A1(new_n651), .A2(new_n645), .A3(new_n649), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n652), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2096), .B(G2100), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1991), .B(G1996), .Z(new_n659));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT82), .ZN(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT83), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n661), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(new_n666), .B2(new_n665), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT20), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n665), .A2(new_n661), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n663), .A2(new_n664), .ZN(new_n671));
  MUX2_X1   g246(.A(new_n670), .B(new_n661), .S(new_n671), .Z(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n673), .B1(new_n669), .B2(new_n672), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n659), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n676), .ZN(new_n678));
  INV_X1    g253(.A(new_n659), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n678), .A2(new_n679), .A3(new_n674), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  AND3_X1   g256(.A1(new_n677), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n681), .B1(new_n677), .B2(new_n680), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(G229));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  NOR2_X1   g260(.A1(G171), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(G5), .B2(new_n685), .ZN(new_n687));
  INV_X1    g262(.A(G1961), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT31), .B(G11), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT101), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT102), .B(G28), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n692), .A2(KEYINPUT30), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(KEYINPUT30), .ZN(new_n694));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI221_X1 g271(.A(new_n691), .B1(new_n693), .B2(new_n696), .C1(new_n626), .C2(new_n695), .ZN(new_n697));
  INV_X1    g272(.A(G2084), .ZN(new_n698));
  NAND2_X1  g273(.A1(G160), .A2(G29), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT24), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n700), .A2(G34), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n695), .B1(new_n700), .B2(G34), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n697), .B1(new_n698), .B2(new_n703), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n687), .A2(new_n688), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n695), .A2(G35), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G162), .B2(new_n695), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT29), .B(G2090), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  AND4_X1   g284(.A1(new_n689), .A2(new_n704), .A3(new_n705), .A4(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT98), .ZN(new_n711));
  NAND4_X1  g286(.A1(new_n465), .A2(new_n467), .A3(G129), .A4(G2105), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT97), .ZN(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT26), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n465), .A2(new_n467), .A3(G141), .A4(new_n473), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n475), .A2(G105), .ZN(new_n718));
  AND3_X1   g293(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n711), .B1(new_n713), .B2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n713), .A2(new_n719), .A3(new_n711), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(new_n695), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(KEYINPUT99), .ZN(new_n725));
  INV_X1    g300(.A(G32), .ZN(new_n726));
  AOI21_X1  g301(.A(KEYINPUT99), .B1(new_n695), .B2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n725), .B1(new_n724), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT27), .B(G1996), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n685), .A2(G21), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G168), .B2(new_n685), .ZN(new_n734));
  INV_X1    g309(.A(G1966), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n695), .A2(G27), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G164), .B2(new_n695), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(new_n443), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n710), .A2(new_n732), .A3(new_n736), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n685), .A2(G20), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT23), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n572), .B2(new_n685), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1956), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n695), .A2(G33), .ZN(new_n746));
  NAND2_X1  g321(.A1(G115), .A2(G2104), .ZN(new_n747));
  INV_X1    g322(.A(G127), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n468), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G2105), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT25), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n480), .A2(G139), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n750), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT95), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n746), .B1(new_n758), .B2(G29), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(new_n442), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT96), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n725), .B(new_n730), .C1(new_n724), .C2(new_n728), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n703), .A2(new_n698), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n759), .B2(new_n442), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(KEYINPUT100), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT96), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n760), .B(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT100), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n768), .A2(new_n769), .A3(new_n762), .A4(new_n764), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n745), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n685), .A2(G22), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G166), .B2(new_n685), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G1971), .ZN(new_n775));
  NOR2_X1   g350(.A1(G6), .A2(G16), .ZN(new_n776));
  INV_X1    g351(.A(G305), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(G16), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT32), .B(G1981), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n775), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(G288), .A2(KEYINPUT87), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT87), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n575), .A2(new_n576), .A3(new_n783), .A4(new_n577), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  MUX2_X1   g360(.A(G23), .B(new_n785), .S(G16), .Z(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT33), .B(G1976), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n781), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT34), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n781), .A2(new_n788), .A3(KEYINPUT34), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G107), .B2(new_n473), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT84), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n480), .A2(G131), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n479), .A2(G119), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n803), .A2(new_n695), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G25), .B2(new_n695), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT35), .B(G1991), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT85), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n805), .A2(new_n807), .B1(KEYINPUT88), .B2(KEYINPUT36), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n685), .A2(G24), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT86), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G290), .B2(G16), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1986), .ZN(new_n813));
  AND3_X1   g388(.A1(new_n808), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  AND3_X1   g389(.A1(new_n793), .A2(new_n795), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n795), .B1(new_n793), .B2(new_n814), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n601), .A2(G16), .ZN(new_n818));
  INV_X1    g393(.A(G4), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(G16), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n820), .A2(G1348), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n685), .A2(G19), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n542), .B2(new_n685), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT89), .B(G1341), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT90), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n823), .B(new_n825), .Z(new_n826));
  NOR2_X1   g401(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(G116), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n464), .B1(new_n828), .B2(G2105), .ZN(new_n829));
  OAI21_X1  g404(.A(KEYINPUT91), .B1(G104), .B2(G2105), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NOR3_X1   g406(.A1(KEYINPUT91), .A2(G104), .A3(G2105), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n829), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n465), .A2(new_n467), .A3(G140), .A4(new_n473), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n465), .A2(new_n467), .A3(G128), .A4(G2105), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G29), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT92), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n695), .A2(G26), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT28), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT93), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G2067), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n820), .A2(G1348), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n827), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(KEYINPUT94), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT94), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n827), .A2(new_n843), .A3(new_n847), .A4(new_n844), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n772), .A2(new_n817), .A3(KEYINPUT103), .A4(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT103), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n745), .A2(new_n771), .A3(new_n846), .A4(new_n848), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n793), .A2(new_n814), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(new_n794), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n793), .A2(new_n795), .A3(new_n814), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n851), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n850), .A2(new_n857), .ZN(G311));
  NAND3_X1  g433(.A1(new_n772), .A2(new_n817), .A3(new_n849), .ZN(G150));
  XOR2_X1   g434(.A(KEYINPUT107), .B(G860), .Z(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(G67), .ZN(new_n862));
  OR2_X1    g437(.A1(KEYINPUT5), .A2(G543), .ZN(new_n863));
  NAND2_X1  g438(.A1(KEYINPUT5), .A2(G543), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(G80), .A2(G543), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT104), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT104), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n869), .B(new_n866), .C1(new_n501), .C2(new_n862), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(G651), .A3(new_n870), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n518), .B(G93), .C1(new_n520), .C2(new_n521), .ZN(new_n872));
  OAI211_X1 g447(.A(G55), .B(G543), .C1(new_n520), .C2(new_n521), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT105), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n874), .B1(new_n872), .B2(new_n873), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n871), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(KEYINPUT106), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT106), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n879), .B(new_n871), .C1(new_n875), .C2(new_n876), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n542), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n877), .A2(new_n541), .A3(KEYINPUT106), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n602), .A2(G559), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT39), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n861), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n887), .B2(new_n886), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n877), .A2(new_n861), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n890), .B(KEYINPUT37), .Z(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(G145));
  NAND2_X1  g467(.A1(new_n480), .A2(G142), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n479), .A2(G130), .ZN(new_n894));
  OR2_X1    g469(.A1(G106), .A2(G2105), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n895), .B(G2104), .C1(G118), .C2(new_n473), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n616), .ZN(new_n898));
  INV_X1    g473(.A(new_n836), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n497), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n836), .A2(new_n490), .A3(new_n494), .A4(new_n496), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(new_n721), .A3(new_n722), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n713), .A2(new_n719), .A3(new_n711), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n901), .B(new_n900), .C1(new_n904), .C2(new_n720), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n756), .A2(new_n757), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n713), .A2(new_n719), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n900), .A2(new_n713), .A3(new_n719), .A4(new_n901), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n754), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n802), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n907), .A2(new_n802), .A3(new_n911), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n898), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n914), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n916), .A2(new_n616), .A3(new_n912), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n897), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n626), .B(G160), .ZN(new_n919));
  XOR2_X1   g494(.A(new_n919), .B(G162), .Z(new_n920));
  OAI21_X1  g495(.A(new_n616), .B1(new_n916), .B2(new_n912), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n913), .A2(new_n898), .A3(new_n914), .ZN(new_n922));
  INV_X1    g497(.A(new_n897), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n918), .A2(new_n920), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n918), .A2(KEYINPUT108), .A3(new_n920), .A4(new_n924), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n920), .B1(new_n918), .B2(new_n924), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n930), .A2(G37), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n929), .A2(KEYINPUT40), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT40), .B1(new_n929), .B2(new_n931), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(G395));
  OR2_X1    g509(.A1(new_n877), .A2(G868), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n785), .A2(G290), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n589), .A2(new_n590), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(new_n784), .A3(new_n782), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT111), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT111), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n937), .A2(new_n939), .A3(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(G303), .B(G305), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n941), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n944), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n946), .A2(KEYINPUT111), .A3(new_n940), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT42), .ZN(new_n949));
  OR2_X1    g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(KEYINPUT112), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT41), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n561), .A2(KEYINPUT109), .A3(new_n571), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n600), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT109), .B1(new_n561), .B2(new_n571), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI211_X1 g532(.A(KEYINPUT109), .B(new_n600), .C1(new_n561), .C2(new_n571), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n953), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n572), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n961), .A2(new_n600), .A3(new_n954), .ZN(new_n962));
  INV_X1    g537(.A(new_n958), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(new_n963), .A3(KEYINPUT41), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n959), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n608), .B(new_n883), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(KEYINPUT110), .A3(new_n966), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n965), .A2(new_n966), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n962), .A2(new_n963), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n969), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n952), .B(new_n967), .C1(new_n968), .C2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT112), .B1(new_n950), .B2(new_n951), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n972), .B(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n936), .B1(new_n974), .B2(G868), .ZN(G295));
  AOI21_X1  g550(.A(new_n936), .B1(new_n974), .B2(G868), .ZN(G331));
  INV_X1    g551(.A(new_n970), .ZN(new_n977));
  XNOR2_X1  g552(.A(G168), .B(G301), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n881), .A2(new_n882), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n978), .B1(new_n881), .B2(new_n882), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT114), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n978), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n883), .A2(KEYINPUT114), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n977), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n980), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n881), .A2(new_n882), .A3(new_n978), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n959), .A2(new_n964), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n985), .A2(new_n948), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G37), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n985), .A2(new_n989), .A3(KEYINPUT116), .A4(new_n948), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n945), .A2(new_n995), .A3(new_n947), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n995), .B1(new_n945), .B2(new_n947), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n959), .A2(new_n964), .A3(new_n988), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n986), .A2(KEYINPUT114), .A3(new_n987), .ZN(new_n1001));
  INV_X1    g576(.A(new_n984), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n970), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n999), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n992), .A2(new_n993), .A3(new_n994), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT43), .ZN(new_n1006));
  AOI21_X1  g581(.A(G37), .B1(new_n990), .B2(new_n991), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n959), .A2(new_n1001), .A3(new_n1002), .A4(new_n964), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(new_n970), .B2(new_n988), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n999), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT43), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1007), .A2(new_n1010), .A3(new_n1011), .A4(new_n994), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1006), .A2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g588(.A(KEYINPUT113), .B(KEYINPUT44), .Z(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1007), .A2(new_n1011), .A3(new_n994), .A4(new_n1004), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n1007), .A2(new_n994), .A3(new_n1010), .ZN(new_n1017));
  OAI211_X1 g592(.A(KEYINPUT44), .B(new_n1016), .C1(new_n1017), .C2(new_n1011), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1015), .A2(new_n1018), .ZN(G397));
  INV_X1    g594(.A(G1384), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT45), .B1(new_n497), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n470), .A2(G2105), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1022), .A2(G40), .A3(new_n476), .A4(new_n474), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  OR3_X1    g600(.A1(new_n1025), .A2(KEYINPUT117), .A3(G1996), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT117), .B1(new_n1025), .B2(G1996), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g603(.A(new_n1028), .B(KEYINPUT46), .Z(new_n1029));
  INV_X1    g604(.A(new_n1025), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n836), .B(G2067), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1030), .B1(new_n908), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT47), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1028), .A2(new_n721), .A3(new_n722), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1031), .B1(G1996), .B2(new_n908), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(new_n1025), .B2(new_n1036), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n803), .A2(new_n807), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n803), .A2(new_n807), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1025), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1025), .A2(G1986), .A3(G290), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1041), .B(KEYINPUT48), .ZN(new_n1042));
  OR3_X1    g617(.A1(new_n1037), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n1039), .B(KEYINPUT127), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1037), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n836), .A2(G2067), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1030), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1034), .A2(new_n1043), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n1020), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n1024), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n735), .B1(new_n1052), .B2(new_n1021), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n497), .A2(new_n1020), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT50), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT50), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n497), .A2(new_n1056), .A3(new_n1020), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1055), .A2(new_n698), .A3(new_n1024), .A4(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1053), .A2(G168), .A3(new_n1058), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1059), .A2(G8), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1053), .A2(new_n1058), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G286), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1050), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1059), .A2(new_n1050), .A3(G8), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT62), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1062), .A2(G8), .A3(new_n1059), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1064), .B1(new_n1066), .B2(KEYINPUT51), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT62), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G8), .ZN(new_n1070));
  INV_X1    g645(.A(G1971), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1052), .B2(new_n1021), .ZN(new_n1072));
  INV_X1    g647(.A(G2090), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1055), .A2(new_n1073), .A3(new_n1024), .A4(new_n1057), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1070), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n1077));
  NOR3_X1   g652(.A1(G166), .A2(new_n1077), .A3(new_n1070), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1076), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n782), .A2(G1976), .A3(new_n784), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(G8), .B1(new_n1054), .B2(new_n1023), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT52), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n497), .A2(new_n1020), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n1024), .ZN(new_n1087));
  INV_X1    g662(.A(G1976), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT52), .B1(G288), .B2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1087), .A2(new_n1082), .A3(G8), .A4(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1085), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(G305), .A2(G1981), .ZN(new_n1092));
  INV_X1    g667(.A(G1981), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n582), .A2(new_n1093), .A3(new_n583), .A4(new_n584), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT49), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT118), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1092), .A2(new_n1098), .A3(KEYINPUT49), .A4(new_n1094), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1084), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1091), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1080), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1075), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1081), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT45), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1054), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1108), .A2(new_n443), .A3(new_n1024), .A4(new_n1051), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1055), .A2(new_n1024), .A3(new_n1057), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1106), .A2(new_n1109), .B1(new_n1110), .B2(new_n688), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1051), .A2(new_n1024), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1112), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n1108), .ZN(new_n1113));
  AOI21_X1  g688(.A(G301), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1105), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1065), .A2(new_n1069), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1118));
  NOR2_X1   g693(.A1(G288), .A2(G1976), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1118), .A2(new_n1119), .B1(new_n1093), .B2(new_n777), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1118), .A2(new_n1085), .A3(new_n1090), .ZN(new_n1121));
  OAI22_X1  g696(.A1(new_n1120), .A2(new_n1084), .B1(new_n1121), .B2(new_n1104), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1075), .A2(new_n1103), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  AOI211_X1 g699(.A(new_n1070), .B(G286), .C1(new_n1053), .C2(new_n1058), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(KEYINPUT63), .A3(new_n1104), .A4(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1081), .A2(new_n1102), .A3(new_n1104), .A4(new_n1125), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT63), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1122), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1067), .A2(new_n1105), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1109), .A2(new_n1106), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1110), .A2(new_n688), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1133), .A2(new_n1113), .A3(new_n1134), .A4(G301), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1111), .A2(KEYINPUT124), .A3(G301), .A4(new_n1113), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1132), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT125), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1114), .A2(new_n1140), .ZN(new_n1141));
  AOI211_X1 g716(.A(KEYINPUT125), .B(G301), .C1(new_n1111), .C2(new_n1113), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1139), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1115), .A2(new_n1135), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n1132), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1131), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(G1956), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1110), .A2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(KEYINPUT56), .B(G2072), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1112), .A2(new_n1108), .A3(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n566), .A2(new_n570), .A3(new_n550), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT57), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1151), .B(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1148), .A2(new_n1150), .A3(new_n1153), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1087), .A2(G2067), .ZN(new_n1155));
  INV_X1    g730(.A(G1348), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1110), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1154), .A2(new_n1158), .A3(new_n602), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1159), .B1(new_n1153), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT60), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n602), .B1(new_n1158), .B2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1155), .A2(new_n1157), .A3(new_n601), .A4(KEYINPUT60), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1163), .A2(KEYINPUT123), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT123), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1166), .B(new_n602), .C1(new_n1158), .C2(new_n1162), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1158), .A2(new_n1162), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1170), .A2(KEYINPUT122), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1154), .B(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT59), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1173), .A2(KEYINPUT120), .ZN(new_n1174));
  MUX2_X1   g749(.A(new_n1174), .B(new_n1173), .S(KEYINPUT121), .Z(new_n1175));
  XOR2_X1   g750(.A(KEYINPUT58), .B(G1341), .Z(new_n1176));
  NAND2_X1  g751(.A1(new_n1087), .A2(new_n1176), .ZN(new_n1177));
  XOR2_X1   g752(.A(KEYINPUT119), .B(G1996), .Z(new_n1178));
  INV_X1    g753(.A(new_n1178), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1108), .A2(new_n1024), .A3(new_n1051), .A4(new_n1179), .ZN(new_n1180));
  AOI211_X1 g755(.A(new_n541), .B(new_n1175), .C1(new_n1177), .C2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n542), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1181), .B1(new_n1183), .B2(new_n1174), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1172), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1161), .B1(new_n1169), .B2(new_n1185), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1117), .B(new_n1130), .C1(new_n1146), .C2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n1188));
  XNOR2_X1  g763(.A(G290), .B(G1986), .ZN(new_n1189));
  AOI211_X1 g764(.A(new_n1040), .B(new_n1037), .C1(new_n1030), .C2(new_n1189), .ZN(new_n1190));
  AND3_X1   g765(.A1(new_n1187), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1188), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1049), .B1(new_n1191), .B2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g768(.A(G319), .ZN(new_n1195));
  NOR3_X1   g769(.A1(G401), .A2(new_n1195), .A3(G227), .ZN(new_n1196));
  OAI21_X1  g770(.A(new_n1196), .B1(new_n682), .B2(new_n683), .ZN(new_n1197));
  AOI21_X1  g771(.A(new_n1197), .B1(new_n929), .B2(new_n931), .ZN(new_n1198));
  AND2_X1   g772(.A1(new_n1198), .A2(new_n1013), .ZN(G308));
  NAND2_X1  g773(.A1(new_n1198), .A2(new_n1013), .ZN(G225));
endmodule


