

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725;

  XNOR2_X1 U364 ( .A(n441), .B(G107), .ZN(n464) );
  OR2_X2 U365 ( .A1(n544), .A2(n656), .ZN(n498) );
  XNOR2_X2 U366 ( .A(n393), .B(KEYINPUT22), .ZN(n549) );
  NOR2_X2 U367 ( .A1(n544), .A2(n347), .ZN(n393) );
  NOR2_X2 U368 ( .A1(n541), .A2(n719), .ZN(n542) );
  XNOR2_X2 U369 ( .A(G110), .B(G104), .ZN(n441) );
  XNOR2_X2 U370 ( .A(n405), .B(n490), .ZN(n690) );
  XNOR2_X2 U371 ( .A(n407), .B(n406), .ZN(n490) );
  NOR2_X1 U372 ( .A1(n651), .A2(n650), .ZN(n388) );
  NOR2_X1 U373 ( .A1(G953), .A2(n670), .ZN(n673) );
  XNOR2_X1 U374 ( .A(n540), .B(n539), .ZN(n719) );
  XNOR2_X1 U375 ( .A(n438), .B(n346), .ZN(n533) );
  XNOR2_X1 U376 ( .A(n445), .B(n444), .ZN(n571) );
  XNOR2_X1 U377 ( .A(n474), .B(n391), .ZN(n517) );
  XNOR2_X1 U378 ( .A(n443), .B(n442), .ZN(n604) );
  INV_X2 U379 ( .A(KEYINPUT68), .ZN(n399) );
  XNOR2_X1 U380 ( .A(n483), .B(n482), .ZN(n576) );
  XNOR2_X2 U381 ( .A(n532), .B(KEYINPUT35), .ZN(n717) );
  NOR2_X2 U382 ( .A1(n572), .A2(n531), .ZN(n532) );
  XNOR2_X2 U383 ( .A(n705), .B(G146), .ZN(n492) );
  XNOR2_X2 U384 ( .A(n459), .B(n400), .ZN(n705) );
  NAND2_X1 U385 ( .A1(n343), .A2(n416), .ZN(n414) );
  XNOR2_X1 U386 ( .A(n480), .B(n380), .ZN(n482) );
  NOR2_X1 U387 ( .A1(G902), .A2(n687), .ZN(n483) );
  XNOR2_X1 U388 ( .A(n481), .B(KEYINPUT75), .ZN(n380) );
  NOR2_X1 U389 ( .A1(G953), .A2(G237), .ZN(n516) );
  XNOR2_X1 U390 ( .A(n511), .B(n458), .ZN(n459) );
  XNOR2_X1 U391 ( .A(G116), .B(G113), .ZN(n406) );
  XNOR2_X1 U392 ( .A(n440), .B(G101), .ZN(n407) );
  XNOR2_X1 U393 ( .A(KEYINPUT3), .B(G119), .ZN(n440) );
  XOR2_X1 U394 ( .A(G146), .B(G125), .Z(n474) );
  NOR2_X1 U395 ( .A1(n675), .A2(n604), .ZN(n445) );
  NOR2_X1 U396 ( .A1(n562), .A2(n454), .ZN(n456) );
  XNOR2_X1 U397 ( .A(n379), .B(n378), .ZN(n484) );
  INV_X1 U398 ( .A(KEYINPUT20), .ZN(n378) );
  NOR2_X1 U399 ( .A1(n604), .A2(n479), .ZN(n379) );
  XOR2_X1 U400 ( .A(KEYINPUT5), .B(KEYINPUT91), .Z(n488) );
  NAND2_X1 U401 ( .A1(n412), .A2(n411), .ZN(n410) );
  INV_X1 U402 ( .A(KEYINPUT104), .ZN(n431) );
  NOR2_X1 U403 ( .A1(n706), .A2(n409), .ZN(n408) );
  INV_X1 U404 ( .A(n604), .ZN(n409) );
  NAND2_X1 U405 ( .A1(n565), .A2(KEYINPUT82), .ZN(n426) );
  INV_X1 U406 ( .A(KEYINPUT33), .ZN(n527) );
  OR2_X1 U407 ( .A1(n611), .A2(G902), .ZN(n494) );
  XNOR2_X1 U408 ( .A(n518), .B(n517), .ZN(n680) );
  XNOR2_X1 U409 ( .A(n383), .B(n514), .ZN(n518) );
  XNOR2_X1 U410 ( .A(n515), .B(n350), .ZN(n383) );
  XNOR2_X1 U411 ( .A(n492), .B(n465), .ZN(n678) );
  XNOR2_X1 U412 ( .A(n690), .B(n435), .ZN(n675) );
  XNOR2_X1 U413 ( .A(n394), .B(n436), .ZN(n435) );
  XNOR2_X1 U414 ( .A(n397), .B(n395), .ZN(n394) );
  XNOR2_X1 U415 ( .A(n591), .B(KEYINPUT39), .ZN(n595) );
  INV_X1 U416 ( .A(n582), .ZN(n385) );
  XNOR2_X1 U417 ( .A(n390), .B(n478), .ZN(n687) );
  XNOR2_X1 U418 ( .A(n508), .B(n507), .ZN(n683) );
  INV_X1 U419 ( .A(KEYINPUT95), .ZN(n416) );
  INV_X1 U420 ( .A(KEYINPUT70), .ZN(n401) );
  NOR2_X1 U421 ( .A1(n724), .A2(n725), .ZN(n377) );
  NOR2_X1 U422 ( .A1(n343), .A2(n416), .ZN(n411) );
  NAND2_X1 U423 ( .A1(G234), .A2(G237), .ZN(n449) );
  XOR2_X1 U424 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n450) );
  INV_X1 U425 ( .A(KEYINPUT15), .ZN(n442) );
  XNOR2_X1 U426 ( .A(G902), .B(KEYINPUT86), .ZN(n443) );
  XNOR2_X1 U427 ( .A(n486), .B(n485), .ZN(n557) );
  INV_X1 U428 ( .A(KEYINPUT48), .ZN(n434) );
  XNOR2_X1 U429 ( .A(G143), .B(G113), .ZN(n437) );
  XOR2_X1 U430 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n513) );
  XNOR2_X1 U431 ( .A(G104), .B(G122), .ZN(n512) );
  XNOR2_X1 U432 ( .A(G101), .B(KEYINPUT76), .ZN(n460) );
  XNOR2_X1 U433 ( .A(KEYINPUT18), .B(KEYINPUT87), .ZN(n396) );
  OR2_X1 U434 ( .A1(G237), .A2(G902), .ZN(n446) );
  XNOR2_X1 U435 ( .A(n558), .B(KEYINPUT1), .ZN(n651) );
  XNOR2_X1 U436 ( .A(n388), .B(n387), .ZN(n526) );
  INV_X1 U437 ( .A(KEYINPUT73), .ZN(n387) );
  NAND2_X1 U438 ( .A1(n345), .A2(n648), .ZN(n360) );
  OR2_X1 U439 ( .A1(n680), .A2(G902), .ZN(n438) );
  XNOR2_X1 U440 ( .A(n492), .B(n491), .ZN(n611) );
  INV_X1 U441 ( .A(G227), .ZN(n709) );
  XNOR2_X1 U442 ( .A(n464), .B(n349), .ZN(n405) );
  INV_X1 U443 ( .A(KEYINPUT45), .ZN(n428) );
  XNOR2_X1 U444 ( .A(n469), .B(n468), .ZN(n473) );
  XNOR2_X1 U445 ( .A(G119), .B(G110), .ZN(n468) );
  XOR2_X1 U446 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n469) );
  XNOR2_X1 U447 ( .A(n471), .B(n470), .ZN(n472) );
  INV_X1 U448 ( .A(KEYINPUT23), .ZN(n470) );
  XNOR2_X1 U449 ( .A(G137), .B(G128), .ZN(n471) );
  XNOR2_X1 U450 ( .A(n392), .B(KEYINPUT10), .ZN(n391) );
  INV_X1 U451 ( .A(G140), .ZN(n392) );
  XNOR2_X1 U452 ( .A(G116), .B(G107), .ZN(n499) );
  NAND2_X1 U453 ( .A1(n424), .A2(n423), .ZN(n422) );
  AND2_X1 U454 ( .A1(n427), .A2(n426), .ZN(n425) );
  NOR2_X1 U455 ( .A1(n565), .A2(KEYINPUT82), .ZN(n423) );
  AND2_X1 U456 ( .A1(n626), .A2(n579), .ZN(n368) );
  BUF_X1 U457 ( .A(n571), .Z(n600) );
  AND2_X1 U458 ( .A1(n569), .A2(n375), .ZN(n590) );
  AND2_X1 U459 ( .A1(n568), .A2(n376), .ZN(n375) );
  INV_X1 U460 ( .A(n570), .ZN(n376) );
  XNOR2_X1 U461 ( .A(n510), .B(n509), .ZN(n534) );
  XNOR2_X1 U462 ( .A(KEYINPUT101), .B(G478), .ZN(n509) );
  NOR2_X1 U463 ( .A1(n537), .A2(n385), .ZN(n384) );
  XNOR2_X1 U464 ( .A(n418), .B(n417), .ZN(n720) );
  NOR2_X1 U465 ( .A1(n550), .A2(n577), .ZN(n419) );
  XNOR2_X1 U466 ( .A(n688), .B(n687), .ZN(n356) );
  XNOR2_X1 U467 ( .A(n685), .B(n684), .ZN(n357) );
  INV_X1 U468 ( .A(KEYINPUT60), .ZN(n366) );
  INV_X1 U469 ( .A(KEYINPUT120), .ZN(n361) );
  INV_X1 U470 ( .A(KEYINPUT56), .ZN(n364) );
  NOR2_X1 U471 ( .A1(n544), .A2(n543), .ZN(n343) );
  XOR2_X1 U472 ( .A(n493), .B(G472), .Z(n344) );
  AND2_X1 U473 ( .A1(n374), .A2(n579), .ZN(n345) );
  XOR2_X1 U474 ( .A(n520), .B(n519), .Z(n346) );
  OR2_X1 U475 ( .A1(n637), .A2(n645), .ZN(n347) );
  XOR2_X1 U476 ( .A(n377), .B(n593), .Z(n348) );
  XOR2_X1 U477 ( .A(KEYINPUT16), .B(G122), .Z(n349) );
  AND2_X1 U478 ( .A1(G214), .A2(n516), .ZN(n350) );
  XOR2_X1 U479 ( .A(n675), .B(n674), .Z(n351) );
  XOR2_X1 U480 ( .A(n678), .B(n677), .Z(n352) );
  XOR2_X1 U481 ( .A(n611), .B(n610), .Z(n353) );
  XNOR2_X1 U482 ( .A(n680), .B(KEYINPUT59), .ZN(n354) );
  INV_X1 U483 ( .A(n689), .ZN(n372) );
  XNOR2_X1 U484 ( .A(n614), .B(KEYINPUT83), .ZN(n355) );
  NAND2_X1 U485 ( .A1(n594), .A2(n348), .ZN(n381) );
  XNOR2_X1 U486 ( .A(n381), .B(n434), .ZN(n433) );
  INV_X1 U487 ( .A(n576), .ZN(n374) );
  NOR2_X1 U488 ( .A1(n356), .A2(n689), .ZN(G66) );
  NOR2_X1 U489 ( .A1(n357), .A2(n689), .ZN(G63) );
  NAND2_X1 U490 ( .A1(n358), .A2(n408), .ZN(n389) );
  INV_X1 U491 ( .A(n694), .ZN(n358) );
  XNOR2_X2 U492 ( .A(n429), .B(n428), .ZN(n694) );
  XNOR2_X1 U493 ( .A(n360), .B(n359), .ZN(n560) );
  INV_X1 U494 ( .A(KEYINPUT28), .ZN(n359) );
  XNOR2_X1 U495 ( .A(n362), .B(n361), .ZN(G54) );
  NAND2_X1 U496 ( .A1(n371), .A2(n372), .ZN(n362) );
  XNOR2_X1 U497 ( .A(n363), .B(n355), .ZN(G57) );
  NAND2_X1 U498 ( .A1(n369), .A2(n372), .ZN(n363) );
  XNOR2_X1 U499 ( .A(n365), .B(n364), .ZN(G51) );
  NAND2_X1 U500 ( .A1(n370), .A2(n372), .ZN(n365) );
  XNOR2_X1 U501 ( .A(n367), .B(n366), .ZN(G60) );
  NAND2_X1 U502 ( .A1(n373), .A2(n372), .ZN(n367) );
  NAND2_X1 U503 ( .A1(n433), .A2(n603), .ZN(n706) );
  NAND2_X1 U504 ( .A1(n526), .A2(n577), .ZN(n528) );
  XNOR2_X1 U505 ( .A(n473), .B(n472), .ZN(n475) );
  XNOR2_X1 U506 ( .A(n475), .B(n517), .ZN(n390) );
  NAND2_X1 U507 ( .A1(n578), .A2(n368), .ZN(n598) );
  XNOR2_X1 U508 ( .A(n612), .B(n353), .ZN(n369) );
  XNOR2_X1 U509 ( .A(n676), .B(n351), .ZN(n370) );
  XNOR2_X1 U510 ( .A(n679), .B(n352), .ZN(n371) );
  XNOR2_X1 U511 ( .A(n681), .B(n354), .ZN(n373) );
  AND2_X1 U512 ( .A1(n648), .A2(n633), .ZN(n567) );
  XNOR2_X2 U513 ( .A(n607), .B(KEYINPUT65), .ZN(n609) );
  XNOR2_X1 U514 ( .A(n585), .B(KEYINPUT69), .ZN(n594) );
  NAND2_X1 U515 ( .A1(n382), .A2(n722), .ZN(n585) );
  XNOR2_X1 U516 ( .A(n402), .B(n401), .ZN(n382) );
  NOR2_X1 U517 ( .A1(n564), .A2(KEYINPUT47), .ZN(n563) );
  NAND2_X1 U518 ( .A1(n621), .A2(n638), .ZN(n564) );
  NAND2_X1 U519 ( .A1(n386), .A2(n384), .ZN(n540) );
  INV_X1 U520 ( .A(n538), .ZN(n386) );
  NAND2_X1 U521 ( .A1(n389), .A2(n606), .ZN(n607) );
  NAND2_X1 U522 ( .A1(n484), .A2(G217), .ZN(n480) );
  NAND2_X1 U523 ( .A1(n576), .A2(n557), .ZN(n650) );
  XNOR2_X2 U524 ( .A(n467), .B(n466), .ZN(n558) );
  INV_X1 U525 ( .A(n708), .ZN(n552) );
  XNOR2_X1 U526 ( .A(n439), .B(n396), .ZN(n395) );
  NOR2_X1 U527 ( .A1(n708), .A2(n398), .ZN(n397) );
  INV_X1 U528 ( .A(G224), .ZN(n398) );
  XNOR2_X2 U529 ( .A(n399), .B(G131), .ZN(n511) );
  XNOR2_X1 U530 ( .A(n400), .B(n505), .ZN(n508) );
  XNOR2_X2 U531 ( .A(n457), .B(G134), .ZN(n400) );
  NAND2_X1 U532 ( .A1(n404), .A2(n403), .ZN(n402) );
  XNOR2_X1 U533 ( .A(n575), .B(KEYINPUT79), .ZN(n403) );
  XNOR2_X1 U534 ( .A(n563), .B(KEYINPUT71), .ZN(n404) );
  NOR2_X1 U535 ( .A1(n694), .A2(n706), .ZN(n631) );
  NAND2_X1 U536 ( .A1(n413), .A2(n410), .ZN(n421) );
  INV_X1 U537 ( .A(n545), .ZN(n412) );
  AND2_X1 U538 ( .A1(n415), .A2(n414), .ZN(n413) );
  NAND2_X1 U539 ( .A1(n545), .A2(n416), .ZN(n415) );
  NAND2_X1 U540 ( .A1(n420), .A2(n720), .ZN(n551) );
  INV_X1 U541 ( .A(KEYINPUT103), .ZN(n417) );
  NAND2_X1 U542 ( .A1(n549), .A2(n419), .ZN(n418) );
  NAND2_X1 U543 ( .A1(n421), .A2(n638), .ZN(n420) );
  XNOR2_X2 U544 ( .A(n456), .B(n455), .ZN(n544) );
  OR2_X2 U545 ( .A1(n678), .A2(G902), .ZN(n467) );
  NOR2_X2 U546 ( .A1(n588), .A2(n562), .ZN(n621) );
  XNOR2_X2 U547 ( .A(n580), .B(n448), .ZN(n562) );
  NAND2_X2 U548 ( .A1(n425), .A2(n422), .ZN(n580) );
  INV_X1 U549 ( .A(n571), .ZN(n424) );
  NAND2_X1 U550 ( .A1(n571), .A2(KEYINPUT82), .ZN(n427) );
  NAND2_X1 U551 ( .A1(n432), .A2(n430), .ZN(n429) );
  XNOR2_X1 U552 ( .A(n551), .B(n431), .ZN(n430) );
  XNOR2_X1 U553 ( .A(n542), .B(KEYINPUT44), .ZN(n432) );
  XNOR2_X1 U554 ( .A(n457), .B(n474), .ZN(n436) );
  XNOR2_X1 U555 ( .A(n511), .B(n437), .ZN(n515) );
  INV_X1 U556 ( .A(n533), .ZN(n524) );
  BUF_X1 U557 ( .A(n682), .Z(n686) );
  NOR2_X1 U558 ( .A1(n580), .A2(n598), .ZN(n581) );
  AND2_X1 U559 ( .A1(n577), .A2(n644), .ZN(n578) );
  AND2_X1 U560 ( .A1(n708), .A2(n613), .ZN(n689) );
  XNOR2_X2 U561 ( .A(G143), .B(G128), .ZN(n457) );
  XNOR2_X2 U562 ( .A(KEYINPUT64), .B(G953), .ZN(n708) );
  XNOR2_X1 U563 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n439) );
  AND2_X1 U564 ( .A1(G210), .A2(n446), .ZN(n444) );
  NAND2_X1 U565 ( .A1(n446), .A2(G214), .ZN(n447) );
  XNOR2_X1 U566 ( .A(KEYINPUT88), .B(n447), .ZN(n633) );
  INV_X1 U567 ( .A(n633), .ZN(n565) );
  INV_X1 U568 ( .A(KEYINPUT19), .ZN(n448) );
  XOR2_X1 U569 ( .A(n450), .B(n449), .Z(n451) );
  NAND2_X1 U570 ( .A1(G952), .A2(n451), .ZN(n663) );
  NOR2_X1 U571 ( .A1(G953), .A2(n663), .ZN(n555) );
  NAND2_X1 U572 ( .A1(n451), .A2(G902), .ZN(n553) );
  INV_X1 U573 ( .A(G898), .ZN(n697) );
  NAND2_X1 U574 ( .A1(G953), .A2(n697), .ZN(n691) );
  NOR2_X1 U575 ( .A1(n553), .A2(n691), .ZN(n452) );
  NOR2_X1 U576 ( .A1(n555), .A2(n452), .ZN(n453) );
  XOR2_X1 U577 ( .A(KEYINPUT89), .B(n453), .Z(n454) );
  INV_X1 U578 ( .A(KEYINPUT0), .ZN(n455) );
  XNOR2_X1 U579 ( .A(KEYINPUT4), .B(G137), .ZN(n458) );
  OR2_X1 U580 ( .A1(n708), .A2(n709), .ZN(n462) );
  XNOR2_X1 U581 ( .A(n460), .B(G140), .ZN(n461) );
  XNOR2_X1 U582 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U583 ( .A(n464), .B(n463), .ZN(n465) );
  INV_X1 U584 ( .A(G469), .ZN(n466) );
  XOR2_X1 U585 ( .A(KEYINPUT80), .B(KEYINPUT8), .Z(n477) );
  NAND2_X1 U586 ( .A1(G234), .A2(n552), .ZN(n476) );
  XNOR2_X1 U587 ( .A(n477), .B(n476), .ZN(n506) );
  NAND2_X1 U588 ( .A1(G221), .A2(n506), .ZN(n478) );
  XOR2_X1 U589 ( .A(KEYINPUT74), .B(KEYINPUT25), .Z(n481) );
  INV_X1 U590 ( .A(G234), .ZN(n479) );
  NAND2_X1 U591 ( .A1(n484), .A2(G221), .ZN(n486) );
  INV_X1 U592 ( .A(KEYINPUT21), .ZN(n485) );
  NAND2_X1 U593 ( .A1(n516), .A2(G210), .ZN(n487) );
  XOR2_X1 U594 ( .A(n488), .B(n487), .Z(n489) );
  XNOR2_X1 U595 ( .A(n490), .B(n489), .ZN(n491) );
  INV_X1 U596 ( .A(KEYINPUT92), .ZN(n493) );
  XNOR2_X2 U597 ( .A(n494), .B(n344), .ZN(n648) );
  NAND2_X1 U598 ( .A1(n526), .A2(n648), .ZN(n496) );
  INV_X1 U599 ( .A(KEYINPUT93), .ZN(n495) );
  XNOR2_X1 U600 ( .A(n496), .B(n495), .ZN(n656) );
  XNOR2_X1 U601 ( .A(KEYINPUT94), .B(KEYINPUT31), .ZN(n497) );
  XNOR2_X2 U602 ( .A(n498), .B(n497), .ZN(n545) );
  XOR2_X1 U603 ( .A(KEYINPUT7), .B(KEYINPUT99), .Z(n500) );
  XNOR2_X1 U604 ( .A(n500), .B(n499), .ZN(n504) );
  XOR2_X1 U605 ( .A(KEYINPUT98), .B(KEYINPUT9), .Z(n502) );
  XNOR2_X1 U606 ( .A(G122), .B(KEYINPUT100), .ZN(n501) );
  XNOR2_X1 U607 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U608 ( .A(n504), .B(n503), .Z(n505) );
  NAND2_X1 U609 ( .A1(G217), .A2(n506), .ZN(n507) );
  NOR2_X1 U610 ( .A1(n683), .A2(G902), .ZN(n510) );
  XNOR2_X1 U611 ( .A(n513), .B(n512), .ZN(n514) );
  INV_X1 U612 ( .A(n517), .ZN(n704) );
  XOR2_X1 U613 ( .A(KEYINPUT13), .B(KEYINPUT96), .Z(n520) );
  XNOR2_X1 U614 ( .A(KEYINPUT97), .B(G475), .ZN(n519) );
  AND2_X1 U615 ( .A1(n534), .A2(n524), .ZN(n622) );
  NAND2_X1 U616 ( .A1(n545), .A2(n622), .ZN(n522) );
  XOR2_X1 U617 ( .A(G116), .B(KEYINPUT113), .Z(n521) );
  XNOR2_X1 U618 ( .A(n522), .B(n521), .ZN(G18) );
  NOR2_X1 U619 ( .A1(n534), .A2(n524), .ZN(n626) );
  NAND2_X1 U620 ( .A1(n545), .A2(n626), .ZN(n523) );
  XNOR2_X1 U621 ( .A(n523), .B(G113), .ZN(G15) );
  NAND2_X1 U622 ( .A1(n533), .A2(n534), .ZN(n525) );
  XOR2_X1 U623 ( .A(KEYINPUT105), .B(n525), .Z(n572) );
  INV_X1 U624 ( .A(n648), .ZN(n566) );
  XNOR2_X1 U625 ( .A(n566), .B(KEYINPUT6), .ZN(n577) );
  XNOR2_X2 U626 ( .A(n528), .B(n527), .ZN(n632) );
  NOR2_X1 U627 ( .A1(n632), .A2(n544), .ZN(n530) );
  XNOR2_X1 U628 ( .A(KEYINPUT34), .B(KEYINPUT77), .ZN(n529) );
  XNOR2_X1 U629 ( .A(n530), .B(n529), .ZN(n531) );
  NOR2_X1 U630 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U631 ( .A(KEYINPUT102), .B(n535), .Z(n637) );
  INV_X1 U632 ( .A(n576), .ZN(n644) );
  NAND2_X1 U633 ( .A1(n549), .A2(n644), .ZN(n538) );
  NAND2_X1 U634 ( .A1(n385), .A2(n566), .ZN(n536) );
  OR2_X1 U635 ( .A1(n538), .A2(n536), .ZN(n620) );
  NAND2_X1 U636 ( .A1(n717), .A2(n620), .ZN(n541) );
  INV_X1 U637 ( .A(n577), .ZN(n548) );
  XOR2_X1 U638 ( .A(KEYINPUT78), .B(n548), .Z(n537) );
  INV_X1 U639 ( .A(n651), .ZN(n582) );
  XOR2_X1 U640 ( .A(KEYINPUT66), .B(KEYINPUT32), .Z(n539) );
  NOR2_X1 U641 ( .A1(n650), .A2(n558), .ZN(n568) );
  NAND2_X1 U642 ( .A1(n568), .A2(n566), .ZN(n543) );
  INV_X1 U643 ( .A(n626), .ZN(n547) );
  INV_X1 U644 ( .A(n622), .ZN(n546) );
  NAND2_X1 U645 ( .A1(n547), .A2(n546), .ZN(n638) );
  OR2_X1 U646 ( .A1(n582), .A2(n644), .ZN(n550) );
  OR2_X1 U647 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U648 ( .A1(G900), .A2(n554), .ZN(n556) );
  NOR2_X1 U649 ( .A1(n556), .A2(n555), .ZN(n570) );
  INV_X1 U650 ( .A(n557), .ZN(n645) );
  NOR2_X1 U651 ( .A1(n570), .A2(n645), .ZN(n579) );
  INV_X1 U652 ( .A(n558), .ZN(n559) );
  NAND2_X1 U653 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U654 ( .A(n561), .B(KEYINPUT106), .ZN(n588) );
  NAND2_X1 U655 ( .A1(n564), .A2(KEYINPUT47), .ZN(n574) );
  XNOR2_X1 U656 ( .A(KEYINPUT30), .B(n567), .ZN(n569) );
  NOR2_X1 U657 ( .A1(n600), .A2(n572), .ZN(n573) );
  NAND2_X1 U658 ( .A1(n590), .A2(n573), .ZN(n625) );
  NAND2_X1 U659 ( .A1(n574), .A2(n625), .ZN(n575) );
  XNOR2_X1 U660 ( .A(KEYINPUT36), .B(n581), .ZN(n583) );
  NAND2_X1 U661 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U662 ( .A(n584), .B(KEYINPUT108), .ZN(n722) );
  XNOR2_X1 U663 ( .A(KEYINPUT38), .B(n600), .ZN(n634) );
  NAND2_X1 U664 ( .A1(n634), .A2(n633), .ZN(n639) );
  NOR2_X1 U665 ( .A1(n637), .A2(n639), .ZN(n587) );
  XOR2_X1 U666 ( .A(KEYINPUT41), .B(KEYINPUT107), .Z(n586) );
  XNOR2_X1 U667 ( .A(n587), .B(n586), .ZN(n664) );
  NOR2_X1 U668 ( .A1(n664), .A2(n588), .ZN(n589) );
  XNOR2_X1 U669 ( .A(n589), .B(KEYINPUT42), .ZN(n725) );
  NAND2_X1 U670 ( .A1(n590), .A2(n634), .ZN(n591) );
  NAND2_X1 U671 ( .A1(n626), .A2(n595), .ZN(n592) );
  XOR2_X1 U672 ( .A(KEYINPUT40), .B(n592), .Z(n724) );
  XNOR2_X1 U673 ( .A(KEYINPUT46), .B(KEYINPUT81), .ZN(n593) );
  NAND2_X1 U674 ( .A1(n595), .A2(n622), .ZN(n596) );
  XNOR2_X1 U675 ( .A(n596), .B(KEYINPUT109), .ZN(n718) );
  NAND2_X1 U676 ( .A1(n385), .A2(n633), .ZN(n597) );
  OR2_X1 U677 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U678 ( .A(n599), .B(KEYINPUT43), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n601), .A2(n600), .ZN(n629) );
  INV_X1 U680 ( .A(n629), .ZN(n602) );
  NOR2_X1 U681 ( .A1(n718), .A2(n602), .ZN(n603) );
  NAND2_X1 U682 ( .A1(n604), .A2(KEYINPUT2), .ZN(n605) );
  XOR2_X1 U683 ( .A(KEYINPUT67), .B(n605), .Z(n606) );
  AND2_X1 U684 ( .A1(n631), .A2(KEYINPUT2), .ZN(n608) );
  NOR2_X4 U685 ( .A1(n609), .A2(n608), .ZN(n682) );
  NAND2_X1 U686 ( .A1(n682), .A2(G472), .ZN(n612) );
  XNOR2_X1 U687 ( .A(KEYINPUT84), .B(KEYINPUT62), .ZN(n610) );
  INV_X1 U688 ( .A(G952), .ZN(n613) );
  XNOR2_X1 U689 ( .A(KEYINPUT85), .B(KEYINPUT63), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n343), .A2(n626), .ZN(n615) );
  XNOR2_X1 U691 ( .A(n615), .B(G104), .ZN(G6) );
  XOR2_X1 U692 ( .A(KEYINPUT26), .B(KEYINPUT111), .Z(n617) );
  NAND2_X1 U693 ( .A1(n343), .A2(n622), .ZN(n616) );
  XNOR2_X1 U694 ( .A(n617), .B(n616), .ZN(n619) );
  XOR2_X1 U695 ( .A(G107), .B(KEYINPUT27), .Z(n618) );
  XNOR2_X1 U696 ( .A(n619), .B(n618), .ZN(G9) );
  XNOR2_X1 U697 ( .A(G110), .B(n620), .ZN(G12) );
  XOR2_X1 U698 ( .A(G128), .B(KEYINPUT29), .Z(n624) );
  NAND2_X1 U699 ( .A1(n621), .A2(n622), .ZN(n623) );
  XNOR2_X1 U700 ( .A(n624), .B(n623), .ZN(G30) );
  XNOR2_X1 U701 ( .A(G143), .B(n625), .ZN(G45) );
  NAND2_X1 U702 ( .A1(n621), .A2(n626), .ZN(n627) );
  XNOR2_X1 U703 ( .A(n627), .B(KEYINPUT112), .ZN(n628) );
  XNOR2_X1 U704 ( .A(G146), .B(n628), .ZN(G48) );
  XNOR2_X1 U705 ( .A(G140), .B(KEYINPUT114), .ZN(n630) );
  XNOR2_X1 U706 ( .A(n630), .B(n629), .ZN(G42) );
  XNOR2_X1 U707 ( .A(n631), .B(KEYINPUT2), .ZN(n668) );
  NOR2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U709 ( .A(n635), .B(KEYINPUT116), .ZN(n636) );
  NOR2_X1 U710 ( .A1(n637), .A2(n636), .ZN(n642) );
  INV_X1 U711 ( .A(n638), .ZN(n640) );
  NOR2_X1 U712 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U713 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U714 ( .A1(n632), .A2(n643), .ZN(n660) );
  XOR2_X1 U715 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n647) );
  NAND2_X1 U716 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U717 ( .A(n647), .B(n646), .ZN(n649) );
  NOR2_X1 U718 ( .A1(n649), .A2(n648), .ZN(n654) );
  NAND2_X1 U719 ( .A1(n385), .A2(n650), .ZN(n652) );
  XNOR2_X1 U720 ( .A(n652), .B(KEYINPUT50), .ZN(n653) );
  NAND2_X1 U721 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U722 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U723 ( .A(n657), .B(KEYINPUT51), .ZN(n658) );
  NOR2_X1 U724 ( .A1(n658), .A2(n664), .ZN(n659) );
  NOR2_X1 U725 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U726 ( .A(n661), .B(KEYINPUT52), .ZN(n662) );
  NOR2_X1 U727 ( .A1(n663), .A2(n662), .ZN(n666) );
  NOR2_X1 U728 ( .A1(n632), .A2(n664), .ZN(n665) );
  NOR2_X1 U729 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U730 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U731 ( .A(KEYINPUT117), .B(n669), .Z(n670) );
  XOR2_X1 U732 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n671) );
  XNOR2_X1 U733 ( .A(KEYINPUT118), .B(n671), .ZN(n672) );
  XNOR2_X1 U734 ( .A(n673), .B(n672), .ZN(G75) );
  NAND2_X1 U735 ( .A1(n682), .A2(G210), .ZN(n676) );
  XOR2_X1 U736 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n674) );
  NAND2_X1 U737 ( .A1(n682), .A2(G469), .ZN(n679) );
  XOR2_X1 U738 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n677) );
  NAND2_X1 U739 ( .A1(n682), .A2(G475), .ZN(n681) );
  NAND2_X1 U740 ( .A1(n686), .A2(G478), .ZN(n685) );
  XOR2_X1 U741 ( .A(KEYINPUT121), .B(n683), .Z(n684) );
  NAND2_X1 U742 ( .A1(n686), .A2(G217), .ZN(n688) );
  XNOR2_X1 U743 ( .A(n690), .B(KEYINPUT124), .ZN(n692) );
  NAND2_X1 U744 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U745 ( .A(n693), .B(KEYINPUT125), .ZN(n703) );
  OR2_X1 U746 ( .A1(n694), .A2(G953), .ZN(n701) );
  XOR2_X1 U747 ( .A(KEYINPUT122), .B(KEYINPUT61), .Z(n696) );
  NAND2_X1 U748 ( .A1(G224), .A2(G953), .ZN(n695) );
  XNOR2_X1 U749 ( .A(n696), .B(n695), .ZN(n698) );
  NOR2_X1 U750 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U751 ( .A(n699), .B(KEYINPUT123), .ZN(n700) );
  NAND2_X1 U752 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U753 ( .A(n703), .B(n702), .ZN(G69) );
  XNOR2_X1 U754 ( .A(n705), .B(n704), .ZN(n710) );
  XNOR2_X1 U755 ( .A(n706), .B(n710), .ZN(n707) );
  NOR2_X1 U756 ( .A1(n708), .A2(n707), .ZN(n715) );
  XNOR2_X1 U757 ( .A(n710), .B(n709), .ZN(n711) );
  NAND2_X1 U758 ( .A1(n711), .A2(G900), .ZN(n712) );
  NAND2_X1 U759 ( .A1(G953), .A2(n712), .ZN(n713) );
  XOR2_X1 U760 ( .A(KEYINPUT126), .B(n713), .Z(n714) );
  NOR2_X1 U761 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U762 ( .A(KEYINPUT127), .B(n716), .ZN(G72) );
  XNOR2_X1 U763 ( .A(n717), .B(G122), .ZN(G24) );
  XOR2_X1 U764 ( .A(G134), .B(n718), .Z(G36) );
  XOR2_X1 U765 ( .A(G119), .B(n719), .Z(G21) );
  XNOR2_X1 U766 ( .A(G101), .B(KEYINPUT110), .ZN(n721) );
  XNOR2_X1 U767 ( .A(n721), .B(n720), .ZN(G3) );
  XOR2_X1 U768 ( .A(n722), .B(G125), .Z(n723) );
  XNOR2_X1 U769 ( .A(KEYINPUT37), .B(n723), .ZN(G27) );
  XOR2_X1 U770 ( .A(G131), .B(n724), .Z(G33) );
  XOR2_X1 U771 ( .A(G137), .B(n725), .Z(G39) );
endmodule

