//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n789, new_n790, new_n792, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT76), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT76), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n207), .A2(G155gat), .A3(G162gat), .ZN(new_n208));
  INV_X1    g007(.A(G155gat), .ZN(new_n209));
  INV_X1    g008(.A(G162gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n206), .A2(new_n208), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G148gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G141gat), .ZN(new_n214));
  INV_X1    g013(.A(G141gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n207), .A2(KEYINPUT2), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n212), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT77), .B1(new_n215), .B2(G148gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT77), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(new_n213), .A3(G141gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n223), .A3(new_n216), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n205), .B1(new_n211), .B2(KEYINPUT2), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n220), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT3), .ZN(new_n228));
  XNOR2_X1  g027(.A(G197gat), .B(G204gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(G211gat), .A2(G218gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT72), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT22), .ZN(new_n232));
  AND3_X1   g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n231), .B1(new_n230), .B2(new_n232), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n229), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  XOR2_X1   g034(.A(G211gat), .B(G218gat), .Z(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n235), .B(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT29), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n206), .A2(new_n208), .A3(new_n211), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n240), .B1(new_n217), .B2(new_n218), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n224), .A2(new_n225), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n239), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n228), .B1(new_n238), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT82), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n228), .B(KEYINPUT82), .C1(new_n238), .C2(new_n243), .ZN(new_n247));
  INV_X1    g046(.A(G228gat), .ZN(new_n248));
  INV_X1    g047(.A(G233gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n212), .A2(new_n219), .B1(new_n224), .B2(new_n225), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT78), .B(KEYINPUT3), .Z(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n239), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(new_n238), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n246), .A2(new_n247), .A3(new_n250), .A4(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n250), .ZN(new_n257));
  INV_X1    g056(.A(new_n255), .ZN(new_n258));
  OAI22_X1  g057(.A1(new_n238), .A2(new_n243), .B1(new_n251), .B2(new_n252), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G22gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n256), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT83), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n261), .B1(new_n256), .B2(new_n260), .ZN(new_n265));
  NOR3_X1   g064(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n256), .A2(new_n260), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G22gat), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT83), .B1(new_n268), .B2(new_n262), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n204), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n264), .B1(new_n263), .B2(new_n265), .ZN(new_n271));
  INV_X1    g070(.A(new_n204), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n275));
  XNOR2_X1  g074(.A(G127gat), .B(G134gat), .ZN(new_n276));
  INV_X1    g075(.A(G120gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G113gat), .ZN(new_n278));
  INV_X1    g077(.A(G113gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G120gat), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT1), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n276), .B1(new_n281), .B2(KEYINPUT69), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(KEYINPUT69), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n284));
  XNOR2_X1  g083(.A(G113gat), .B(G120gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n284), .B1(new_n285), .B2(KEYINPUT1), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n282), .B1(new_n287), .B2(new_n276), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT25), .ZN(new_n289));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT23), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n290), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n292), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT66), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT65), .B(KEYINPUT23), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(KEYINPUT66), .A3(new_n292), .ZN(new_n302));
  AOI211_X1 g101(.A(new_n289), .B(new_n294), .C1(new_n300), .C2(new_n302), .ZN(new_n303));
  XOR2_X1   g102(.A(KEYINPUT67), .B(G183gat), .Z(new_n304));
  INV_X1    g103(.A(KEYINPUT68), .ZN(new_n305));
  INV_X1    g104(.A(G190gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT67), .B(G183gat), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT68), .B1(new_n308), .B2(G190gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT24), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n307), .A2(new_n309), .A3(new_n310), .A4(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n294), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT64), .ZN(new_n316));
  OR2_X1    g115(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n310), .A2(new_n316), .ZN(new_n318));
  INV_X1    g117(.A(G183gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(new_n306), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n317), .A2(new_n318), .A3(new_n320), .A4(new_n313), .ZN(new_n321));
  INV_X1    g120(.A(new_n302), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT66), .B1(new_n301), .B2(new_n292), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n315), .B(new_n321), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n303), .A2(new_n314), .B1(new_n324), .B2(new_n289), .ZN(new_n325));
  NOR2_X1   g124(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n328));
  AOI21_X1  g127(.A(G190gat), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT28), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n292), .A2(KEYINPUT26), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(new_n290), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n292), .A2(KEYINPUT26), .ZN(new_n333));
  OAI221_X1 g132(.A(new_n311), .B1(new_n329), .B2(new_n330), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n326), .B1(new_n308), .B2(KEYINPUT27), .ZN(new_n335));
  NOR3_X1   g134(.A1(new_n335), .A2(KEYINPUT28), .A3(G190gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n288), .B1(new_n325), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n324), .A2(new_n289), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n294), .B1(new_n300), .B2(new_n302), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n314), .A2(new_n340), .A3(KEYINPUT25), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n337), .ZN(new_n343));
  INV_X1    g142(.A(new_n288), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n338), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G227gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n347), .A2(new_n249), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT34), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT34), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n346), .A2(new_n352), .A3(new_n349), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n345), .A3(new_n348), .ZN(new_n355));
  XOR2_X1   g154(.A(G15gat), .B(G43gat), .Z(new_n356));
  XNOR2_X1  g155(.A(G71gat), .B(G99gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT33), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n355), .A2(KEYINPUT32), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT70), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT70), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n355), .A2(new_n362), .A3(KEYINPUT32), .A4(new_n359), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n355), .A2(KEYINPUT32), .ZN(new_n365));
  INV_X1    g164(.A(new_n355), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n365), .B(new_n358), .C1(new_n366), .C2(KEYINPUT33), .ZN(new_n367));
  AOI211_X1 g166(.A(new_n275), .B(new_n354), .C1(new_n364), .C2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n351), .A2(new_n353), .A3(KEYINPUT71), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n352), .B1(new_n346), .B2(new_n349), .ZN(new_n370));
  AOI211_X1 g169(.A(KEYINPUT34), .B(new_n348), .C1(new_n338), .C2(new_n345), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n275), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n364), .A2(new_n369), .A3(new_n372), .A4(new_n367), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n274), .B1(new_n368), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT89), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n287), .A2(new_n276), .ZN(new_n378));
  INV_X1    g177(.A(new_n282), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(new_n251), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT4), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT4), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n288), .A2(new_n382), .A3(new_n251), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n378), .A2(new_n379), .B1(new_n251), .B2(new_n252), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n381), .A2(new_n383), .B1(new_n228), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G225gat), .A2(G233gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  XOR2_X1   g186(.A(KEYINPUT79), .B(KEYINPUT5), .Z(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G1gat), .B(G29gat), .ZN(new_n391));
  INV_X1    g190(.A(G85gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT0), .B(G57gat), .ZN(new_n394));
  XOR2_X1   g193(.A(new_n393), .B(new_n394), .Z(new_n395));
  NAND2_X1  g194(.A1(new_n344), .A2(new_n227), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n386), .B1(new_n396), .B2(new_n380), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n397), .B1(new_n385), .B2(new_n386), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n390), .B(new_n395), .C1(new_n389), .C2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT80), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n397), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n388), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n404), .A2(KEYINPUT80), .A3(new_n390), .A4(new_n395), .ZN(new_n405));
  INV_X1    g204(.A(new_n395), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n398), .A2(new_n389), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n388), .B1(new_n385), .B2(new_n386), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT6), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n401), .A2(new_n405), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n399), .A2(new_n410), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(G226gat), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n415), .A2(new_n249), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n239), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n342), .B2(new_n343), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n342), .A2(new_n343), .A3(new_n416), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n238), .A3(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n235), .B(new_n236), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n325), .A2(new_n337), .A3(new_n417), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n423), .B1(new_n424), .B2(new_n419), .ZN(new_n425));
  XNOR2_X1  g224(.A(G8gat), .B(G36gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(G64gat), .B(G92gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n422), .A2(new_n425), .A3(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT74), .B(KEYINPUT30), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n432), .A2(KEYINPUT75), .ZN(new_n433));
  XOR2_X1   g232(.A(new_n428), .B(KEYINPUT73), .Z(new_n434));
  AOI21_X1  g233(.A(new_n238), .B1(new_n420), .B2(new_n421), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n424), .A2(new_n419), .A3(new_n423), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT30), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n437), .B1(new_n438), .B2(new_n430), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT75), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n440), .B1(new_n430), .B2(new_n431), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n433), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n414), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT81), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n414), .A2(new_n442), .A3(KEYINPUT81), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n364), .A2(new_n372), .A3(new_n367), .ZN(new_n447));
  INV_X1    g246(.A(new_n369), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n373), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n450), .A2(KEYINPUT89), .A3(new_n274), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n377), .A2(new_n445), .A3(new_n446), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT35), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT90), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n452), .A2(KEYINPUT90), .A3(KEYINPUT35), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n409), .A2(new_n410), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT85), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n458), .B1(new_n407), .B2(new_n408), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n404), .A2(KEYINPUT85), .A3(new_n390), .ZN(new_n460));
  XOR2_X1   g259(.A(new_n395), .B(KEYINPUT84), .Z(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n459), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n413), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n465), .A2(KEYINPUT88), .A3(new_n442), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT88), .B1(new_n465), .B2(new_n442), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT35), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n450), .A2(new_n468), .A3(new_n274), .ZN(new_n469));
  NOR3_X1   g268(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n471), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n270), .A2(new_n273), .ZN(new_n473));
  INV_X1    g272(.A(new_n442), .ZN(new_n474));
  OR3_X1    g273(.A1(new_n385), .A2(KEYINPUT39), .A3(new_n386), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n461), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT40), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n385), .A2(new_n386), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n396), .A2(new_n386), .A3(new_n380), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT39), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  OR3_X1    g280(.A1(new_n476), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n477), .B1(new_n476), .B2(new_n481), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n463), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n473), .B1(new_n474), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n422), .A2(new_n425), .A3(KEYINPUT86), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n486), .B(KEYINPUT37), .C1(KEYINPUT86), .C2(new_n425), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT38), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT37), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n422), .A2(new_n425), .A3(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n487), .A2(new_n488), .A3(new_n434), .A4(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT87), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n430), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n494), .B1(new_n491), .B2(new_n492), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n490), .A2(new_n428), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n489), .B1(new_n422), .B2(new_n425), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT38), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n493), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n485), .B1(new_n499), .B2(new_n465), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n450), .B(KEYINPUT36), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n274), .B1(new_n445), .B2(new_n446), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n472), .A2(new_n505), .ZN(new_n506));
  OR3_X1    g305(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(G29gat), .ZN(new_n510));
  INV_X1    g309(.A(G36gat), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G50gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(G43gat), .ZN(new_n514));
  INV_X1    g313(.A(G43gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(G50gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT91), .ZN(new_n518));
  XNOR2_X1  g317(.A(G43gat), .B(G50gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT91), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n518), .A2(new_n521), .A3(KEYINPUT15), .ZN(new_n522));
  INV_X1    g321(.A(new_n516), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT15), .B1(new_n523), .B2(KEYINPUT92), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT92), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n512), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n507), .A2(new_n508), .B1(G29gat), .B2(G36gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT15), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n530), .B1(new_n517), .B2(KEYINPUT91), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n529), .B1(new_n531), .B2(new_n521), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT17), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(G15gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n261), .ZN(new_n535));
  INV_X1    g334(.A(G1gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(G15gat), .A2(G22gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n535), .A2(new_n537), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n536), .A2(KEYINPUT16), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(G8gat), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n542), .B1(new_n538), .B2(KEYINPUT93), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n541), .B(new_n543), .Z(new_n544));
  NAND2_X1  g343(.A1(new_n522), .A2(new_n512), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n531), .A2(new_n521), .B1(new_n524), .B2(new_n526), .ZN(new_n547));
  OAI211_X1 g346(.A(new_n545), .B(new_n546), .C1(new_n547), .C2(new_n512), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n544), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n545), .B1(new_n547), .B2(new_n512), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n541), .B(new_n543), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n549), .A2(new_n550), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT18), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n549), .A2(new_n554), .A3(KEYINPUT18), .A4(new_n550), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n544), .A2(new_n551), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT94), .B(KEYINPUT13), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(new_n550), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n557), .A2(new_n558), .A3(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(G197gat), .ZN(new_n567));
  XOR2_X1   g366(.A(KEYINPUT11), .B(G169gat), .Z(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT12), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n557), .A2(new_n558), .A3(new_n564), .A4(new_n570), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n506), .A2(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(G127gat), .B(G155gat), .Z(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G71gat), .A2(G78gat), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT9), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OR2_X1    g381(.A1(G57gat), .A2(G64gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(G57gat), .A2(G64gat), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT95), .ZN(new_n586));
  XNOR2_X1  g385(.A(G71gat), .B(G78gat), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n587), .B1(new_n585), .B2(new_n586), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT21), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n587), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n594));
  AND2_X1   g393(.A1(G57gat), .A2(G64gat), .ZN(new_n595));
  NOR2_X1   g394(.A1(G57gat), .A2(G64gat), .ZN(new_n596));
  NOR3_X1   g395(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n593), .B1(new_n597), .B2(KEYINPUT95), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n600), .A2(KEYINPUT21), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n544), .B1(new_n592), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT96), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(new_n319), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(G211gat), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n553), .B1(KEYINPUT21), .B2(new_n600), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n602), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n606), .B1(new_n602), .B2(new_n607), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n579), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n602), .A2(new_n607), .ZN(new_n611));
  INV_X1    g410(.A(new_n606), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n602), .A2(new_n606), .A3(new_n607), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(new_n578), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G134gat), .B(G162gat), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT41), .ZN(new_n618));
  INV_X1    g417(.A(G232gat), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n618), .B1(new_n619), .B2(new_n249), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n617), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(KEYINPUT97), .B(KEYINPUT98), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G99gat), .A2(G106gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT8), .ZN(new_n626));
  NAND2_X1  g425(.A1(G85gat), .A2(G92gat), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT7), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(G92gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n392), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n626), .A2(new_n629), .A3(new_n631), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G99gat), .B(G106gat), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  AND3_X1   g435(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI22_X1  g438(.A1(KEYINPUT8), .A2(new_n625), .B1(new_n392), .B2(new_n630), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n634), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n533), .B(new_n548), .C1(new_n636), .C2(new_n641), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n618), .A2(new_n619), .A3(new_n249), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n636), .A2(new_n641), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n643), .B1(new_n552), .B2(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(G190gat), .B(G218gat), .Z(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n642), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n647), .B1(new_n642), .B2(new_n645), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n624), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n650), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n652), .A2(new_n623), .A3(new_n648), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n616), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT99), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n639), .A2(new_n634), .A3(new_n640), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n633), .A2(new_n635), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n660), .B(new_n661), .C1(new_n588), .C2(new_n589), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT10), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n659), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n598), .B(new_n599), .C1(new_n636), .C2(new_n641), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n662), .A2(new_n665), .A3(new_n663), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n644), .A2(new_n600), .A3(KEYINPUT99), .A4(KEYINPUT10), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(G230gat), .A2(G233gat), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(KEYINPUT100), .Z(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n662), .A2(new_n665), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n670), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n658), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n672), .A2(new_n674), .A3(new_n658), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n654), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n575), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n414), .A2(KEYINPUT101), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n414), .A2(KEYINPUT101), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(G1gat), .ZN(G1324gat));
  INV_X1    g486(.A(KEYINPUT42), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n506), .A2(new_n574), .A3(new_n474), .A4(new_n679), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT102), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n470), .B1(new_n453), .B2(new_n454), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n504), .B1(new_n691), .B2(new_n456), .ZN(new_n692));
  INV_X1    g491(.A(new_n574), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n694), .A2(new_n695), .A3(new_n474), .A4(new_n679), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n690), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT16), .B(G8gat), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n688), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n689), .A2(new_n688), .A3(new_n698), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n697), .B2(G8gat), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n699), .A2(new_n701), .A3(KEYINPUT103), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(G1325gat));
  AOI21_X1  g505(.A(G15gat), .B1(new_n681), .B2(new_n450), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n501), .A2(new_n534), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(new_n681), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1326gat));
  NAND2_X1  g510(.A1(new_n681), .A2(new_n473), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT105), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT43), .B(G22gat), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n712), .B(KEYINPUT105), .ZN(new_n717));
  INV_X1    g516(.A(new_n715), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n716), .A2(new_n719), .ZN(G1327gat));
  NOR2_X1   g519(.A1(new_n678), .A2(new_n616), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n653), .A2(new_n651), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT106), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n575), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n725), .A2(new_n510), .A3(new_n685), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT45), .ZN(new_n727));
  INV_X1    g526(.A(new_n573), .ZN(new_n728));
  AOI22_X1  g527(.A1(new_n555), .A2(new_n556), .B1(new_n560), .B2(new_n563), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n570), .B1(new_n729), .B2(new_n558), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT107), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n572), .A2(new_n732), .A3(new_n573), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n721), .ZN(new_n735));
  INV_X1    g534(.A(new_n722), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT44), .B1(new_n692), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n452), .A2(KEYINPUT90), .A3(KEYINPUT35), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT90), .B1(new_n452), .B2(KEYINPUT35), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n739), .A2(new_n740), .A3(new_n470), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n738), .B(new_n722), .C1(new_n741), .C2(new_n504), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n735), .B1(new_n737), .B2(new_n742), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n743), .A2(new_n685), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n727), .B1(new_n744), .B2(new_n510), .ZN(G1328gat));
  NAND3_X1  g544(.A1(new_n725), .A2(new_n511), .A3(new_n474), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT46), .Z(new_n747));
  AND2_X1   g546(.A1(new_n743), .A2(new_n474), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(new_n511), .ZN(G1329gat));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n750));
  INV_X1    g549(.A(new_n501), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n743), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n752), .B2(new_n515), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n725), .A2(new_n515), .A3(new_n450), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n752), .B2(new_n515), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT47), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n753), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  OAI221_X1 g556(.A(new_n754), .B1(new_n750), .B2(KEYINPUT47), .C1(new_n752), .C2(new_n515), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(G1330gat));
  INV_X1    g558(.A(KEYINPUT48), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n725), .A2(new_n513), .A3(new_n473), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n513), .B1(new_n743), .B2(new_n473), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n762), .B2(KEYINPUT109), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT109), .ZN(new_n764));
  AOI211_X1 g563(.A(new_n764), .B(new_n513), .C1(new_n743), .C2(new_n473), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n760), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n743), .A2(KEYINPUT110), .A3(new_n473), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G50gat), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT110), .B1(new_n743), .B2(new_n473), .ZN(new_n769));
  OAI211_X1 g568(.A(KEYINPUT48), .B(new_n761), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n766), .A2(new_n770), .ZN(G1331gat));
  INV_X1    g570(.A(new_n677), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n675), .ZN(new_n773));
  NOR4_X1   g572(.A1(new_n692), .A2(new_n654), .A3(new_n773), .A4(new_n734), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n685), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g575(.A1(new_n442), .A2(KEYINPUT111), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n442), .A2(KEYINPUT111), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT49), .ZN(new_n780));
  INV_X1    g579(.A(G64gat), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n782), .B(KEYINPUT112), .Z(new_n783));
  NAND2_X1  g582(.A1(new_n774), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n780), .A2(new_n781), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n784), .B(new_n785), .ZN(G1333gat));
  NAND2_X1  g585(.A1(new_n774), .A2(new_n751), .ZN(new_n787));
  INV_X1    g586(.A(new_n450), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(G71gat), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n787), .A2(G71gat), .B1(new_n774), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n473), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(G78gat), .ZN(G1335gat));
  INV_X1    g592(.A(new_n734), .ZN(new_n794));
  INV_X1    g593(.A(new_n616), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT113), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n506), .A2(new_n722), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n506), .A2(KEYINPUT51), .A3(new_n722), .A4(new_n798), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(KEYINPUT115), .A3(new_n802), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n802), .A2(KEYINPUT115), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n684), .A2(G85gat), .A3(new_n773), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n737), .A2(new_n742), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n797), .A2(new_n773), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(new_n810), .A3(new_n685), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(G85gat), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n810), .B1(new_n809), .B2(new_n685), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n806), .B1(new_n812), .B2(new_n813), .ZN(G1336gat));
  AOI21_X1  g613(.A(new_n630), .B1(new_n809), .B2(new_n474), .ZN(new_n815));
  INV_X1    g614(.A(new_n779), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n816), .A2(G92gat), .A3(new_n773), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n818), .B1(new_n801), .B2(new_n802), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT52), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT116), .B1(new_n809), .B2(new_n779), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n807), .A2(KEYINPUT116), .A3(new_n779), .A4(new_n808), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G92gat), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n803), .A2(new_n804), .A3(new_n817), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n820), .B1(new_n824), .B2(new_n827), .ZN(G1337gat));
  NAND2_X1  g627(.A1(new_n809), .A2(new_n751), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(G99gat), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n788), .A2(G99gat), .A3(new_n773), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n803), .A2(new_n804), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(G1338gat));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n274), .A2(G106gat), .A3(new_n773), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n803), .A2(new_n804), .A3(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n809), .A2(new_n473), .ZN(new_n837));
  INV_X1    g636(.A(G106gat), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n834), .B(new_n836), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n809), .B2(new_n473), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n835), .B(KEYINPUT117), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n841), .B1(new_n801), .B2(new_n802), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT53), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n839), .A2(new_n843), .ZN(G1339gat));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n794), .A2(new_n845), .A3(new_n679), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT118), .B1(new_n680), .B2(new_n734), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n668), .A2(new_n849), .A3(new_n671), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n850), .A2(new_n657), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n664), .A2(new_n666), .A3(new_n670), .A4(new_n667), .ZN(new_n852));
  AND4_X1   g651(.A1(KEYINPUT119), .A2(new_n672), .A3(KEYINPUT54), .A4(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n849), .B1(new_n668), .B2(new_n671), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT119), .B1(new_n854), .B2(new_n852), .ZN(new_n855));
  OAI211_X1 g654(.A(KEYINPUT55), .B(new_n851), .C1(new_n853), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n677), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n672), .A2(KEYINPUT54), .A3(new_n852), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n854), .A2(KEYINPUT119), .A3(new_n852), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT55), .B1(new_n862), .B2(new_n851), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n857), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n560), .A2(new_n563), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n550), .B1(new_n549), .B2(new_n554), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n569), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n864), .A2(new_n573), .A3(new_n722), .A4(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n573), .A2(new_n867), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT120), .B1(new_n869), .B2(new_n773), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n678), .A2(new_n871), .A3(new_n573), .A4(new_n867), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n873), .B1(new_n864), .B2(new_n734), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n868), .B1(new_n874), .B2(new_n722), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n848), .B1(new_n875), .B2(new_n795), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n377), .A2(new_n451), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n684), .A2(new_n779), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n279), .A3(new_n734), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n876), .A2(new_n375), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n885), .A2(new_n693), .A3(new_n881), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n883), .B1(new_n279), .B2(new_n886), .ZN(G1340gat));
  NAND3_X1  g686(.A1(new_n882), .A2(new_n277), .A3(new_n678), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n885), .A2(new_n773), .A3(new_n881), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(new_n277), .ZN(G1341gat));
  AOI21_X1  g689(.A(G127gat), .B1(new_n882), .B2(new_n616), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n885), .A2(new_n881), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n616), .A2(G127gat), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(G1342gat));
  INV_X1    g693(.A(new_n879), .ZN(new_n895));
  INV_X1    g694(.A(G134gat), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n474), .A2(new_n736), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n895), .A2(new_n896), .A3(new_n685), .A4(new_n897), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT56), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n896), .B1(new_n892), .B2(new_n722), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n899), .A2(new_n900), .ZN(G1343gat));
  NAND3_X1  g700(.A1(new_n877), .A2(new_n473), .A3(new_n501), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n880), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(G141gat), .A3(new_n693), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n905), .A2(KEYINPUT58), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n851), .B1(new_n853), .B2(new_n855), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT55), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n909), .A2(new_n574), .A3(new_n677), .A4(new_n856), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n678), .A2(new_n573), .A3(new_n867), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n736), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT121), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n722), .B1(new_n910), .B2(new_n911), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT121), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n915), .A2(new_n868), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n848), .B1(new_n918), .B2(new_n795), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n473), .A2(KEYINPUT57), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT122), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n868), .B1(new_n916), .B2(KEYINPUT121), .ZN(new_n922));
  AOI211_X1 g721(.A(new_n914), .B(new_n722), .C1(new_n910), .C2(new_n911), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n795), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n848), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n920), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT57), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n929), .B1(new_n876), .B2(new_n274), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n921), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n881), .A2(new_n751), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n931), .A2(new_n574), .A3(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n906), .B1(new_n215), .B2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n936), .B1(new_n931), .B2(new_n932), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n930), .B1(new_n926), .B2(new_n927), .ZN(new_n938));
  AOI211_X1 g737(.A(KEYINPUT122), .B(new_n920), .C1(new_n924), .C2(new_n925), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n936), .B(new_n932), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n734), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n905), .B1(new_n942), .B2(G141gat), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT58), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n935), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(KEYINPUT124), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n947), .B(new_n935), .C1(new_n943), .C2(new_n944), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(G1344gat));
  OR2_X1    g748(.A1(new_n937), .A2(new_n941), .ZN(new_n950));
  AOI211_X1 g749(.A(KEYINPUT59), .B(new_n213), .C1(new_n950), .C2(new_n678), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT59), .ZN(new_n952));
  OAI21_X1  g751(.A(KEYINPUT57), .B1(new_n876), .B2(new_n274), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n616), .B1(new_n913), .B2(new_n868), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n680), .A2(new_n574), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n929), .B(new_n473), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n957), .A2(new_n678), .A3(new_n932), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n952), .B1(new_n958), .B2(G148gat), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n678), .A2(new_n213), .ZN(new_n960));
  OAI22_X1  g759(.A1(new_n951), .A2(new_n959), .B1(new_n904), .B2(new_n960), .ZN(G1345gat));
  NOR2_X1   g760(.A1(new_n795), .A2(new_n209), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n903), .A2(new_n616), .A3(new_n880), .ZN(new_n963));
  AOI22_X1  g762(.A1(new_n950), .A2(new_n962), .B1(new_n209), .B2(new_n963), .ZN(G1346gat));
  NAND4_X1  g763(.A1(new_n903), .A2(new_n210), .A3(new_n685), .A4(new_n897), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n950), .A2(new_n722), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n965), .B1(new_n966), .B2(new_n210), .ZN(G1347gat));
  INV_X1    g766(.A(G169gat), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n685), .A2(new_n442), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n970), .A2(new_n885), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n968), .B1(new_n971), .B2(new_n574), .ZN(new_n972));
  XOR2_X1   g771(.A(new_n972), .B(KEYINPUT125), .Z(new_n973));
  NOR2_X1   g772(.A1(new_n685), .A2(new_n816), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n895), .A2(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n976), .A2(new_n968), .A3(new_n734), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n973), .A2(new_n977), .ZN(G1348gat));
  AOI21_X1  g777(.A(G176gat), .B1(new_n976), .B2(new_n678), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n678), .A2(G176gat), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n979), .B1(new_n971), .B2(new_n980), .ZN(G1349gat));
  AOI211_X1 g780(.A(new_n795), .B(new_n975), .C1(new_n327), .C2(new_n328), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n304), .B1(new_n971), .B2(new_n616), .ZN(new_n983));
  NOR3_X1   g782(.A1(new_n982), .A2(KEYINPUT126), .A3(new_n983), .ZN(new_n984));
  XOR2_X1   g783(.A(new_n984), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g784(.A(new_n306), .B1(new_n971), .B2(new_n722), .ZN(new_n986));
  XOR2_X1   g785(.A(new_n986), .B(KEYINPUT61), .Z(new_n987));
  NAND3_X1  g786(.A1(new_n976), .A2(new_n306), .A3(new_n722), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(G1351gat));
  NOR2_X1   g788(.A1(new_n970), .A2(new_n751), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(new_n957), .ZN(new_n991));
  OAI21_X1  g790(.A(G197gat), .B1(new_n991), .B2(new_n693), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n903), .A2(new_n974), .ZN(new_n993));
  OR2_X1    g792(.A1(new_n794), .A2(G197gat), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(G1352gat));
  NOR3_X1   g794(.A1(new_n993), .A2(G204gat), .A3(new_n773), .ZN(new_n996));
  INV_X1    g795(.A(new_n996), .ZN(new_n997));
  OR3_X1    g796(.A1(new_n997), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(KEYINPUT62), .ZN(new_n999));
  OAI21_X1  g798(.A(KEYINPUT127), .B1(new_n997), .B2(KEYINPUT62), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n990), .A2(new_n957), .A3(new_n678), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1001), .A2(G204gat), .ZN(new_n1002));
  NAND4_X1  g801(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .A4(new_n1002), .ZN(G1353gat));
  NAND3_X1  g802(.A1(new_n990), .A2(new_n957), .A3(new_n616), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n1004), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1005));
  INV_X1    g804(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g805(.A(KEYINPUT63), .B1(new_n1004), .B2(G211gat), .ZN(new_n1007));
  OR2_X1    g806(.A1(new_n795), .A2(G211gat), .ZN(new_n1008));
  OAI22_X1  g807(.A1(new_n1006), .A2(new_n1007), .B1(new_n993), .B2(new_n1008), .ZN(G1354gat));
  INV_X1    g808(.A(G218gat), .ZN(new_n1010));
  NOR3_X1   g809(.A1(new_n991), .A2(new_n1010), .A3(new_n736), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n903), .A2(new_n722), .A3(new_n974), .ZN(new_n1012));
  AOI21_X1  g811(.A(new_n1011), .B1(new_n1010), .B2(new_n1012), .ZN(G1355gat));
endmodule


