//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n581, new_n582, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n633, new_n634, new_n635, new_n636, new_n639,
    new_n641, new_n642, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1242, new_n1243, new_n1244;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT67), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n460), .B1(new_n453), .B2(G2106), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT69), .Z(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G101), .ZN(new_n465));
  OAI21_X1  g040(.A(KEYINPUT73), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT73), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n467), .A2(new_n463), .A3(G101), .A4(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT72), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n470), .B1(new_n471), .B2(KEYINPUT3), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(KEYINPUT72), .A3(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n471), .A2(KEYINPUT3), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n472), .A2(new_n474), .A3(new_n463), .A4(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n469), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n473), .A2(G2104), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n479), .A2(new_n475), .A3(G125), .ZN(new_n480));
  INV_X1    g055(.A(G113), .ZN(new_n481));
  OAI21_X1  g056(.A(KEYINPUT70), .B1(new_n481), .B2(new_n471), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n483), .A2(G113), .A3(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(G2105), .B1(new_n480), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT71), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n479), .A2(new_n475), .ZN(new_n488));
  INV_X1    g063(.A(G125), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n482), .B(new_n484), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n490), .A2(new_n491), .A3(G2105), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n478), .B1(new_n487), .B2(new_n492), .ZN(G160));
  NAND4_X1  g068(.A1(new_n472), .A2(new_n474), .A3(G2105), .A4(new_n475), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G124), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n463), .A2(G112), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OR2_X1    g074(.A1(new_n476), .A2(KEYINPUT74), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n476), .A2(KEYINPUT74), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n499), .B1(new_n502), .B2(G136), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT75), .ZN(new_n504));
  XNOR2_X1  g079(.A(new_n503), .B(new_n504), .ZN(G162));
  AND2_X1   g080(.A1(new_n474), .A2(new_n475), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT77), .ZN(new_n507));
  INV_X1    g082(.A(G138), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n508), .A2(G2105), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n506), .A2(new_n507), .A3(new_n472), .A4(new_n509), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n472), .A2(new_n474), .A3(new_n509), .A4(new_n475), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT77), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n510), .A2(KEYINPUT4), .A3(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT4), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n509), .A2(new_n479), .A3(new_n475), .A4(new_n514), .ZN(new_n515));
  OAI21_X1  g090(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n517), .B1(G114), .B2(new_n463), .ZN(new_n518));
  INV_X1    g093(.A(G126), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n494), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT76), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT76), .ZN(new_n522));
  OAI211_X1 g097(.A(new_n518), .B(new_n522), .C1(new_n494), .C2(new_n519), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n513), .A2(new_n515), .B1(new_n521), .B2(new_n523), .ZN(G164));
  NAND2_X1  g099(.A1(G75), .A2(G543), .ZN(new_n525));
  AND2_X1   g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G62), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n525), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G651), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT6), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT78), .B1(new_n532), .B2(G651), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT78), .ZN(new_n534));
  INV_X1    g109(.A(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT6), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n533), .A2(new_n536), .B1(new_n532), .B2(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT5), .B(G543), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n537), .A2(G88), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n533), .A2(new_n536), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n532), .A2(G651), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n540), .A2(G50), .A3(G543), .A4(new_n541), .ZN(new_n542));
  AND3_X1   g117(.A1(new_n539), .A2(new_n542), .A3(KEYINPUT79), .ZN(new_n543));
  AOI21_X1  g118(.A(KEYINPUT79), .B1(new_n539), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n531), .B1(new_n543), .B2(new_n544), .ZN(G303));
  INV_X1    g120(.A(G303), .ZN(G166));
  NAND3_X1  g121(.A1(new_n540), .A2(G543), .A3(new_n541), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(KEYINPUT80), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT80), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n537), .A2(new_n549), .A3(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n551), .A2(G51), .ZN(new_n552));
  NAND3_X1  g127(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT7), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n538), .A2(G63), .A3(G651), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n540), .A2(new_n538), .A3(new_n541), .ZN(new_n556));
  INV_X1    g131(.A(G89), .ZN(new_n557));
  OAI211_X1 g132(.A(new_n554), .B(new_n555), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n552), .A2(new_n558), .ZN(G168));
  NAND2_X1  g134(.A1(new_n551), .A2(G52), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n538), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(new_n535), .ZN(new_n562));
  INV_X1    g137(.A(new_n556), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G90), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n560), .A2(new_n562), .A3(new_n564), .ZN(G301));
  INV_X1    g140(.A(G301), .ZN(G171));
  INV_X1    g141(.A(G43), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n548), .B2(new_n550), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G68), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G56), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n528), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G651), .ZN(new_n573));
  INV_X1    g148(.A(G81), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n574), .B2(new_n556), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G860), .ZN(G153));
  NAND4_X1  g154(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g155(.A1(G1), .A2(G3), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT8), .ZN(new_n582));
  NAND4_X1  g157(.A1(G319), .A2(G483), .A3(G661), .A4(new_n582), .ZN(G188));
  AND3_X1   g158(.A1(new_n537), .A2(G53), .A3(G543), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT9), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n584), .B(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G78), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G65), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n528), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G651), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT81), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n589), .A2(KEYINPUT81), .A3(G651), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n592), .A2(new_n593), .B1(new_n563), .B2(G91), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n586), .A2(new_n594), .ZN(G299));
  INV_X1    g170(.A(G168), .ZN(G286));
  NAND3_X1  g171(.A1(new_n537), .A2(G49), .A3(G543), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n538), .B2(G74), .ZN(new_n598));
  INV_X1    g173(.A(G87), .ZN(new_n599));
  OAI211_X1 g174(.A(new_n597), .B(new_n598), .C1(new_n599), .C2(new_n556), .ZN(G288));
  NAND3_X1  g175(.A1(new_n537), .A2(G86), .A3(new_n538), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n537), .A2(G48), .A3(G543), .ZN(new_n602));
  OAI21_X1  g177(.A(G61), .B1(new_n526), .B2(new_n527), .ZN(new_n603));
  NAND2_X1  g178(.A1(G73), .A2(G543), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(KEYINPUT82), .B1(new_n605), .B2(G651), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT82), .ZN(new_n607));
  AOI211_X1 g182(.A(new_n607), .B(new_n535), .C1(new_n603), .C2(new_n604), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n601), .B(new_n602), .C1(new_n606), .C2(new_n608), .ZN(G305));
  NAND2_X1  g184(.A1(G72), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G60), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n528), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G651), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT83), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n551), .A2(G47), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n563), .A2(G85), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(G290));
  NAND2_X1  g193(.A1(G301), .A2(G868), .ZN(new_n619));
  NAND4_X1  g194(.A1(new_n540), .A2(G92), .A3(new_n538), .A4(new_n541), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT84), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT10), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n620), .A2(KEYINPUT84), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n620), .A2(KEYINPUT84), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(KEYINPUT10), .A3(new_n625), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n538), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n627), .A2(new_n535), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(new_n551), .B2(G54), .ZN(new_n629));
  AND3_X1   g204(.A1(new_n623), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n619), .B1(new_n630), .B2(G868), .ZN(G284));
  OAI21_X1  g206(.A(new_n619), .B1(new_n630), .B2(G868), .ZN(G321));
  NAND2_X1  g207(.A1(G286), .A2(G868), .ZN(new_n633));
  INV_X1    g208(.A(new_n594), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n584), .B(KEYINPUT9), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n633), .B1(G868), .B2(new_n636), .ZN(G297));
  XOR2_X1   g212(.A(G297), .B(KEYINPUT85), .Z(G280));
  INV_X1    g213(.A(G559), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n630), .B1(new_n639), .B2(G860), .ZN(G148));
  NAND2_X1  g215(.A1(new_n630), .A2(new_n639), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(G868), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(G868), .B2(new_n578), .ZN(G323));
  XNOR2_X1  g218(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g219(.A1(new_n502), .A2(G135), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n495), .A2(G123), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n463), .A2(G111), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n645), .B(new_n646), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n649), .A2(G2096), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(G2096), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT12), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT13), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(G2100), .Z(new_n655));
  NAND3_X1  g230(.A1(new_n650), .A2(new_n651), .A3(new_n655), .ZN(G156));
  XOR2_X1   g231(.A(G1341), .B(G1348), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT86), .ZN(new_n658));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT14), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2427), .B(G2438), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2430), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT15), .B(G2435), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n666), .B1(new_n665), .B2(new_n664), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n661), .B(new_n667), .Z(new_n668));
  XNOR2_X1  g243(.A(G2443), .B(G2446), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(G14), .A3(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G401));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT17), .Z(new_n675));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  XOR2_X1   g251(.A(G2084), .B(G2090), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n675), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT87), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(new_n676), .ZN(new_n681));
  INV_X1    g256(.A(new_n674), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n681), .B(new_n678), .C1(new_n682), .C2(new_n676), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n682), .A2(new_n676), .A3(new_n677), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT18), .Z(new_n685));
  NAND3_X1  g260(.A1(new_n680), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G2096), .B(G2100), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G227));
  XOR2_X1   g264(.A(G1971), .B(G1976), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  XOR2_X1   g266(.A(G1956), .B(G2474), .Z(new_n692));
  XOR2_X1   g267(.A(G1961), .B(G1966), .Z(new_n693));
  AND2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT20), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n692), .A2(new_n693), .ZN(new_n697));
  NOR3_X1   g272(.A1(new_n691), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n691), .B2(new_n697), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G1981), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT88), .B(KEYINPUT89), .Z(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n701), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1991), .B(G1996), .ZN(new_n706));
  INV_X1    g281(.A(G1986), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n705), .B(new_n708), .ZN(G229));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G35), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G162), .B2(new_n710), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT103), .B(KEYINPUT29), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT104), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n712), .B(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G2090), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n710), .A2(G32), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n502), .A2(G141), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT98), .ZN(new_n720));
  NAND3_X1  g295(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT26), .Z(new_n722));
  INV_X1    g297(.A(G105), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(new_n464), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G129), .B2(new_n495), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n718), .B1(new_n727), .B2(new_n710), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT99), .Z(new_n729));
  XOR2_X1   g304(.A(KEYINPUT27), .B(G1996), .Z(new_n730));
  AOI21_X1  g305(.A(new_n717), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT31), .B(G11), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT30), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n733), .A2(G28), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n710), .B1(new_n733), .B2(G28), .ZN(new_n735));
  OAI221_X1 g310(.A(new_n732), .B1(new_n734), .B2(new_n735), .C1(new_n649), .C2(new_n710), .ZN(new_n736));
  INV_X1    g311(.A(G2084), .ZN(new_n737));
  NAND2_X1  g312(.A1(G160), .A2(G29), .ZN(new_n738));
  AND2_X1   g313(.A1(KEYINPUT24), .A2(G34), .ZN(new_n739));
  NOR2_X1   g314(.A1(KEYINPUT24), .A2(G34), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n710), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT97), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n736), .B1(new_n737), .B2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G16), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G21), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G168), .B2(new_n745), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n744), .B1(G1966), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n745), .A2(G20), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT23), .Z(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G299), .B2(G16), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(G1956), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n710), .A2(G26), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT28), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n502), .A2(G140), .ZN(new_n755));
  NOR2_X1   g330(.A1(G104), .A2(G2105), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT94), .ZN(new_n757));
  INV_X1    g332(.A(G116), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n471), .B1(new_n758), .B2(G2105), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n495), .A2(G128), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n754), .B1(new_n762), .B2(new_n710), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G2067), .ZN(new_n764));
  NOR3_X1   g339(.A1(new_n748), .A2(new_n752), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(G301), .A2(G16), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n745), .A2(G5), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G1961), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n769), .A2(new_n770), .B1(new_n747), .B2(G1966), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n745), .A2(G19), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n577), .B2(G16), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1341), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n630), .A2(G16), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G4), .B2(G16), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT93), .B(G1348), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n771), .B(new_n774), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n768), .A2(G1961), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT101), .Z(new_n780));
  AOI211_X1 g355(.A(new_n778), .B(new_n780), .C1(new_n776), .C2(new_n777), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n710), .A2(G27), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G164), .B2(new_n710), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT102), .ZN(new_n784));
  INV_X1    g359(.A(G2078), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n715), .B2(new_n716), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n731), .A2(new_n765), .A3(new_n781), .A4(new_n787), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n710), .A2(G33), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n502), .A2(G139), .ZN(new_n790));
  NAND2_X1  g365(.A1(G115), .A2(G2104), .ZN(new_n791));
  INV_X1    g366(.A(G127), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n488), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n463), .B1(new_n793), .B2(KEYINPUT95), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(KEYINPUT95), .B2(new_n793), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT25), .Z(new_n797));
  NAND3_X1  g372(.A1(new_n790), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n789), .B1(new_n798), .B2(G29), .ZN(new_n799));
  INV_X1    g374(.A(G2072), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT96), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(KEYINPUT96), .B1(new_n799), .B2(new_n800), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n738), .A2(G2084), .A3(new_n742), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n799), .B2(new_n800), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g383(.A(KEYINPUT100), .B(new_n808), .C1(new_n729), .C2(new_n730), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT100), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n728), .A2(KEYINPUT99), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n728), .A2(KEYINPUT99), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n730), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n808), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n810), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n809), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n788), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT91), .ZN(new_n818));
  MUX2_X1   g393(.A(G6), .B(G305), .S(G16), .Z(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT32), .B(G1981), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  MUX2_X1   g396(.A(G23), .B(G288), .S(G16), .Z(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT33), .Z(new_n823));
  AOI21_X1  g398(.A(new_n821), .B1(G1976), .B2(new_n823), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n823), .A2(G1976), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n745), .A2(G22), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G166), .B2(new_n745), .ZN(new_n827));
  INV_X1    g402(.A(G1971), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n824), .A2(new_n825), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT34), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT34), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n824), .A2(new_n825), .A3(new_n832), .A4(new_n829), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n745), .A2(G24), .ZN(new_n834));
  INV_X1    g409(.A(G290), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(new_n745), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G1986), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n710), .A2(G25), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n502), .A2(G131), .ZN(new_n839));
  OAI21_X1  g414(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n840));
  INV_X1    g415(.A(G107), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n840), .B1(new_n841), .B2(G2105), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT90), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(G119), .B2(new_n495), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n838), .B1(new_n846), .B2(new_n710), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT35), .B(G1991), .Z(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n847), .B(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n837), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n831), .A2(new_n833), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n818), .B1(new_n852), .B2(KEYINPUT92), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n853), .A2(KEYINPUT36), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n853), .B(KEYINPUT36), .C1(new_n818), .C2(new_n852), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n817), .A2(new_n854), .A3(new_n855), .ZN(G311));
  NAND3_X1  g431(.A1(new_n817), .A2(new_n854), .A3(new_n855), .ZN(G150));
  NAND3_X1  g432(.A1(new_n623), .A2(new_n626), .A3(new_n629), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n858), .A2(new_n639), .ZN(new_n859));
  XNOR2_X1  g434(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(G55), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(new_n548), .B2(new_n550), .ZN(new_n863));
  NAND2_X1  g438(.A1(G80), .A2(G543), .ZN(new_n864));
  INV_X1    g439(.A(G67), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n864), .B1(new_n528), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(G651), .ZN(new_n867));
  INV_X1    g442(.A(G93), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n867), .B1(new_n868), .B2(new_n556), .ZN(new_n869));
  NOR4_X1   g444(.A1(new_n568), .A2(new_n863), .A3(new_n575), .A4(new_n869), .ZN(new_n870));
  OAI22_X1  g445(.A1(new_n568), .A2(new_n575), .B1(new_n863), .B2(new_n869), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n861), .B(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n874), .A2(KEYINPUT39), .ZN(new_n875));
  INV_X1    g450(.A(G860), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(KEYINPUT39), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n863), .A2(new_n869), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n879), .A2(new_n876), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT37), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT106), .ZN(G145));
  XNOR2_X1  g458(.A(new_n845), .B(KEYINPUT107), .ZN(new_n884));
  INV_X1    g459(.A(new_n653), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT107), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n845), .B(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n653), .ZN(new_n889));
  OR2_X1    g464(.A1(G106), .A2(G2105), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n890), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n891));
  INV_X1    g466(.A(G130), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n891), .B1(new_n494), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n893), .B1(new_n502), .B2(G142), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n886), .A2(new_n889), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n894), .B1(new_n886), .B2(new_n889), .ZN(new_n897));
  OAI21_X1  g472(.A(KEYINPUT108), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n726), .A2(new_n761), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n720), .A2(new_n762), .A3(new_n725), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n520), .B1(new_n513), .B2(new_n515), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n902), .B1(new_n899), .B2(new_n900), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n904), .A2(new_n905), .A3(new_n798), .ZN(new_n906));
  INV_X1    g481(.A(new_n798), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n899), .A2(new_n900), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n901), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n907), .B1(new_n909), .B2(new_n903), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n898), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n798), .B1(new_n904), .B2(new_n905), .ZN(new_n912));
  INV_X1    g487(.A(new_n897), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n895), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n909), .A2(new_n903), .A3(new_n907), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n912), .A2(new_n914), .A3(new_n915), .A4(KEYINPUT108), .ZN(new_n916));
  XNOR2_X1  g491(.A(G162), .B(new_n649), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(G160), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n911), .A2(new_n916), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n914), .B1(new_n906), .B2(new_n910), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n912), .A2(new_n915), .A3(new_n895), .A4(new_n913), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n922), .A3(new_n918), .ZN(new_n923));
  INV_X1    g498(.A(G37), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n920), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g501(.A(G305), .B(G288), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n929));
  NAND2_X1  g504(.A1(G303), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g505(.A(KEYINPUT110), .B(new_n531), .C1(new_n543), .C2(new_n544), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(G290), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(G290), .B1(new_n930), .B2(new_n931), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n928), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n934), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(new_n927), .A3(new_n932), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n938), .B(KEYINPUT42), .Z(new_n939));
  XOR2_X1   g514(.A(new_n641), .B(new_n873), .Z(new_n940));
  NAND2_X1  g515(.A1(new_n630), .A2(new_n636), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n858), .A2(G299), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT109), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT41), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n941), .A2(new_n942), .A3(KEYINPUT41), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n945), .B1(new_n940), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n940), .A2(KEYINPUT109), .A3(new_n944), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n939), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n939), .B1(new_n951), .B2(new_n950), .ZN(new_n953));
  OAI21_X1  g528(.A(G868), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(G868), .B2(new_n879), .ZN(G295));
  OAI21_X1  g530(.A(new_n954), .B1(G868), .B2(new_n879), .ZN(G331));
  OAI21_X1  g531(.A(G171), .B1(new_n870), .B2(new_n872), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n551), .A2(G55), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n563), .A2(G93), .B1(new_n866), .B2(G651), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n569), .A2(new_n958), .A3(new_n576), .A4(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n960), .A2(new_n871), .A3(G301), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n957), .A2(G168), .A3(new_n961), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n960), .A2(new_n871), .A3(G301), .ZN(new_n963));
  AOI21_X1  g538(.A(G301), .B1(new_n960), .B2(new_n871), .ZN(new_n964));
  OAI21_X1  g539(.A(G286), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n944), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT112), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n947), .A2(new_n948), .A3(new_n962), .A4(new_n965), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n966), .A2(new_n970), .A3(new_n944), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n968), .A2(new_n938), .A3(new_n969), .A4(new_n971), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n972), .A2(new_n924), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT113), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n967), .A2(new_n969), .ZN(new_n975));
  INV_X1    g550(.A(new_n938), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI211_X1 g552(.A(KEYINPUT113), .B(new_n938), .C1(new_n967), .C2(new_n969), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  XOR2_X1   g554(.A(KEYINPUT111), .B(KEYINPUT43), .Z(new_n980));
  NAND3_X1  g555(.A1(new_n973), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n982));
  INV_X1    g557(.A(new_n980), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n972), .A2(new_n924), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n971), .A2(new_n969), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n938), .B1(new_n985), .B2(new_n968), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n983), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n981), .A2(new_n982), .A3(new_n987), .ZN(new_n988));
  AND4_X1   g563(.A1(new_n947), .A2(new_n948), .A3(new_n962), .A4(new_n965), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n943), .B1(new_n962), .B2(new_n965), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n976), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT113), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n975), .A2(new_n974), .A3(new_n976), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT43), .B1(new_n994), .B2(new_n984), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n985), .A2(new_n968), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n976), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n973), .A2(new_n997), .A3(new_n980), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n982), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n988), .A2(new_n999), .ZN(G397));
  NAND2_X1  g575(.A1(G303), .A2(G8), .ZN(new_n1001));
  XNOR2_X1  g576(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1005), .A2(KEYINPUT55), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1004), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n1008));
  INV_X1    g583(.A(G1384), .ZN(new_n1009));
  INV_X1    g584(.A(new_n515), .ZN(new_n1010));
  AND4_X1   g585(.A1(new_n472), .A2(new_n474), .A3(new_n509), .A4(new_n475), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n514), .B1(new_n1011), .B2(new_n507), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1010), .B1(new_n1012), .B2(new_n512), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1008), .B(new_n1009), .C1(new_n1013), .C2(new_n520), .ZN(new_n1014));
  INV_X1    g589(.A(G40), .ZN(new_n1015));
  AOI211_X1 g590(.A(new_n1015), .B(new_n478), .C1(new_n487), .C2(new_n492), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n521), .A2(new_n523), .ZN(new_n1018));
  INV_X1    g593(.A(new_n512), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT4), .B1(new_n511), .B2(KEYINPUT77), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n515), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1008), .B1(new_n1022), .B2(new_n1009), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1017), .A2(new_n1023), .A3(G2090), .ZN(new_n1024));
  INV_X1    g599(.A(new_n478), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n486), .A2(KEYINPUT71), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n491), .B1(new_n490), .B2(G2105), .ZN(new_n1027));
  OAI211_X1 g602(.A(G40), .B(new_n1025), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n520), .ZN(new_n1029));
  AOI21_X1  g604(.A(G1384), .B1(new_n1021), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1028), .B1(new_n1030), .B2(KEYINPUT45), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT45), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(G164), .B2(G1384), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1971), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1007), .B(G8), .C1(new_n1024), .C2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT49), .ZN(new_n1036));
  INV_X1    g611(.A(G1981), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n538), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n607), .B1(new_n1038), .B2(new_n535), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n605), .A2(KEYINPUT82), .A3(G651), .ZN(new_n1040));
  INV_X1    g615(.A(new_n547), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1039), .A2(new_n1040), .B1(new_n1041), .B2(G48), .ZN(new_n1042));
  XOR2_X1   g617(.A(KEYINPUT116), .B(G86), .Z(new_n1043));
  NAND2_X1  g618(.A1(new_n563), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1037), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(G305), .A2(G1981), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1036), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1044), .B(new_n602), .C1(new_n606), .C2(new_n608), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G1981), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1042), .A2(new_n1037), .A3(new_n601), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(new_n1050), .A3(KEYINPUT49), .ZN(new_n1051));
  INV_X1    g626(.A(G8), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n1016), .B2(new_n1030), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1047), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1976), .ZN(new_n1055));
  OR2_X1    g630(.A1(G288), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1009), .B1(new_n1013), .B2(new_n520), .ZN(new_n1057));
  OAI211_X1 g632(.A(G8), .B(new_n1056), .C1(new_n1057), .C2(new_n1028), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT52), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT52), .B1(G288), .B2(new_n1055), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1053), .A2(new_n1056), .A3(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1054), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(G288), .A2(G1976), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1046), .B1(new_n1054), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1053), .ZN(new_n1065));
  OAI22_X1  g640(.A1(new_n1035), .A2(new_n1062), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g641(.A(KEYINPUT45), .B(new_n1009), .C1(new_n1013), .C2(new_n520), .ZN(new_n1067));
  AOI21_X1  g642(.A(G1384), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1067), .B(new_n1016), .C1(new_n1068), .C2(KEYINPUT45), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n828), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1028), .B1(new_n1030), .B2(new_n1008), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n1072), .A3(new_n716), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1052), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1062), .B1(new_n1074), .B2(new_n1007), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT63), .ZN(new_n1076));
  OAI21_X1  g651(.A(G8), .B1(new_n1024), .B2(new_n1034), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1007), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1966), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1016), .B1(new_n1030), .B2(KEYINPUT45), .ZN(new_n1081));
  AOI211_X1 g656(.A(new_n1032), .B(G1384), .C1(new_n1018), .C2(new_n1021), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1071), .A2(new_n1072), .A3(KEYINPUT117), .A4(new_n737), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1014), .B(new_n1016), .C1(new_n1068), .C2(new_n1008), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(new_n1087), .B2(G2084), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1052), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1075), .A2(new_n1079), .A3(new_n1089), .A4(G168), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1022), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT50), .B1(new_n901), .B2(G1384), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(new_n1092), .A3(new_n1016), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(G2090), .ZN(new_n1094));
  OAI21_X1  g669(.A(G8), .B1(new_n1094), .B2(new_n1034), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1078), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1075), .A2(new_n1089), .A3(new_n1096), .A4(G168), .ZN(new_n1097));
  AOI22_X1  g672(.A1(KEYINPUT118), .A2(new_n1090), .B1(new_n1097), .B2(new_n1076), .ZN(new_n1098));
  OR2_X1    g673(.A1(new_n1090), .A2(KEYINPUT118), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1066), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT119), .B(G1956), .Z(new_n1101));
  NAND2_X1  g676(.A1(new_n1093), .A2(new_n1101), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n634), .A2(new_n635), .A3(KEYINPUT57), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n586), .B2(new_n594), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  XOR2_X1   g681(.A(KEYINPUT56), .B(G2072), .Z(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1031), .A2(new_n1033), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1102), .A2(new_n1106), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(G1348), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1057), .A2(G2067), .A3(new_n1028), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n630), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1102), .A2(new_n1109), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1110), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n1122));
  XOR2_X1   g697(.A(KEYINPUT58), .B(G1341), .Z(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n1057), .B2(new_n1028), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n1069), .B2(G1996), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(KEYINPUT121), .B(new_n1124), .C1(new_n1069), .C2(G1996), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1122), .B1(new_n1129), .B2(new_n578), .ZN(new_n1130));
  AOI211_X1 g705(.A(KEYINPUT59), .B(new_n577), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT60), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1133), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n630), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n1136));
  INV_X1    g711(.A(G1348), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1112), .B1(new_n1087), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1136), .B1(new_n1138), .B2(KEYINPUT60), .ZN(new_n1139));
  NOR4_X1   g714(.A1(new_n1111), .A2(KEYINPUT123), .A3(new_n1133), .A4(new_n1112), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1135), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1137), .B1(new_n1017), .B2(new_n1023), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1112), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1142), .A2(KEYINPUT60), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT123), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1142), .A2(new_n1136), .A3(new_n1143), .A4(KEYINPUT60), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1145), .A2(new_n630), .A3(new_n1134), .A4(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1102), .A2(new_n1106), .A3(new_n1109), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1106), .B1(new_n1102), .B2(new_n1109), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1148), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1118), .A2(new_n1110), .A3(new_n1152), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1141), .A2(new_n1147), .A3(new_n1151), .A4(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1121), .B1(new_n1132), .B2(new_n1154), .ZN(new_n1155));
  XOR2_X1   g730(.A(KEYINPUT125), .B(KEYINPUT54), .Z(new_n1156));
  NAND3_X1  g731(.A1(new_n1031), .A2(new_n1033), .A3(new_n785), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT53), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1087), .A2(new_n770), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1057), .A2(KEYINPUT114), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT114), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1030), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1161), .A2(new_n1032), .A3(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1158), .A2(G2078), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1025), .A2(G40), .A3(new_n486), .A4(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1166), .B1(new_n1030), .B2(KEYINPUT45), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  AND4_X1   g743(.A1(G301), .A2(new_n1159), .A3(new_n1160), .A4(new_n1168), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1157), .A2(new_n1158), .B1(new_n1087), .B2(new_n770), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n1165), .ZN(new_n1172));
  AOI21_X1  g747(.A(G301), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1156), .B1(new_n1169), .B2(new_n1173), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1054), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1035), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1028), .B1(new_n1068), .B2(new_n1008), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1177), .A2(new_n716), .A3(new_n1092), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1070), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1007), .B1(new_n1179), .B2(G8), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1176), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1159), .A2(new_n1168), .A3(new_n1160), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(G171), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1170), .A2(G301), .A3(new_n1172), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1183), .A2(KEYINPUT54), .A3(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1174), .A2(new_n1181), .A3(new_n1185), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1088), .A2(G168), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT51), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1052), .B1(KEYINPUT124), .B2(new_n1188), .ZN(new_n1189));
  OR2_X1    g764(.A1(new_n1188), .A2(KEYINPUT124), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1187), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1088), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1193));
  OAI211_X1 g768(.A(G8), .B(G286), .C1(new_n1192), .C2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1191), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1190), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1186), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1155), .A2(new_n1198), .ZN(new_n1199));
  OR3_X1    g774(.A1(new_n1195), .A2(KEYINPUT62), .A3(new_n1196), .ZN(new_n1200));
  OAI21_X1  g775(.A(KEYINPUT62), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1200), .A2(new_n1201), .A3(new_n1173), .A4(new_n1181), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1100), .A2(new_n1199), .A3(new_n1202), .ZN(new_n1203));
  OR2_X1    g778(.A1(new_n1164), .A2(new_n1028), .ZN(new_n1204));
  INV_X1    g779(.A(new_n1204), .ZN(new_n1205));
  OR2_X1    g780(.A1(new_n761), .A2(G2067), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n761), .A2(G2067), .ZN(new_n1207));
  AND2_X1   g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n845), .B(new_n848), .ZN(new_n1209));
  NOR2_X1   g784(.A1(new_n727), .A2(G1996), .ZN(new_n1210));
  AND3_X1   g785(.A1(new_n720), .A2(G1996), .A3(new_n725), .ZN(new_n1211));
  OAI211_X1 g786(.A(new_n1208), .B(new_n1209), .C1(new_n1210), .C2(new_n1211), .ZN(new_n1212));
  XNOR2_X1  g787(.A(G290), .B(G1986), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1205), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1203), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT47), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1204), .A2(G1996), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT46), .ZN(new_n1218));
  XNOR2_X1  g793(.A(new_n1217), .B(new_n1218), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n727), .A2(new_n1208), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1205), .A2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g796(.A1(new_n1219), .A2(KEYINPUT126), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g797(.A(new_n1222), .ZN(new_n1223));
  AOI21_X1  g798(.A(KEYINPUT126), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1216), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g800(.A1(new_n845), .A2(new_n849), .ZN(new_n1226));
  OAI211_X1 g801(.A(new_n1208), .B(new_n1226), .C1(new_n1210), .C2(new_n1211), .ZN(new_n1227));
  AOI21_X1  g802(.A(new_n1204), .B1(new_n1227), .B2(new_n1206), .ZN(new_n1228));
  AND3_X1   g803(.A1(new_n1212), .A2(KEYINPUT127), .A3(new_n1205), .ZN(new_n1229));
  AOI21_X1  g804(.A(KEYINPUT127), .B1(new_n1212), .B2(new_n1205), .ZN(new_n1230));
  NOR2_X1   g805(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NOR3_X1   g806(.A1(new_n1204), .A2(G1986), .A3(G290), .ZN(new_n1232));
  XOR2_X1   g807(.A(new_n1232), .B(KEYINPUT48), .Z(new_n1233));
  AOI21_X1  g808(.A(new_n1228), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1235));
  INV_X1    g810(.A(KEYINPUT126), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g812(.A1(new_n1237), .A2(KEYINPUT47), .A3(new_n1222), .ZN(new_n1238));
  AND3_X1   g813(.A1(new_n1225), .A2(new_n1234), .A3(new_n1238), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1215), .A2(new_n1239), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g815(.A1(new_n981), .A2(new_n987), .ZN(new_n1242));
  NAND3_X1  g816(.A1(G319), .A2(new_n672), .A3(new_n688), .ZN(new_n1243));
  NOR2_X1   g817(.A1(G229), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g818(.A1(new_n1242), .A2(new_n925), .A3(new_n1244), .ZN(G225));
  INV_X1    g819(.A(G225), .ZN(G308));
endmodule


