//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0004(.A(G50), .B1(G58), .B2(G68), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT64), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n211), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n210), .B1(new_n219), .B2(KEYINPUT0), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G97), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n217), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT67), .Z(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n227));
  INV_X1    g0027(.A(G50), .ZN(new_n228));
  INV_X1    g0028(.A(G226), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT65), .B(G238), .Z(new_n230));
  INV_X1    g0030(.A(G68), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n226), .B1(KEYINPUT66), .B2(new_n232), .ZN(new_n233));
  AND2_X1   g0033(.A1(new_n232), .A2(KEYINPUT66), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n214), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT1), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n220), .B(new_n236), .C1(KEYINPUT0), .C2(new_n219), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(G97), .B(G107), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(KEYINPUT76), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT14), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT13), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT70), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT70), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G1698), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(new_n263), .A3(G226), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G232), .A3(G1698), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G97), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G1), .A3(G13), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G1), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n272), .B1(G41), .B2(G45), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n269), .A2(G238), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT69), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT69), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G45), .ZN(new_n278));
  AOI21_X1  g0078(.A(G41), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n272), .A2(G274), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n274), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n257), .B1(new_n271), .B2(new_n282), .ZN(new_n283));
  AOI211_X1 g0083(.A(KEYINPUT13), .B(new_n281), .C1(new_n267), .C2(new_n270), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G169), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n256), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI221_X1 g0087(.A(G169), .B1(new_n254), .B2(new_n255), .C1(new_n283), .C2(new_n284), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n271), .A2(new_n282), .A3(new_n257), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT75), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n291), .B1(new_n285), .B2(new_n290), .ZN(new_n292));
  INV_X1    g0092(.A(G179), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n287), .B(new_n288), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n207), .ZN(new_n296));
  INV_X1    g0096(.A(G33), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(G20), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n299), .A2(new_n202), .B1(new_n208), .B2(G68), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n208), .A2(new_n297), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(new_n228), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n296), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT11), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n272), .A2(G13), .A3(G20), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT72), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n272), .A2(KEYINPUT72), .A3(G13), .A4(G20), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n231), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT12), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n272), .A2(G20), .ZN(new_n313));
  INV_X1    g0113(.A(new_n296), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n309), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n304), .B(new_n312), .C1(new_n231), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n294), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G200), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n285), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(new_n316), .ZN(new_n320));
  INV_X1    g0120(.A(G190), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n292), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G150), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n201), .A2(new_n208), .B1(new_n301), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n222), .A2(KEYINPUT8), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n222), .A2(KEYINPUT8), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n326), .B1(new_n327), .B2(KEYINPUT71), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(KEYINPUT71), .B2(new_n326), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n325), .B1(new_n329), .B2(new_n298), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(new_n314), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n310), .A2(new_n228), .ZN(new_n333));
  INV_X1    g0133(.A(new_n315), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G50), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n332), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n262), .A2(new_n263), .A3(G222), .ZN(new_n337));
  INV_X1    g0137(.A(G223), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n263), .A2(G1698), .ZN(new_n339));
  OAI221_X1 g0139(.A(new_n337), .B1(new_n202), .B2(new_n263), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n270), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n279), .A2(new_n280), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n269), .A2(new_n273), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n342), .B1(G226), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n336), .B1(new_n347), .B2(G169), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n346), .A2(G179), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n347), .A2(KEYINPUT74), .A3(G190), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT74), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n346), .B2(new_n321), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n335), .A2(new_n333), .ZN(new_n355));
  OR3_X1    g0155(.A1(new_n355), .A2(KEYINPUT9), .A3(new_n331), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT9), .B1(new_n355), .B2(new_n331), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n346), .A2(G200), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n354), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT10), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT10), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n354), .A2(new_n358), .A3(new_n362), .A4(new_n359), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n350), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n262), .A2(new_n263), .A3(G232), .ZN(new_n365));
  INV_X1    g0165(.A(G107), .ZN(new_n366));
  OAI221_X1 g0166(.A(new_n365), .B1(new_n366), .B2(new_n263), .C1(new_n230), .C2(new_n339), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n270), .ZN(new_n368));
  INV_X1    g0168(.A(G244), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n279), .A2(new_n280), .B1(new_n343), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n334), .A2(G77), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G20), .A2(G77), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT15), .B(G87), .ZN(new_n375));
  INV_X1    g0175(.A(new_n326), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n376), .A2(new_n327), .ZN(new_n377));
  OAI221_X1 g0177(.A(new_n374), .B1(new_n375), .B2(new_n299), .C1(new_n377), .C2(new_n301), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n378), .A2(new_n296), .B1(new_n202), .B2(new_n310), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n372), .A2(new_n286), .B1(new_n373), .B2(new_n379), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n372), .A2(KEYINPUT73), .A3(G179), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT73), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n370), .B1(new_n367), .B2(new_n270), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n382), .B1(new_n383), .B2(new_n293), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n380), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n373), .B(new_n379), .C1(new_n372), .C2(new_n321), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n383), .A2(new_n318), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n323), .A2(new_n364), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n342), .B1(G232), .B2(new_n344), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT70), .B(G1698), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n394), .A2(new_n338), .B1(new_n229), .B2(new_n258), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT3), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G33), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  XNOR2_X1  g0198(.A(KEYINPUT77), .B(G33), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n398), .B1(new_n399), .B2(KEYINPUT3), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n395), .A2(new_n400), .B1(G33), .B2(G87), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT81), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n270), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n262), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n404));
  AND2_X1   g0204(.A1(KEYINPUT77), .A2(G33), .ZN(new_n405));
  NOR2_X1   g0205(.A1(KEYINPUT77), .A2(G33), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT3), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n397), .ZN(new_n408));
  INV_X1    g0208(.A(G87), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n404), .A2(new_n408), .B1(new_n297), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n410), .A2(KEYINPUT81), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n293), .B(new_n393), .C1(new_n403), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT82), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n269), .B1(new_n410), .B2(KEYINPUT81), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n401), .A2(new_n402), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT82), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n416), .A2(new_n417), .A3(new_n293), .A4(new_n393), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n393), .B1(new_n403), .B2(new_n411), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n286), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n413), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT7), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n400), .B2(G20), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT78), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n408), .A2(new_n425), .A3(KEYINPUT7), .A4(new_n208), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(G20), .B1(new_n407), .B2(new_n397), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n425), .B1(new_n428), .B2(KEYINPUT7), .ZN(new_n429));
  OAI21_X1  g0229(.A(G68), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n222), .A2(new_n231), .ZN(new_n431));
  NOR2_X1   g0231(.A1(G58), .A2(G68), .ZN(new_n432));
  OAI21_X1  g0232(.A(G20), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G159), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n433), .B1(new_n434), .B2(new_n301), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT79), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n433), .B(KEYINPUT79), .C1(new_n434), .C2(new_n301), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n430), .A2(KEYINPUT16), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT16), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n423), .A2(G20), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT3), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n297), .A2(KEYINPUT3), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n443), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n423), .B1(new_n263), .B2(G20), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n231), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n442), .B1(new_n439), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n441), .A2(new_n296), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n315), .A2(new_n329), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n329), .B2(new_n310), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT80), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT80), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n452), .B(new_n455), .C1(new_n329), .C2(new_n310), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n451), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n422), .A2(KEYINPUT18), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT18), .ZN(new_n461));
  OR2_X1    g0261(.A1(KEYINPUT77), .A2(G33), .ZN(new_n462));
  NAND2_X1  g0262(.A1(KEYINPUT77), .A2(G33), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n396), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g0264(.A(KEYINPUT7), .B(new_n208), .C1(new_n464), .C2(new_n398), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT78), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(new_n424), .A3(new_n426), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n439), .B1(new_n467), .B2(G68), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n314), .B1(new_n468), .B2(KEYINPUT16), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n457), .B1(new_n469), .B2(new_n450), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n461), .B1(new_n470), .B2(new_n421), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT17), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n321), .B(new_n393), .C1(new_n403), .C2(new_n411), .ZN(new_n473));
  INV_X1    g0273(.A(new_n393), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n474), .B1(new_n414), .B2(new_n415), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n473), .B1(new_n475), .B2(G200), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n470), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n451), .A2(new_n476), .A3(new_n458), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT17), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n460), .A2(new_n471), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT83), .B1(new_n392), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT83), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT18), .B1(new_n422), .B2(new_n459), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n470), .A2(new_n421), .A3(new_n461), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n472), .B1(new_n470), .B2(new_n476), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n478), .A2(KEYINPUT17), .ZN(new_n486));
  OAI22_X1  g0286(.A1(new_n483), .A2(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR3_X1   g0287(.A1(new_n391), .A2(new_n482), .A3(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n481), .A2(new_n488), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n272), .A2(KEYINPUT84), .A3(G33), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT84), .B1(new_n272), .B2(G33), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n309), .A2(new_n314), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n375), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n407), .A2(new_n208), .A3(G68), .A4(new_n397), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT19), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n208), .B1(new_n266), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n409), .A2(new_n224), .A3(new_n366), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n208), .A2(G33), .A3(G97), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n498), .A2(new_n499), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n296), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n309), .A2(new_n494), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n495), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n269), .B(G250), .C1(G1), .C2(new_n275), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n275), .A2(G1), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G274), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G116), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n399), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(G238), .ZN(new_n514));
  OAI22_X1  g0314(.A1(new_n394), .A2(new_n514), .B1(new_n369), .B2(new_n258), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n513), .B1(new_n515), .B2(new_n400), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n293), .B(new_n511), .C1(new_n516), .C2(new_n269), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n405), .A2(new_n406), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G116), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n262), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n519), .B1(new_n520), .B2(new_n408), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n510), .B1(new_n521), .B2(new_n270), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n506), .B(new_n517), .C1(G169), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(G190), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n511), .B1(new_n516), .B2(new_n269), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G200), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n309), .A2(new_n492), .A3(new_n314), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n527), .A2(new_n409), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n314), .B1(new_n496), .B2(new_n501), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n528), .A2(new_n529), .A3(new_n504), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n524), .A2(new_n526), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT22), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n397), .A2(new_n445), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n208), .A2(G87), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n366), .A2(G20), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT23), .ZN(new_n537));
  XNOR2_X1  g0337(.A(new_n536), .B(new_n537), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n532), .A2(new_n409), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n513), .B1(new_n400), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n539), .B(KEYINPUT24), .C1(new_n541), .C2(G20), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT24), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n407), .A2(new_n397), .A3(new_n540), .ZN(new_n544));
  AOI21_X1  g0344(.A(G20), .B1(new_n544), .B2(new_n519), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n535), .A2(new_n538), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n543), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n542), .A2(new_n547), .A3(new_n296), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT25), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n309), .B2(G107), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n310), .A2(KEYINPUT25), .A3(new_n366), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n550), .A2(new_n551), .B1(new_n493), .B2(G107), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT5), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n272), .B(G45), .C1(new_n554), .C2(G41), .ZN(new_n555));
  INV_X1    g0355(.A(G41), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(KEYINPUT5), .ZN(new_n557));
  OAI211_X1 g0357(.A(G264), .B(new_n269), .C1(new_n555), .C2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n557), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n556), .A2(KEYINPUT5), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n559), .A2(G274), .A3(new_n508), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  OAI22_X1  g0363(.A1(new_n394), .A2(new_n211), .B1(new_n217), .B2(new_n258), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n564), .A2(new_n400), .B1(G294), .B2(new_n518), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n563), .B1(new_n565), .B2(new_n269), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G200), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n518), .A2(G294), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n217), .A2(new_n258), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n569), .B1(new_n262), .B2(G250), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n568), .B1(new_n570), .B2(new_n408), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n562), .B1(new_n571), .B2(new_n270), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(G190), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n567), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n523), .B(new_n531), .C1(new_n553), .C2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n394), .A2(new_n369), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT4), .B1(new_n400), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g0377(.A1(KEYINPUT4), .A2(G244), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n262), .A2(new_n263), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n263), .A2(G250), .A3(G1698), .ZN(new_n580));
  NAND2_X1  g0380(.A1(G33), .A2(G283), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n270), .B1(new_n577), .B2(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(G257), .B(new_n269), .C1(new_n555), .C2(new_n557), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n583), .A2(new_n321), .A3(new_n561), .A4(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(new_n561), .A3(new_n584), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n318), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n366), .B1(new_n447), .B2(new_n448), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n366), .A2(G97), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT6), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n590), .B2(new_n251), .ZN(new_n592));
  OAI22_X1  g0392(.A1(new_n592), .A2(new_n208), .B1(new_n202), .B2(new_n301), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n296), .B1(new_n588), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n309), .A2(G97), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n595), .B1(new_n493), .B2(G97), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n596), .A3(KEYINPUT85), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT85), .ZN(new_n598));
  INV_X1    g0398(.A(new_n443), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n462), .A2(new_n396), .A3(new_n463), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n599), .B1(new_n600), .B2(new_n445), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT7), .B1(new_n533), .B2(new_n208), .ZN(new_n602));
  OAI21_X1  g0402(.A(G107), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n301), .A2(new_n202), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n224), .A2(G107), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n589), .A2(new_n605), .A3(new_n590), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n590), .B2(new_n589), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n604), .B1(new_n607), .B2(G20), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n314), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n595), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n527), .B2(new_n224), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n598), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n585), .A2(new_n587), .B1(new_n597), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n586), .A2(G169), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n583), .A2(G179), .A3(new_n561), .A4(new_n584), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n614), .A2(new_n615), .B1(new_n594), .B2(new_n596), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n575), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT86), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n310), .A2(new_n512), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n309), .A2(new_n492), .A3(new_n314), .A4(G116), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n295), .A2(new_n207), .B1(G20), .B2(new_n512), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n581), .B(new_n208), .C1(G33), .C2(new_n224), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT20), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT20), .B1(new_n622), .B2(new_n623), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n618), .B1(new_n621), .B2(new_n628), .ZN(new_n629));
  XNOR2_X1  g0429(.A(new_n624), .B(new_n625), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n630), .A2(KEYINPUT86), .A3(new_n620), .A4(new_n619), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  OAI22_X1  g0432(.A1(new_n394), .A2(new_n217), .B1(new_n218), .B2(new_n258), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n633), .A2(new_n400), .ZN(new_n634));
  INV_X1    g0434(.A(G303), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n263), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n270), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  OAI211_X1 g0437(.A(G270), .B(new_n269), .C1(new_n555), .C2(new_n557), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n638), .A2(new_n561), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n286), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n632), .A2(KEYINPUT21), .A3(new_n640), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n633), .A2(new_n400), .B1(G303), .B2(new_n533), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n639), .B1(new_n642), .B2(new_n269), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(new_n293), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n632), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT21), .B1(new_n632), .B2(new_n640), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n318), .B1(new_n637), .B2(new_n639), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n643), .A2(new_n321), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n632), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n646), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT87), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n572), .B2(new_n286), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n566), .A2(KEYINPUT87), .A3(G169), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n653), .B(new_n654), .C1(new_n293), .C2(new_n566), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n553), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n617), .A2(new_n651), .A3(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n489), .A2(new_n657), .ZN(G372));
  INV_X1    g0458(.A(new_n350), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n317), .A2(new_n385), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n477), .A2(new_n479), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(new_n661), .A3(new_n322), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n460), .A2(new_n471), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n361), .A2(new_n363), .ZN(new_n665));
  OAI211_X1 g0465(.A(KEYINPUT88), .B(new_n659), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT88), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n665), .B1(new_n662), .B2(new_n663), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n667), .B1(new_n668), .B2(new_n350), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n614), .A2(new_n615), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n594), .A2(new_n596), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n531), .A2(new_n523), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT26), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n531), .A2(new_n523), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n597), .A2(new_n612), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n676), .A2(new_n677), .A3(new_n679), .A4(new_n671), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n675), .A2(new_n680), .A3(new_n523), .ZN(new_n681));
  INV_X1    g0481(.A(new_n646), .ZN(new_n682));
  INV_X1    g0482(.A(new_n647), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(new_n656), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n617), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n670), .B1(new_n489), .B2(new_n686), .ZN(G369));
  NAND3_X1  g0487(.A1(new_n272), .A2(new_n208), .A3(G13), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT89), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n688), .A2(new_n689), .A3(KEYINPUT27), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n689), .B1(new_n688), .B2(KEYINPUT27), .ZN(new_n691));
  OAI221_X1 g0491(.A(G213), .B1(KEYINPUT27), .B2(new_n688), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(G343), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n632), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n651), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n646), .A2(new_n647), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n696), .B1(new_n697), .B2(new_n695), .ZN(new_n698));
  XOR2_X1   g0498(.A(KEYINPUT90), .B(G330), .Z(new_n699));
  AND2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n656), .A2(new_n694), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n553), .A2(new_n694), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n553), .B2(new_n574), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n701), .B1(new_n656), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n694), .B1(new_n682), .B2(new_n683), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n700), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n704), .A2(new_n705), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(new_n701), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n707), .A2(new_n709), .ZN(G399));
  NOR2_X1   g0510(.A1(new_n216), .A2(G41), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n499), .A2(G116), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n711), .A2(new_n272), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n206), .B2(new_n711), .ZN(new_n715));
  XOR2_X1   g0515(.A(new_n715), .B(KEYINPUT28), .Z(new_n716));
  AOI21_X1  g0516(.A(new_n678), .B1(new_n614), .B2(new_n615), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n676), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT26), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n676), .A2(new_n677), .A3(new_n616), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n719), .A2(new_n523), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n684), .A2(KEYINPUT92), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT92), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n697), .A2(new_n723), .A3(new_n656), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n722), .A2(new_n617), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n694), .B1(new_n721), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT29), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n694), .B1(new_n681), .B2(new_n685), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n728), .A2(KEYINPUT29), .ZN(new_n729));
  INV_X1    g0529(.A(new_n694), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n617), .A2(new_n651), .A3(new_n656), .A4(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT30), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n522), .A2(new_n572), .A3(new_n583), .A4(new_n584), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n637), .A2(G179), .A3(new_n639), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n522), .A2(G179), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n736), .A2(new_n586), .A3(new_n643), .A4(new_n566), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(KEYINPUT91), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n566), .A2(new_n525), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n740), .A2(new_n644), .A3(new_n584), .A4(new_n583), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n741), .A2(new_n732), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT91), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n735), .A2(new_n743), .A3(new_n737), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n739), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT31), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n730), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n741), .A2(new_n732), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n694), .B1(new_n749), .B2(new_n738), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n746), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n731), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n727), .A2(new_n729), .B1(new_n699), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n716), .B1(new_n753), .B2(G1), .ZN(G364));
  INV_X1    g0554(.A(new_n711), .ZN(new_n755));
  INV_X1    g0555(.A(G13), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n272), .B1(new_n757), .B2(G45), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n700), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(new_n699), .B2(new_n698), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n207), .B1(G20), .B2(new_n286), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n293), .A2(new_n318), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n208), .A2(new_n321), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n208), .A2(G190), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n293), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n767), .A2(new_n228), .B1(new_n770), .B2(new_n202), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n318), .A2(G179), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n766), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n768), .A2(new_n772), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G87), .A2(new_n774), .B1(new_n776), .B2(G107), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n766), .A2(new_n769), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n777), .B(new_n263), .C1(new_n222), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n765), .A2(new_n768), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n771), .B(new_n779), .C1(G68), .C2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n293), .A2(new_n318), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT93), .ZN(new_n784));
  INV_X1    g0584(.A(new_n768), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G159), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT32), .Z(new_n788));
  OAI21_X1  g0588(.A(G20), .B1(new_n784), .B2(new_n321), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n782), .B(new_n788), .C1(new_n224), .C2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n773), .B(KEYINPUT94), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n793), .A2(G303), .B1(G329), .B2(new_n786), .ZN(new_n794));
  INV_X1    g0594(.A(G311), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n533), .B1(new_n770), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(G326), .ZN(new_n797));
  INV_X1    g0597(.A(G322), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n767), .A2(new_n797), .B1(new_n778), .B2(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n796), .B(new_n799), .C1(G283), .C2(new_n776), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT95), .B(KEYINPUT33), .Z(new_n801));
  AOI21_X1  g0601(.A(new_n780), .B1(new_n801), .B2(G317), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(G317), .B2(new_n801), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n789), .A2(G294), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n794), .A2(new_n800), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n764), .B1(new_n791), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n216), .A2(new_n533), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G355), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(G116), .B2(new_n215), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n216), .A2(new_n400), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n276), .A2(new_n278), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n811), .B1(new_n206), .B2(new_n812), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n249), .A2(new_n275), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n809), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(G13), .A2(G33), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(G20), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n763), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n760), .B1(new_n815), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n806), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n818), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n698), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n762), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G396));
  NAND2_X1  g0626(.A1(new_n379), .A2(new_n373), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n694), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n387), .B2(new_n388), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n385), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT100), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n380), .B(new_n730), .C1(new_n381), .C2(new_n384), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n831), .B1(new_n830), .B2(new_n832), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n728), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n752), .A2(new_n699), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n760), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n838), .B2(new_n837), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n764), .A2(new_n817), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n760), .B1(G77), .B2(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT96), .ZN(new_n843));
  INV_X1    g0643(.A(new_n778), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n263), .B1(new_n844), .B2(G294), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n845), .B1(new_n409), .B2(new_n775), .C1(new_n792), .C2(new_n366), .ZN(new_n846));
  INV_X1    g0646(.A(new_n767), .ZN(new_n847));
  INV_X1    g0647(.A(new_n770), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n847), .A2(G303), .B1(new_n848), .B2(G116), .ZN(new_n849));
  INV_X1    g0649(.A(G283), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n849), .B1(new_n850), .B2(new_n780), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT97), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n851), .A2(new_n852), .B1(G97), .B2(new_n789), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n852), .B2(new_n851), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n846), .B(new_n854), .C1(G311), .C2(new_n786), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n847), .A2(G137), .B1(new_n848), .B2(G159), .ZN(new_n856));
  INV_X1    g0656(.A(G143), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n856), .B1(new_n857), .B2(new_n778), .C1(new_n324), .C2(new_n780), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT34), .Z(new_n859));
  OAI21_X1  g0659(.A(new_n400), .B1(new_n231), .B2(new_n775), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(G132), .B2(new_n786), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n861), .B1(new_n228), .B2(new_n792), .C1(new_n222), .C2(new_n790), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n859), .B1(KEYINPUT98), .B2(new_n862), .ZN(new_n863));
  OR2_X1    g0663(.A1(new_n862), .A2(KEYINPUT98), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n855), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n843), .B1(new_n865), .B2(new_n764), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n866), .B(KEYINPUT99), .Z(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n817), .B2(new_n836), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n840), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(G384));
  OR2_X1    g0670(.A1(new_n607), .A2(KEYINPUT35), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n871), .A2(G116), .A3(new_n209), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(KEYINPUT35), .B2(new_n607), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n873), .A2(KEYINPUT36), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(KEYINPUT36), .ZN(new_n875));
  OAI21_X1  g0675(.A(G77), .B1(new_n222), .B2(new_n231), .ZN(new_n876));
  OAI22_X1  g0676(.A1(new_n876), .A2(new_n205), .B1(G50), .B2(new_n231), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(G1), .A3(new_n756), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n874), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT101), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n287), .A2(new_n288), .ZN(new_n881));
  INV_X1    g0681(.A(new_n283), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(new_n290), .A3(new_n289), .ZN(new_n883));
  INV_X1    g0683(.A(new_n291), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n293), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n316), .B(new_n694), .C1(new_n881), .C2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT102), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n294), .A2(KEYINPUT102), .A3(new_n316), .A4(new_n694), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n316), .A2(new_n694), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n317), .A2(new_n322), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(KEYINPUT31), .B(new_n694), .C1(new_n749), .C2(new_n738), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n731), .A2(new_n751), .A3(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT40), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT106), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n893), .A2(new_n895), .A3(new_n836), .A4(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n692), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n459), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT105), .B1(new_n480), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT105), .ZN(new_n902));
  INV_X1    g0702(.A(new_n900), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n487), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n478), .B1(new_n470), .B2(new_n692), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n470), .A2(new_n421), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT37), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n478), .B(new_n900), .C1(new_n906), .C2(KEYINPUT104), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT37), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n422), .A2(new_n459), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT104), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n907), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n901), .A2(new_n904), .A3(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT38), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n441), .A2(new_n296), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n468), .A2(KEYINPUT16), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n458), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT103), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT103), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n921), .B(new_n458), .C1(new_n917), .C2(new_n918), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n920), .A2(new_n899), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n920), .A2(new_n422), .A3(new_n922), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(new_n924), .A3(new_n478), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT37), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT104), .B1(new_n422), .B2(new_n459), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n927), .A2(new_n905), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT37), .B1(new_n906), .B2(KEYINPUT104), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n480), .A2(new_n923), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n931), .A2(KEYINPUT38), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n898), .B1(new_n916), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT38), .B1(new_n931), .B2(new_n933), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n925), .A2(KEYINPUT37), .B1(new_n929), .B2(new_n928), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n937), .A2(new_n915), .A3(new_n932), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n895), .A2(new_n836), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n323), .A2(new_n891), .B1(new_n888), .B2(new_n889), .ZN(new_n941));
  OAI21_X1  g0741(.A(KEYINPUT106), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n898), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n935), .A2(new_n896), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n895), .B1(new_n481), .B2(new_n488), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n944), .B(new_n945), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n946), .A2(new_n699), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n294), .A2(new_n316), .A3(new_n730), .ZN(new_n948));
  OAI21_X1  g0748(.A(KEYINPUT39), .B1(new_n936), .B2(new_n938), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT39), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n916), .A2(new_n934), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n948), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n728), .A2(new_n836), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n832), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n893), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n939), .A2(new_n955), .B1(new_n663), .B2(new_n899), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n729), .B(new_n727), .C1(new_n481), .C2(new_n488), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n670), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n957), .B(new_n959), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n947), .A2(new_n960), .B1(new_n272), .B2(new_n757), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n947), .A2(new_n960), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n880), .B1(new_n961), .B2(new_n962), .ZN(G367));
  NAND2_X1  g0763(.A1(new_n245), .A2(new_n810), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n820), .B1(new_n216), .B2(new_n494), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n759), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n730), .A2(new_n530), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT107), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n676), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n523), .B2(new_n969), .ZN(new_n971));
  AOI22_X1  g0771(.A1(G150), .A2(new_n844), .B1(new_n781), .B2(G159), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n222), .B2(new_n773), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n263), .B1(new_n770), .B2(new_n228), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n767), .A2(new_n857), .B1(new_n775), .B2(new_n202), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n789), .A2(G68), .ZN(new_n977));
  INV_X1    g0777(.A(G137), .ZN(new_n978));
  INV_X1    g0778(.A(new_n786), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n976), .B(new_n977), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT113), .Z(new_n981));
  AOI22_X1  g0781(.A1(G97), .A2(new_n776), .B1(new_n848), .B2(G283), .ZN(new_n982));
  INV_X1    g0782(.A(G294), .ZN(new_n983));
  INV_X1    g0783(.A(G317), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n982), .B1(new_n983), .B2(new_n780), .C1(new_n979), .C2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(KEYINPUT46), .B1(new_n774), .B2(G116), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n767), .A2(new_n795), .B1(new_n778), .B2(new_n635), .ZN(new_n987));
  NOR4_X1   g0787(.A1(new_n985), .A2(new_n400), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n793), .A2(KEYINPUT46), .A3(G116), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT112), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n989), .A2(new_n990), .B1(G107), .B2(new_n789), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n988), .B(new_n991), .C1(new_n990), .C2(new_n989), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n981), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n994), .A2(KEYINPUT47), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n763), .B1(new_n994), .B2(KEYINPUT47), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n966), .B1(new_n971), .B2(new_n823), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n758), .B(KEYINPUT111), .Z(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n613), .A2(new_n616), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n678), .B2(new_n730), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n717), .A2(new_n694), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n709), .A2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT45), .Z(new_n1006));
  NOR2_X1   g0806(.A1(new_n709), .A2(new_n1004), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT44), .ZN(new_n1008));
  AOI21_X1  g0808(.A(KEYINPUT109), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(new_n707), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n707), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n700), .A2(new_n706), .ZN(new_n1012));
  NOR3_X1   g0812(.A1(new_n1011), .A2(new_n708), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n753), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT110), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1010), .A2(new_n1015), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1016), .A2(new_n753), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n711), .B(KEYINPUT41), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1000), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1004), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n673), .B1(new_n1021), .B2(new_n656), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n708), .A2(new_n1001), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n730), .A2(new_n1022), .B1(new_n1023), .B2(KEYINPUT42), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(KEYINPUT42), .B2(new_n1023), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1027), .B(new_n1028), .Z(new_n1029));
  NOR2_X1   g0829(.A1(new_n707), .A2(new_n1021), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1031), .B1(new_n1032), .B2(KEYINPUT108), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(KEYINPUT108), .B2(new_n1032), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n998), .B1(new_n1020), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(G387));
  AOI22_X1  g0836(.A1(new_n807), .A2(new_n713), .B1(new_n366), .B2(new_n216), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n377), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n228), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT50), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  AOI211_X1 g0841(.A(G45), .B(new_n713), .C1(G68), .C2(G77), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n811), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT114), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n241), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n1043), .A2(new_n1044), .B1(new_n1045), .B2(new_n812), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1043), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1047), .A2(KEYINPUT114), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1037), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n1049), .A2(KEYINPUT115), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1049), .A2(KEYINPUT115), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n1050), .A2(new_n1051), .A3(new_n820), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n773), .A2(new_n202), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G68), .B2(new_n848), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n228), .B2(new_n778), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n767), .A2(new_n434), .B1(new_n775), .B2(new_n224), .ZN(new_n1056));
  NOR3_X1   g0856(.A1(new_n1055), .A2(new_n408), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n789), .A2(new_n494), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n786), .A2(G150), .B1(new_n329), .B2(new_n781), .ZN(new_n1059));
  AND3_X1   g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n847), .A2(G322), .B1(new_n848), .B2(G303), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n795), .B2(new_n780), .C1(new_n984), .C2(new_n778), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT48), .Z(new_n1063));
  OAI22_X1  g0863(.A1(new_n790), .A2(new_n850), .B1(new_n983), .B2(new_n773), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  XOR2_X1   g0865(.A(KEYINPUT116), .B(KEYINPUT49), .Z(new_n1066));
  OR2_X1    g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n408), .B1(new_n512), .B2(new_n775), .C1(new_n979), .C2(new_n797), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1060), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n760), .B1(new_n1070), .B2(new_n764), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n704), .A2(new_n823), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n1052), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n1013), .B2(new_n999), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1014), .A2(new_n711), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1013), .A2(new_n753), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(G393));
  NAND2_X1  g0877(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(KEYINPUT117), .B2(new_n1011), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1011), .A2(KEYINPUT117), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1079), .B(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1021), .A2(new_n818), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n819), .B1(new_n224), .B2(new_n215), .C1(new_n811), .C2(new_n252), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n760), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G317), .A2(new_n847), .B1(new_n844), .B2(G311), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1086), .A2(KEYINPUT52), .B1(new_n786), .B2(G322), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(KEYINPUT52), .B2(new_n1086), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n780), .A2(new_n635), .B1(new_n770), .B2(new_n983), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G283), .B2(new_n774), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n263), .B1(new_n776), .B2(G107), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(new_n790), .C2(new_n512), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n767), .A2(new_n324), .B1(new_n778), .B2(new_n434), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT51), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n786), .A2(G143), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n1094), .B2(new_n1093), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n789), .A2(G77), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G50), .A2(new_n781), .B1(new_n776), .B2(G87), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1038), .A2(new_n848), .B1(new_n774), .B2(G68), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1097), .A2(new_n400), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1088), .A2(new_n1092), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1085), .B1(new_n1101), .B2(new_n763), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1082), .A2(new_n999), .B1(new_n1083), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1081), .A2(new_n1014), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1104), .A2(new_n711), .A3(new_n1016), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1103), .A2(new_n1105), .ZN(G390));
  NAND2_X1  g0906(.A1(new_n955), .A2(new_n948), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n949), .A2(new_n951), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n916), .A2(new_n934), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n832), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n726), .B2(new_n836), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1109), .B(new_n948), .C1(new_n941), .C2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n893), .A2(new_n895), .A3(G330), .A4(new_n836), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(G330), .B(new_n895), .C1(new_n481), .C2(new_n488), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n958), .A2(new_n1117), .A3(new_n670), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n752), .A2(new_n836), .A3(new_n699), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n941), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n1114), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n954), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT118), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1121), .A2(KEYINPUT118), .A3(new_n954), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  OR2_X1    g0926(.A1(new_n1119), .A2(new_n941), .ZN(new_n1127));
  INV_X1    g0927(.A(G330), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n941), .B1(new_n940), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1127), .A2(new_n1111), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1118), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1108), .A2(new_n1112), .A3(new_n1127), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1116), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(KEYINPUT118), .B1(new_n1121), .B2(new_n954), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1110), .B1(new_n728), .B2(new_n836), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1123), .B(new_n1135), .C1(new_n1120), .C2(new_n1114), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1130), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n958), .A2(new_n1117), .A3(new_n670), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1108), .A2(new_n1127), .A3(new_n1112), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1114), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1133), .A2(new_n1142), .A3(new_n711), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n949), .A2(new_n816), .A3(new_n951), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n760), .B1(new_n329), .B2(new_n841), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n793), .A2(G87), .B1(G294), .B2(new_n786), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n263), .B1(new_n776), .B2(G68), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n767), .A2(new_n850), .B1(new_n780), .B2(new_n366), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n778), .A2(new_n512), .B1(new_n770), .B2(new_n224), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1147), .A2(new_n1097), .A3(new_n1148), .A4(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(G128), .ZN(new_n1153));
  INV_X1    g0953(.A(G132), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n767), .A2(new_n1153), .B1(new_n778), .B2(new_n1154), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT119), .Z(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n434), .B2(new_n790), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n773), .A2(new_n324), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT53), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n786), .A2(G125), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n533), .B1(new_n781), .B2(G137), .ZN(new_n1161));
  XOR2_X1   g0961(.A(KEYINPUT54), .B(G143), .Z(new_n1162));
  AOI22_X1  g0962(.A1(new_n848), .A2(new_n1162), .B1(new_n776), .B2(G50), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .A4(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1152), .B1(new_n1157), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1146), .B1(new_n1165), .B2(new_n763), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1144), .A2(new_n999), .B1(new_n1145), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1143), .A2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT120), .ZN(G378));
  INV_X1    g0969(.A(new_n957), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n336), .A2(new_n899), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n364), .B(new_n1171), .Z(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1172), .B(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n898), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n896), .B1(new_n1109), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n915), .B1(new_n937), .B2(new_n932), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n943), .B1(new_n934), .B2(new_n1177), .ZN(new_n1178));
  OAI211_X1 g0978(.A(G330), .B(new_n1174), .C1(new_n1176), .C2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1174), .B1(new_n944), .B2(G330), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1170), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1174), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1109), .A2(new_n1175), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n934), .A2(new_n1177), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n943), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1184), .A2(KEYINPUT40), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1183), .B1(new_n1187), .B2(new_n1128), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1188), .A2(new_n957), .A3(new_n1179), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1000), .B1(new_n1182), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT121), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1183), .A2(new_n816), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n760), .B1(G50), .B2(new_n841), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n778), .A2(new_n1153), .B1(new_n770), .B2(new_n978), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G125), .B2(new_n847), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G132), .A2(new_n781), .B1(new_n774), .B2(new_n1162), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(new_n790), .C2(new_n324), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(G33), .A2(G41), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n775), .B2(new_n434), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n786), .B2(G124), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1199), .A2(new_n1200), .A3(new_n1203), .ZN(new_n1204));
  AOI211_X1 g1004(.A(G50), .B(new_n1201), .C1(new_n408), .C2(new_n556), .ZN(new_n1205));
  AOI211_X1 g1005(.A(G41), .B(new_n400), .C1(new_n786), .C2(G283), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n767), .A2(new_n512), .B1(new_n780), .B2(new_n224), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n778), .A2(new_n366), .B1(new_n770), .B2(new_n375), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n775), .A2(new_n222), .ZN(new_n1209));
  NOR4_X1   g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1053), .A4(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1206), .A2(new_n1210), .A3(new_n977), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT58), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1205), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1204), .B(new_n1213), .C1(new_n1212), .C2(new_n1211), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1194), .B1(new_n1214), .B2(new_n763), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1193), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1191), .A2(new_n1192), .A3(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1216), .ZN(new_n1218));
  OAI21_X1  g1018(.A(KEYINPUT121), .B1(new_n1190), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(new_n1140), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1221));
  OAI21_X1  g1021(.A(KEYINPUT122), .B1(new_n1221), .B2(new_n1118), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT122), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1133), .A2(new_n1223), .A3(new_n1138), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1222), .A2(new_n1224), .B1(new_n1189), .B2(new_n1182), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n711), .B1(new_n1225), .B2(KEYINPUT57), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1133), .A2(new_n1223), .A3(new_n1138), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1223), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1228));
  OAI21_X1  g1028(.A(KEYINPUT57), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1182), .A2(new_n1189), .A3(KEYINPUT123), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT123), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1188), .A2(new_n1231), .A3(new_n957), .A4(new_n1179), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1229), .A2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1220), .B1(new_n1226), .B2(new_n1234), .ZN(G375));
  NAND3_X1  g1035(.A1(new_n1126), .A2(new_n1118), .A3(new_n1130), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1236), .A2(new_n1139), .A3(new_n1018), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n793), .A2(G97), .B1(G303), .B2(new_n786), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n263), .B1(new_n776), .B2(G77), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n767), .A2(new_n983), .B1(new_n780), .B2(new_n512), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n778), .A2(new_n850), .B1(new_n770), .B2(new_n366), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1238), .A2(new_n1058), .A3(new_n1239), .A4(new_n1242), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n793), .A2(G159), .B1(G128), .B2(new_n786), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n789), .A2(G50), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n767), .A2(new_n1154), .B1(new_n778), .B2(new_n978), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G150), .B2(new_n848), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n408), .B(new_n1209), .C1(new_n781), .C2(new_n1162), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1244), .A2(new_n1245), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1243), .A2(new_n1249), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n760), .B1(G68), .B2(new_n841), .C1(new_n1250), .C2(new_n764), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n941), .B2(new_n816), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1137), .B2(new_n999), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1237), .A2(new_n1253), .ZN(G381));
  OR2_X1    g1054(.A1(G375), .A2(new_n1168), .ZN(new_n1255));
  OR4_X1    g1055(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1256));
  OR4_X1    g1056(.A1(G387), .A2(new_n1255), .A3(G381), .A4(new_n1256), .ZN(G407));
  OAI211_X1 g1057(.A(G407), .B(G213), .C1(G343), .C2(new_n1255), .ZN(G409));
  AND2_X1   g1058(.A1(new_n693), .A2(G213), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1182), .A2(new_n1189), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1018), .B(new_n1260), .C1(new_n1227), .C2(new_n1228), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(KEYINPUT124), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1230), .A2(new_n999), .A3(new_n1232), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1263), .A2(new_n1216), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT124), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1265), .A2(new_n1266), .A3(new_n1018), .A4(new_n1260), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1262), .A2(new_n1264), .A3(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1168), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(G378), .B(new_n1220), .C1(new_n1226), .C2(new_n1234), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1259), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT60), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1236), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(new_n711), .A3(new_n1139), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1236), .A2(new_n1273), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1253), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1277), .A2(new_n869), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n869), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1272), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT126), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1281), .A2(new_n1282), .A3(KEYINPUT62), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT61), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1259), .A2(G2897), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1280), .B(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1284), .B1(new_n1272), .B2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1280), .ZN(new_n1289));
  AOI211_X1 g1089(.A(new_n1259), .B(new_n1289), .C1(new_n1270), .C2(new_n1271), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1283), .A2(new_n1288), .A3(new_n1292), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(G393), .B(new_n825), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G390), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1294), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1103), .A2(new_n1105), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(G387), .A2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1035), .A2(new_n1295), .A3(new_n1297), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1293), .A2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1301), .B1(new_n1290), .B2(KEYINPUT63), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT63), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1281), .A2(new_n1304), .ZN(new_n1305));
  AND4_X1   g1105(.A1(KEYINPUT125), .A2(new_n1303), .A3(new_n1305), .A4(new_n1288), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT63), .B1(new_n1272), .B2(new_n1280), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1287), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT125), .B1(new_n1308), .B2(new_n1303), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1302), .B1(new_n1306), .B2(new_n1309), .ZN(G405));
  XOR2_X1   g1110(.A(new_n1280), .B(KEYINPUT127), .Z(new_n1311));
  AND2_X1   g1111(.A1(G375), .A2(new_n1269), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1271), .ZN(new_n1313));
  OR3_X1    g1113(.A1(new_n1311), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1311), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1301), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(new_n1316), .B(new_n1317), .ZN(G402));
endmodule


