//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT75), .Z(new_n188));
  INV_X1    g002(.A(KEYINPUT32), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  OR2_X1    g004(.A1(KEYINPUT70), .A2(G237), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT70), .A2(G237), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(G210), .A3(new_n194), .ZN(new_n195));
  XOR2_X1   g009(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n196));
  XNOR2_X1  g010(.A(new_n195), .B(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT26), .B(G101), .ZN(new_n198));
  XNOR2_X1  g012(.A(new_n197), .B(new_n198), .ZN(new_n199));
  OR2_X1    g013(.A1(KEYINPUT68), .A2(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT68), .A2(G119), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(G116), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G116), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G119), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT2), .B(G113), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n206), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(new_n202), .A3(new_n204), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT11), .ZN(new_n214));
  INV_X1    g028(.A(G137), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(G134), .ZN(new_n216));
  INV_X1    g030(.A(G134), .ZN(new_n217));
  OAI22_X1  g031(.A1(new_n217), .A2(G137), .B1(KEYINPUT64), .B2(KEYINPUT11), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G131), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n221), .B1(new_n215), .B2(G134), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  AND4_X1   g037(.A1(new_n212), .A2(new_n219), .A3(new_n220), .A4(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n222), .B1(new_n218), .B2(new_n216), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n212), .B1(new_n225), .B2(new_n220), .ZN(new_n226));
  OAI22_X1  g040(.A1(new_n224), .A2(new_n226), .B1(new_n220), .B2(new_n225), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n228));
  XNOR2_X1  g042(.A(G143), .B(G146), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(KEYINPUT0), .A3(G128), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT0), .B(G128), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n227), .A2(new_n228), .A3(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n225), .A2(new_n220), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n219), .A2(new_n220), .A3(new_n223), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT65), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n225), .A2(new_n212), .A3(new_n220), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n235), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT66), .B1(new_n239), .B2(new_n232), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n234), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n215), .A2(G134), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n217), .A2(G137), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n220), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G143), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT1), .B1(new_n247), .B2(G146), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(G146), .ZN(new_n249));
  INV_X1    g063(.A(G146), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(G143), .ZN(new_n251));
  OAI211_X1 g065(.A(G128), .B(new_n248), .C1(new_n249), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n247), .A2(G146), .ZN(new_n254));
  INV_X1    g068(.A(G128), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n253), .B(new_n254), .C1(KEYINPUT1), .C2(new_n255), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n246), .B(new_n257), .C1(new_n224), .C2(new_n226), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n258), .B(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n211), .B1(new_n242), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n227), .A2(new_n233), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n245), .B1(new_n237), .B2(new_n238), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n252), .A2(KEYINPUT69), .A3(new_n256), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT69), .B1(new_n252), .B2(new_n256), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n262), .A2(new_n267), .A3(new_n211), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT28), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n262), .A2(new_n267), .A3(KEYINPUT28), .A4(new_n211), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n199), .B1(new_n261), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT73), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n275), .B(new_n199), .C1(new_n261), .C2(new_n272), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT30), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n258), .A2(new_n259), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT67), .B1(new_n263), .B2(new_n257), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n277), .B1(new_n280), .B2(new_n241), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n262), .A2(new_n267), .A3(KEYINPUT30), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n210), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n199), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n283), .A2(KEYINPUT72), .A3(new_n268), .A4(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT31), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n286), .A2(KEYINPUT72), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n287), .A2(KEYINPUT31), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n268), .ZN(new_n290));
  INV_X1    g104(.A(new_n282), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n240), .B(new_n234), .C1(new_n278), .C2(new_n279), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n291), .B1(new_n292), .B2(new_n277), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n290), .B1(new_n293), .B2(new_n210), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n294), .A2(KEYINPUT72), .A3(KEYINPUT31), .A4(new_n284), .ZN(new_n295));
  AOI221_X4 g109(.A(KEYINPUT74), .B1(new_n274), .B2(new_n276), .C1(new_n289), .C2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n289), .A2(new_n295), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n274), .A2(new_n276), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n190), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G472), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT78), .B(G902), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  XOR2_X1   g118(.A(new_n270), .B(KEYINPUT77), .Z(new_n305));
  INV_X1    g119(.A(KEYINPUT76), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n268), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n262), .A2(new_n267), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n210), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n307), .B(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n305), .B1(new_n310), .B2(KEYINPUT28), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n284), .A2(KEYINPUT29), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n304), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OR2_X1    g127(.A1(new_n294), .A2(new_n284), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n261), .A2(new_n272), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT29), .B1(new_n315), .B2(new_n284), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n302), .B1(new_n313), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n298), .A2(new_n299), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT74), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n298), .A2(new_n299), .A3(new_n297), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n188), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n301), .B(new_n319), .C1(new_n323), .C2(KEYINPUT32), .ZN(new_n324));
  INV_X1    g138(.A(G217), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(new_n303), .B2(G234), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(G140), .ZN(new_n329));
  XNOR2_X1  g143(.A(G125), .B(G140), .ZN(new_n330));
  MUX2_X1   g144(.A(new_n329), .B(new_n330), .S(KEYINPUT16), .Z(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(new_n250), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n200), .A2(G128), .A3(new_n201), .ZN(new_n333));
  INV_X1    g147(.A(G119), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n333), .B1(new_n334), .B2(G128), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT24), .B(G110), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n200), .A2(new_n201), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n255), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n338), .A2(KEYINPUT79), .B1(KEYINPUT23), .B2(new_n333), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n339), .B1(KEYINPUT79), .B2(new_n338), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n255), .A2(KEYINPUT23), .A3(G119), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G110), .ZN(new_n343));
  OAI221_X1 g157(.A(new_n332), .B1(new_n335), .B2(new_n336), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(KEYINPUT80), .ZN(new_n346));
  XOR2_X1   g160(.A(KEYINPUT22), .B(G137), .Z(new_n347));
  XNOR2_X1  g161(.A(new_n346), .B(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n342), .A2(new_n343), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n335), .A2(new_n336), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n330), .A2(new_n250), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n352), .B1(new_n331), .B2(new_n250), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n344), .B(new_n348), .C1(new_n351), .C2(new_n353), .ZN(new_n354));
  XOR2_X1   g168(.A(new_n348), .B(KEYINPUT81), .Z(new_n355));
  AOI21_X1  g169(.A(new_n353), .B1(new_n349), .B2(new_n350), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n342), .A2(new_n343), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n332), .B1(new_n335), .B2(new_n336), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n355), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n354), .A2(new_n360), .A3(new_n303), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT82), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT25), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n327), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT25), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n326), .A2(G902), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n354), .A2(new_n360), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n365), .A2(new_n366), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G902), .ZN(new_n371));
  AND2_X1   g185(.A1(KEYINPUT70), .A2(G237), .ZN(new_n372));
  NOR2_X1   g186(.A1(KEYINPUT70), .A2(G237), .ZN(new_n373));
  OAI211_X1 g187(.A(G214), .B(new_n194), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT91), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n193), .A2(KEYINPUT91), .A3(G214), .A4(new_n194), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(new_n377), .A3(new_n247), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT92), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(G143), .B1(new_n374), .B2(new_n375), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(KEYINPUT92), .A3(new_n377), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  OR3_X1    g197(.A1(new_n374), .A2(KEYINPUT93), .A3(new_n247), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT93), .B1(new_n374), .B2(new_n247), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n220), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n332), .B1(new_n387), .B2(KEYINPUT17), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n381), .A2(KEYINPUT92), .A3(new_n377), .ZN(new_n389));
  AOI21_X1  g203(.A(KEYINPUT92), .B1(new_n381), .B2(new_n377), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n386), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G131), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT17), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n220), .B(new_n386), .C1(new_n389), .C2(new_n390), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n388), .A2(new_n395), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n380), .A2(new_n382), .B1(new_n385), .B2(new_n384), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT94), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT18), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n397), .B(new_n398), .C1(new_n399), .C2(new_n220), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n399), .B(new_n386), .C1(new_n389), .C2(new_n390), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n394), .A2(new_n401), .A3(KEYINPUT94), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n391), .A2(KEYINPUT18), .A3(G131), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n330), .B(new_n250), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n400), .A2(new_n402), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(G113), .B(G122), .ZN(new_n406));
  INV_X1    g220(.A(G104), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n406), .B(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n396), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n408), .B1(new_n396), .B2(new_n405), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n371), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G475), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT20), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n331), .A2(new_n250), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n330), .B(KEYINPUT19), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n415), .B1(new_n250), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n394), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n417), .B1(new_n387), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n405), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n408), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n409), .ZN(new_n423));
  NOR2_X1   g237(.A1(G475), .A2(G902), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n414), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n424), .ZN(new_n426));
  AOI211_X1 g240(.A(KEYINPUT20), .B(new_n426), .C1(new_n422), .C2(new_n409), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n413), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(G234), .A2(G237), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n429), .A2(G952), .A3(new_n194), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n304), .A2(G953), .A3(new_n429), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(G898), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n247), .A2(G128), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n247), .A2(G128), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT13), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n437), .B(KEYINPUT95), .C1(new_n436), .C2(new_n434), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT95), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n439), .B(new_n434), .C1(new_n435), .C2(new_n436), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n438), .A2(G134), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT96), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT96), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n438), .A2(new_n443), .A3(G134), .A4(new_n440), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n435), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(new_n217), .A3(new_n434), .ZN(new_n447));
  OR2_X1    g261(.A1(new_n203), .A2(G122), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n203), .A2(G122), .ZN(new_n449));
  INV_X1    g263(.A(G107), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n450), .B1(new_n448), .B2(new_n449), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n447), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n445), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT97), .B1(new_n449), .B2(KEYINPUT14), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT97), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT14), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n457), .A2(new_n458), .A3(new_n203), .A4(G122), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n449), .A2(KEYINPUT14), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n456), .A2(new_n448), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G107), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT98), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT98), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n461), .A2(new_n464), .A3(G107), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n447), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n217), .B1(new_n446), .B2(new_n434), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(new_n451), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT9), .B(G234), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n472), .A2(new_n325), .A3(G953), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n455), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n473), .ZN(new_n475));
  AOI211_X1 g289(.A(new_n451), .B(new_n469), .C1(new_n463), .C2(new_n465), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n453), .B1(new_n442), .B2(new_n444), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n303), .ZN(new_n480));
  INV_X1    g294(.A(G478), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n481), .A2(KEYINPUT15), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n480), .B(new_n482), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n428), .A2(new_n433), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(G214), .B1(G237), .B2(G902), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n485), .B(KEYINPUT88), .Z(new_n486));
  OAI21_X1  g300(.A(G210), .B1(G237), .B2(G902), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(G110), .B(G122), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(KEYINPUT8), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n202), .A2(KEYINPUT5), .A3(new_n204), .ZN(new_n491));
  OAI21_X1  g305(.A(G113), .B1(new_n202), .B2(KEYINPUT5), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n209), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT83), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n407), .ZN(new_n495));
  NAND2_X1  g309(.A1(KEYINPUT83), .A2(G104), .ZN(new_n496));
  AOI21_X1  g310(.A(G107), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n450), .A2(G104), .ZN(new_n498));
  OAI21_X1  g312(.A(G101), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n407), .A2(KEYINPUT3), .A3(G107), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT3), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n501), .B1(new_n497), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n495), .A2(G107), .A3(new_n496), .ZN(new_n504));
  INV_X1    g318(.A(G101), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n499), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n493), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(KEYINPUT89), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT85), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g325(.A(KEYINPUT85), .B(new_n499), .C1(new_n503), .C2(new_n506), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n493), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n490), .B1(new_n509), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n493), .ZN(new_n515));
  INV_X1    g329(.A(new_n512), .ZN(new_n516));
  AND2_X1   g330(.A1(KEYINPUT83), .A2(G104), .ZN(new_n517));
  NOR2_X1   g331(.A1(KEYINPUT83), .A2(G104), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(G101), .B1(new_n519), .B2(G107), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n450), .B1(new_n517), .B2(new_n518), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT3), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n520), .A2(new_n522), .A3(new_n501), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT85), .B1(new_n523), .B2(new_n499), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n515), .B1(new_n516), .B2(new_n524), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n501), .B(new_n504), .C1(new_n497), .C2(new_n502), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT4), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(new_n527), .A3(G101), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT4), .B1(new_n503), .B2(new_n506), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n500), .B1(new_n521), .B2(KEYINPUT3), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n505), .B1(new_n530), .B2(new_n504), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n210), .B(new_n528), .C1(new_n529), .C2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n525), .A2(new_n532), .A3(new_n489), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n229), .A2(new_n231), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n328), .B1(new_n534), .B2(new_n230), .ZN(new_n535));
  AOI21_X1  g349(.A(G125), .B1(new_n252), .B2(new_n256), .ZN(new_n536));
  OAI211_X1 g350(.A(G224), .B(new_n194), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n232), .A2(G125), .ZN(new_n538));
  INV_X1    g352(.A(new_n536), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n194), .A2(G224), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT7), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n537), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n538), .A2(new_n539), .A3(new_n542), .A4(new_n540), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n514), .A2(new_n533), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT90), .B1(new_n547), .B2(new_n371), .ZN(new_n548));
  INV_X1    g362(.A(new_n490), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT89), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n508), .B(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n549), .B1(new_n551), .B2(new_n525), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n546), .A2(new_n533), .ZN(new_n553));
  OAI211_X1 g367(.A(KEYINPUT90), .B(new_n371), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n489), .ZN(new_n555));
  INV_X1    g369(.A(new_n532), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n555), .B1(new_n556), .B2(new_n513), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(KEYINPUT6), .A3(new_n533), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n537), .A2(new_n541), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT6), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n560), .B(new_n555), .C1(new_n556), .C2(new_n513), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n554), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n488), .B1(new_n548), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n371), .B1(new_n552), .B2(new_n553), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT90), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n567), .A2(new_n487), .A3(new_n562), .A4(new_n554), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n486), .B1(new_n564), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(G221), .B1(new_n472), .B2(G902), .ZN(new_n570));
  INV_X1    g384(.A(G469), .ZN(new_n571));
  XNOR2_X1  g385(.A(G110), .B(G140), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n194), .A2(G227), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT10), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n264), .A2(new_n265), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n516), .B2(new_n524), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT86), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n577), .B(KEYINPUT86), .C1(new_n516), .C2(new_n524), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n233), .B(new_n528), .C1(new_n529), .C2(new_n531), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n523), .A2(new_n257), .A3(new_n499), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT84), .B1(new_n585), .B2(new_n576), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(KEYINPUT84), .A3(new_n576), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n584), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n582), .A2(new_n589), .A3(new_n239), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT87), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n582), .A2(new_n589), .A3(KEYINPUT87), .A4(new_n239), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n582), .A2(new_n589), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n227), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n575), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n252), .A2(new_n256), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n511), .A2(new_n598), .A3(new_n512), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n585), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT12), .B1(new_n600), .B2(new_n227), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT12), .ZN(new_n602));
  AOI211_X1 g416(.A(new_n602), .B(new_n239), .C1(new_n599), .C2(new_n585), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  AOI211_X1 g418(.A(new_n574), .B(new_n604), .C1(new_n592), .C2(new_n593), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n571), .B(new_n303), .C1(new_n597), .C2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n571), .A2(new_n371), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n585), .A2(KEYINPUT84), .A3(new_n576), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n583), .B1(new_n609), .B2(new_n586), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n580), .B2(new_n581), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT87), .B1(new_n611), .B2(new_n239), .ZN(new_n612));
  INV_X1    g426(.A(new_n593), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n596), .B(new_n575), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n604), .B1(new_n592), .B2(new_n593), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n614), .B(G469), .C1(new_n575), .C2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n606), .A2(new_n608), .A3(new_n616), .ZN(new_n617));
  AND4_X1   g431(.A1(new_n484), .A2(new_n569), .A3(new_n570), .A4(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n324), .A2(new_n370), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G101), .ZN(G3));
  OAI21_X1  g434(.A(new_n303), .B1(new_n296), .B2(new_n300), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n321), .A2(new_n322), .ZN(new_n622));
  INV_X1    g436(.A(new_n188), .ZN(new_n623));
  AOI22_X1  g437(.A1(G472), .A2(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n570), .ZN(new_n625));
  INV_X1    g439(.A(new_n604), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n594), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n574), .B1(new_n592), .B2(new_n593), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n627), .A2(new_n574), .B1(new_n628), .B2(new_n596), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n607), .B1(new_n629), .B2(G469), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n625), .B1(new_n630), .B2(new_n606), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n624), .A2(new_n370), .A3(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n633), .B(new_n488), .C1(new_n548), .C2(new_n563), .ZN(new_n634));
  INV_X1    g448(.A(new_n486), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n433), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n564), .A2(KEYINPUT99), .A3(new_n568), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n479), .A2(new_n481), .A3(new_n303), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n476), .A2(new_n477), .A3(new_n475), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n473), .B1(new_n455), .B2(new_n471), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT33), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n474), .A2(new_n478), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n304), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n640), .B1(new_n646), .B2(new_n481), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT100), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT100), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n640), .B(new_n649), .C1(new_n646), .C2(new_n481), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n428), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n639), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n632), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT34), .B(G104), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G6));
  XOR2_X1   g471(.A(new_n433), .B(KEYINPUT101), .Z(new_n658));
  NAND4_X1  g472(.A1(new_n638), .A2(new_n635), .A3(new_n634), .A4(new_n658), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n413), .B(new_n483), .C1(new_n425), .C2(new_n427), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n632), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT35), .B(G107), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G9));
  NAND2_X1  g479(.A1(new_n365), .A2(new_n366), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n356), .A2(new_n359), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n355), .A2(KEYINPUT36), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n667), .B(new_n668), .Z(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n367), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n484), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n624), .A2(new_n569), .A3(new_n631), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT37), .B(G110), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G12));
  NAND3_X1  g492(.A1(new_n617), .A2(new_n671), .A3(new_n570), .ZN(new_n679));
  INV_X1    g493(.A(G900), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n430), .B1(new_n431), .B2(new_n680), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n679), .A2(new_n660), .A3(new_n681), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n638), .A2(new_n635), .A3(new_n634), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n682), .A2(new_n324), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G128), .ZN(G30));
  XOR2_X1   g499(.A(new_n681), .B(KEYINPUT39), .Z(new_n686));
  NAND2_X1  g500(.A1(new_n631), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT40), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n631), .A2(KEYINPUT40), .A3(new_n686), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n294), .A2(new_n284), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n694), .B1(new_n199), .B2(new_n310), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n695), .B2(G902), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n301), .B(new_n696), .C1(new_n323), .C2(KEYINPUT32), .ZN(new_n697));
  AOI22_X1  g511(.A1(new_n365), .A2(new_n366), .B1(new_n367), .B2(new_n669), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n564), .A2(new_n568), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT38), .ZN(new_n701));
  INV_X1    g515(.A(new_n483), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n423), .A2(new_n424), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT20), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n423), .A2(new_n414), .A3(new_n424), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n702), .B1(new_n706), .B2(new_n413), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n701), .A2(new_n635), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n689), .A2(KEYINPUT104), .A3(new_n690), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n693), .A2(new_n699), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G143), .ZN(G45));
  INV_X1    g525(.A(new_n681), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n428), .A2(new_n651), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n679), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n324), .A2(new_n683), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  OAI21_X1  g530(.A(new_n596), .B1(new_n612), .B2(new_n613), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n717), .A2(new_n574), .B1(new_n628), .B2(new_n626), .ZN(new_n718));
  OAI21_X1  g532(.A(G469), .B1(new_n718), .B2(new_n304), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n570), .A3(new_n606), .ZN(new_n720));
  INV_X1    g534(.A(new_n370), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n324), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n654), .ZN(new_n724));
  XOR2_X1   g538(.A(KEYINPUT41), .B(G113), .Z(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NOR2_X1   g540(.A1(new_n723), .A2(new_n662), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n203), .ZN(G18));
  INV_X1    g542(.A(new_n606), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n575), .B(new_n626), .C1(new_n612), .C2(new_n613), .ZN(new_n730));
  AOI22_X1  g544(.A1(new_n592), .A2(new_n593), .B1(new_n227), .B2(new_n595), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n730), .B1(new_n731), .B2(new_n575), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n571), .B1(new_n732), .B2(new_n303), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n734), .A2(KEYINPUT105), .A3(new_n570), .A4(new_n683), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n636), .A2(new_n638), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n736), .B1(new_n720), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n324), .A3(new_n673), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G119), .ZN(G21));
  OR2_X1    g555(.A1(new_n311), .A2(new_n284), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n188), .B1(new_n742), .B2(new_n298), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n721), .B(new_n743), .C1(new_n621), .C2(G472), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n428), .A2(new_n483), .ZN(new_n745));
  INV_X1    g559(.A(new_n658), .ZN(new_n746));
  NOR4_X1   g560(.A1(new_n720), .A2(new_n737), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G122), .ZN(G24));
  AOI211_X1 g563(.A(new_n698), .B(new_n743), .C1(new_n621), .C2(G472), .ZN(new_n750));
  INV_X1    g564(.A(new_n713), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n739), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(KEYINPUT106), .B(G125), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(G27));
  AOI21_X1  g568(.A(new_n318), .B1(new_n622), .B2(new_n190), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n296), .A2(new_n300), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n189), .B1(new_n756), .B2(new_n188), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n721), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n616), .A2(new_n608), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n759), .B1(new_n729), .B2(new_n760), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n700), .A2(new_n486), .A3(new_n625), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n630), .A2(KEYINPUT107), .A3(new_n606), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n713), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(KEYINPUT42), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n758), .A2(new_n765), .A3(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n766), .A2(KEYINPUT42), .ZN(new_n771));
  AOI22_X1  g585(.A1(new_n758), .A2(new_n765), .B1(new_n771), .B2(new_n768), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(new_n220), .ZN(G33));
  NOR2_X1   g588(.A1(new_n660), .A2(new_n681), .ZN(new_n775));
  AND4_X1   g589(.A1(new_n775), .A2(new_n761), .A3(new_n762), .A4(new_n763), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(new_n324), .A3(new_n370), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  INV_X1    g592(.A(new_n624), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n428), .B1(new_n648), .B2(new_n650), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT43), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n779), .A2(new_n781), .A3(new_n671), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n700), .A2(new_n486), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n782), .A2(new_n783), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n629), .A2(KEYINPUT45), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n629), .A2(KEYINPUT45), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(G469), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n608), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT110), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n790), .A2(KEYINPUT46), .A3(new_n608), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT109), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n796), .A3(new_n606), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT110), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n791), .A2(new_n798), .A3(new_n792), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n794), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n796), .B1(new_n795), .B2(new_n606), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n570), .B(new_n686), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n787), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(KEYINPUT111), .B(G137), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n803), .B(new_n804), .ZN(G39));
  OAI21_X1  g619(.A(new_n570), .B1(new_n800), .B2(new_n801), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT47), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(KEYINPUT47), .B(new_n570), .C1(new_n800), .C2(new_n801), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n785), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n324), .A2(new_n370), .A3(new_n713), .A4(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT112), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G140), .ZN(G42));
  NOR2_X1   g629(.A1(new_n697), .A2(new_n721), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n701), .A2(new_n486), .A3(new_n625), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n734), .B(KEYINPUT49), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n816), .A2(new_n780), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n734), .A2(new_n486), .A3(new_n570), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n701), .B1(new_n821), .B2(KEYINPUT116), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n822), .B1(KEYINPUT116), .B2(new_n821), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n744), .A2(new_n781), .A3(new_n430), .ZN(new_n824));
  OR4_X1    g638(.A1(new_n820), .A2(new_n823), .A3(new_n824), .A4(KEYINPUT50), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n734), .A2(new_n430), .A3(new_n762), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n781), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT118), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n781), .A2(new_n829), .A3(new_n826), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n816), .A2(new_n826), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n428), .A2(new_n651), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n831), .A2(new_n750), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(KEYINPUT117), .B(KEYINPUT50), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(new_n823), .B2(new_n824), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n825), .A2(new_n835), .A3(KEYINPUT51), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n734), .A2(new_n625), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n808), .A2(new_n809), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n824), .A2(new_n811), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI211_X1 g656(.A(G952), .B(new_n194), .C1(new_n832), .C2(new_n652), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n824), .B1(new_n738), .B2(new_n735), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT48), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n846), .B1(new_n831), .B2(new_n758), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n324), .A2(new_n370), .ZN(new_n848));
  AOI211_X1 g662(.A(KEYINPUT48), .B(new_n848), .C1(new_n828), .C2(new_n830), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n845), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n842), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n825), .A2(new_n835), .A3(new_n837), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n808), .A2(new_n857), .A3(new_n809), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n856), .A2(new_n858), .A3(new_n839), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n855), .B1(new_n859), .B2(new_n841), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n854), .B1(new_n860), .B2(KEYINPUT51), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n617), .A2(new_n671), .A3(new_n570), .A4(new_n785), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT114), .ZN(new_n863));
  NOR4_X1   g677(.A1(new_n428), .A2(new_n863), .A3(new_n483), .A4(new_n681), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n428), .A2(new_n483), .A3(new_n681), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n866), .A2(KEYINPUT114), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n324), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n758), .A2(new_n776), .B1(new_n765), .B2(new_n750), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n868), .B(new_n869), .C1(new_n770), .C2(new_n772), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n674), .A2(new_n619), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT32), .B1(new_n622), .B2(new_n623), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n301), .A2(new_n319), .ZN(new_n873));
  OAI221_X1 g687(.A(new_n722), .B1(new_n653), .B2(new_n661), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n672), .B1(new_n755), .B2(new_n757), .ZN(new_n875));
  AOI22_X1  g689(.A1(new_n875), .A2(new_n739), .B1(new_n744), .B2(new_n747), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n569), .A2(new_n658), .ZN(new_n877));
  AOI22_X1  g691(.A1(KEYINPUT113), .A2(new_n660), .B1(new_n428), .B2(new_n651), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n660), .A2(KEYINPUT113), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n624), .A2(new_n880), .A3(new_n370), .A4(new_n631), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n871), .A2(new_n874), .A3(new_n876), .A4(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n870), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n713), .B1(new_n735), .B2(new_n738), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n737), .B1(new_n755), .B2(new_n757), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n750), .A2(new_n884), .B1(new_n885), .B2(new_n682), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT52), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n761), .A2(new_n763), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n681), .A2(new_n625), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n683), .A2(new_n707), .A3(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n697), .A2(new_n698), .A3(new_n888), .A4(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n886), .A2(new_n887), .A3(new_n715), .A4(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT53), .ZN(new_n893));
  INV_X1    g707(.A(new_n886), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n894), .B2(KEYINPUT52), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n752), .A2(new_n891), .A3(new_n684), .A4(new_n715), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT52), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n883), .A2(new_n892), .A3(new_n895), .A4(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT54), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n743), .B1(new_n621), .B2(G472), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n900), .A2(new_n671), .A3(new_n751), .A4(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n777), .A2(new_n902), .A3(new_n868), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n768), .A2(new_n771), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n900), .A2(new_n751), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n904), .B1(new_n848), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n903), .B1(new_n906), .B2(new_n769), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n740), .A2(new_n874), .A3(new_n748), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n881), .A2(new_n674), .A3(new_n619), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n907), .A2(new_n892), .A3(new_n897), .A4(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n893), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n898), .A2(new_n899), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT53), .B1(new_n894), .B2(KEYINPUT52), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n899), .B1(new_n916), .B2(new_n912), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n861), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(G952), .A2(G953), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n819), .B1(new_n920), .B2(new_n921), .ZN(G75));
  NAND2_X1  g736(.A1(new_n558), .A2(new_n561), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(new_n559), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n911), .A2(new_n893), .ZN(new_n926));
  INV_X1    g740(.A(new_n895), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n911), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n304), .B(new_n488), .C1(new_n926), .C2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT56), .ZN(new_n930));
  XNOR2_X1  g744(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n929), .B2(new_n930), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n925), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n194), .A2(G952), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT121), .Z(new_n937));
  AOI211_X1 g751(.A(new_n303), .B(new_n487), .C1(new_n898), .C2(new_n912), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n931), .B1(new_n938), .B2(KEYINPUT56), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n939), .A2(new_n924), .A3(new_n940), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n935), .A2(new_n937), .A3(new_n941), .ZN(G51));
  INV_X1    g756(.A(new_n937), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n304), .B1(new_n926), .B2(new_n928), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n944), .A2(new_n790), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT54), .B1(new_n926), .B2(new_n928), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n913), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n607), .B(KEYINPUT57), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n718), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT122), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n945), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n948), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n946), .B2(new_n913), .ZN(new_n953));
  OAI21_X1  g767(.A(KEYINPUT122), .B1(new_n953), .B2(new_n718), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n943), .B1(new_n951), .B2(new_n954), .ZN(G54));
  NAND2_X1  g769(.A1(KEYINPUT58), .A2(G475), .ZN(new_n956));
  OR3_X1    g770(.A1(new_n944), .A2(new_n423), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n423), .B1(new_n944), .B2(new_n956), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n943), .B1(new_n957), .B2(new_n958), .ZN(G60));
  NAND2_X1  g773(.A1(new_n643), .A2(new_n645), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  XOR2_X1   g775(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n962));
  NOR2_X1   g776(.A1(new_n481), .A2(new_n371), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n961), .B1(new_n918), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT124), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n961), .A2(new_n964), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n946), .B2(new_n913), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n966), .B1(new_n969), .B2(new_n943), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n965), .A2(new_n970), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n969), .A2(new_n966), .A3(new_n943), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n971), .A2(new_n972), .ZN(G63));
  INV_X1    g787(.A(KEYINPUT61), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n974), .A2(KEYINPUT125), .ZN(new_n975));
  NAND2_X1  g789(.A1(G217), .A2(G902), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT60), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n898), .B2(new_n912), .ZN(new_n978));
  AOI211_X1 g792(.A(new_n943), .B(new_n975), .C1(new_n978), .C2(new_n669), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n974), .A2(KEYINPUT125), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n978), .A2(new_n369), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n979), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n981), .B1(new_n979), .B2(new_n982), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(G66));
  INV_X1    g799(.A(G224), .ZN(new_n986));
  OAI21_X1  g800(.A(G953), .B1(new_n432), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(new_n910), .B2(G953), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n923), .B1(G898), .B2(new_n194), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT126), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n988), .B(new_n990), .ZN(G69));
  AOI21_X1  g805(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n878), .A2(new_n879), .ZN(new_n993));
  NOR4_X1   g807(.A1(new_n848), .A2(new_n993), .A3(new_n687), .A4(new_n811), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT127), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n803), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n814), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n886), .A2(new_n715), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n710), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT62), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n999), .A2(KEYINPUT62), .A3(new_n710), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(G953), .B1(new_n998), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n293), .B(new_n416), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(new_n773), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n1008), .A2(new_n777), .A3(new_n999), .ZN(new_n1009));
  INV_X1    g823(.A(new_n802), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n1010), .A2(new_n758), .A3(new_n683), .A4(new_n707), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1009), .B(new_n1011), .C1(new_n802), .C2(new_n787), .ZN(new_n1012));
  INV_X1    g826(.A(new_n814), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n1012), .A2(G953), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1006), .B1(new_n680), .B2(new_n194), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n992), .B1(new_n1007), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(new_n992), .ZN(new_n1018));
  OAI221_X1 g832(.A(new_n1018), .B1(new_n1014), .B2(new_n1015), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1017), .A2(new_n1019), .ZN(G72));
  INV_X1    g834(.A(new_n694), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(new_n314), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1004), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n284), .B1(new_n997), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n199), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1024), .A2(new_n1025), .A3(new_n910), .ZN(new_n1026));
  NAND2_X1  g840(.A1(G472), .A2(G902), .ZN(new_n1027));
  XOR2_X1   g841(.A(new_n1027), .B(KEYINPUT63), .Z(new_n1028));
  AOI21_X1  g842(.A(new_n1022), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1022), .A2(new_n1028), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1030), .B1(new_n916), .B2(new_n912), .ZN(new_n1031));
  NOR3_X1   g845(.A1(new_n1029), .A2(new_n943), .A3(new_n1031), .ZN(G57));
endmodule


