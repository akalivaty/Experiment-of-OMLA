//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  NAND3_X1  g0006(.A1(new_n201), .A2(KEYINPUT64), .A3(new_n202), .ZN(new_n207));
  AND3_X1   g0007(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  AND2_X1   g0013(.A1(G107), .A2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n215), .A2(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n214), .B(new_n219), .C1(G68), .C2(G238), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G116), .A2(G270), .ZN(new_n221));
  AND2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G226), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n222), .B1(new_n202), .B2(new_n223), .C1(new_n206), .C2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G58), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n210), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(G50), .B1(G58), .B2(G68), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n213), .B(new_n230), .C1(new_n233), .C2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT65), .B(G264), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n202), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n226), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  XOR2_X1   g0052(.A(KEYINPUT8), .B(G58), .Z(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n253), .A2(new_n254), .B1(G20), .B2(G77), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n232), .A2(G33), .ZN(new_n256));
  XOR2_X1   g0056(.A(KEYINPUT15), .B(G87), .Z(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n255), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n231), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n259), .A2(new_n261), .B1(G77), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n263), .A2(G13), .A3(G20), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(G77), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT68), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT69), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n267), .A2(KEYINPUT69), .A3(new_n270), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT3), .B(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G238), .A2(G1698), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n276), .B(new_n277), .C1(new_n227), .C2(G1698), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n278), .B(new_n281), .C1(G107), .C2(new_n276), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n283));
  INV_X1    g0083(.A(G274), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n280), .A2(new_n283), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n282), .B(new_n286), .C1(new_n224), .C2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G190), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n290), .B1(G200), .B2(new_n288), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n275), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n273), .A2(new_n274), .ZN(new_n293));
  INV_X1    g0093(.A(G169), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n288), .A2(G179), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n254), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n299), .A2(new_n202), .B1(new_n232), .B2(G68), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n256), .A2(new_n206), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n261), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  XOR2_X1   g0102(.A(new_n302), .B(KEYINPUT11), .Z(new_n303));
  INV_X1    g0103(.A(KEYINPUT12), .ZN(new_n304));
  INV_X1    g0104(.A(new_n268), .ZN(new_n305));
  INV_X1    g0105(.A(G68), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n268), .A2(KEYINPUT12), .A3(G68), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n307), .A2(new_n308), .B1(new_n265), .B2(new_n306), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(G226), .A2(G1698), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n227), .B2(G1698), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n276), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G33), .A2(G97), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n280), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT70), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n315), .B(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT13), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n286), .A2(KEYINPUT71), .ZN(new_n319));
  INV_X1    g0119(.A(new_n287), .ZN(new_n320));
  AOI22_X1  g0120(.A1(G238), .A2(new_n320), .B1(new_n286), .B2(KEYINPUT71), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n317), .A2(new_n318), .A3(new_n319), .A4(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n315), .A2(new_n316), .ZN(new_n323));
  AOI211_X1 g0123(.A(KEYINPUT70), .B(new_n280), .C1(new_n313), .C2(new_n314), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n319), .B(new_n321), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT13), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n310), .B1(new_n327), .B2(new_n289), .ZN(new_n328));
  INV_X1    g0128(.A(G200), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n322), .B2(new_n326), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT14), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(new_n327), .B2(G169), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  AOI211_X1 g0134(.A(KEYINPUT14), .B(new_n294), .C1(new_n322), .C2(new_n326), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n327), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n334), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n310), .ZN(new_n341));
  AOI211_X1 g0141(.A(new_n298), .B(new_n331), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT77), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n268), .A2(G50), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n265), .A2(new_n202), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n232), .B1(new_n205), .B2(new_n207), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT8), .B(G58), .ZN(new_n347));
  INV_X1    g0147(.A(G150), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n347), .A2(new_n256), .B1(new_n348), .B2(new_n299), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n261), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  OR2_X1    g0150(.A1(new_n350), .A2(KEYINPUT67), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(KEYINPUT67), .ZN(new_n352));
  AOI211_X1 g0152(.A(new_n344), .B(new_n345), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G1698), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G222), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT66), .B(G223), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n276), .B(new_n355), .C1(new_n356), .C2(new_n354), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n357), .B(new_n281), .C1(G77), .C2(new_n276), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n320), .A2(G226), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(new_n286), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n294), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(G179), .B2(new_n360), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n353), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(G200), .ZN(new_n364));
  INV_X1    g0164(.A(new_n360), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G190), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n344), .B1(new_n351), .B2(new_n352), .ZN(new_n367));
  INV_X1    g0167(.A(new_n345), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT9), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n364), .B(new_n366), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n353), .A2(KEYINPUT9), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT10), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n353), .A2(KEYINPUT9), .B1(G190), .B2(new_n365), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT10), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n369), .A2(new_n370), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .A4(new_n364), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n363), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT74), .ZN(new_n379));
  INV_X1    g0179(.A(G33), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT3), .ZN(new_n381));
  OR2_X1    g0181(.A1(G223), .A2(G1698), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT3), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G33), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n223), .A2(G1698), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n381), .A2(new_n382), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G87), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n285), .B1(new_n388), .B2(new_n281), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n280), .A2(G232), .A3(new_n283), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n294), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n280), .B1(new_n386), .B2(new_n387), .ZN(new_n393));
  NOR4_X1   g0193(.A1(new_n393), .A2(new_n337), .A3(new_n390), .A4(new_n285), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT16), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n383), .A2(KEYINPUT72), .A3(G33), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n381), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT72), .B1(new_n383), .B2(G33), .ZN(new_n399));
  OAI211_X1 g0199(.A(KEYINPUT7), .B(new_n232), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n276), .B2(G20), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n306), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n226), .A2(new_n306), .ZN(new_n404));
  OAI21_X1  g0204(.A(G20), .B1(new_n404), .B2(new_n201), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n254), .A2(G159), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n396), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n381), .A2(new_n384), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(KEYINPUT7), .A3(new_n232), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n402), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G68), .ZN(new_n412));
  INV_X1    g0212(.A(new_n407), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(KEYINPUT16), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n408), .A2(new_n414), .A3(new_n261), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n265), .A2(new_n253), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n347), .A2(new_n268), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n395), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n379), .B1(new_n419), .B2(KEYINPUT18), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT18), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n407), .B1(new_n411), .B2(G68), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n262), .B1(new_n422), .B2(KEYINPUT16), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n423), .A2(new_n408), .B1(new_n416), .B2(new_n417), .ZN(new_n424));
  OAI211_X1 g0224(.A(KEYINPUT74), .B(new_n421), .C1(new_n424), .C2(new_n395), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT73), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n419), .B2(KEYINPUT18), .ZN(new_n428));
  NOR4_X1   g0228(.A1(new_n424), .A2(KEYINPUT73), .A3(new_n395), .A4(new_n421), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n393), .A2(new_n285), .A3(new_n390), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G190), .ZN(new_n432));
  OR2_X1    g0232(.A1(new_n431), .A2(new_n329), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n415), .A2(new_n432), .A3(new_n418), .A4(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT75), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT17), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n435), .B1(new_n434), .B2(KEYINPUT76), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n435), .B(KEYINPUT17), .C1(new_n434), .C2(KEYINPUT76), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n426), .A2(new_n430), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n342), .A2(new_n343), .A3(new_n378), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n340), .A2(new_n341), .ZN(new_n442));
  INV_X1    g0242(.A(new_n331), .ZN(new_n443));
  INV_X1    g0243(.A(new_n298), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n378), .A2(new_n440), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT77), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G303), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n383), .A2(G33), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n380), .A2(KEYINPUT3), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n354), .A2(G257), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G264), .A2(G1698), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n381), .A2(new_n384), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n452), .A2(new_n455), .A3(new_n281), .ZN(new_n456));
  XNOR2_X1  g0256(.A(KEYINPUT5), .B(G41), .ZN(new_n457));
  INV_X1    g0257(.A(G45), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(G1), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(G274), .A3(new_n459), .ZN(new_n460));
  AND2_X1   g0260(.A1(KEYINPUT5), .A2(G41), .ZN(new_n461));
  NOR2_X1   g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(G270), .A3(new_n280), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n456), .A2(new_n460), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT82), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n456), .A2(KEYINPUT82), .A3(new_n460), .A4(new_n464), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n467), .A2(G169), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT83), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(KEYINPUT20), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(KEYINPUT20), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n232), .ZN(new_n476));
  AND2_X1   g0276(.A1(KEYINPUT79), .A2(G97), .ZN(new_n477));
  NOR2_X1   g0277(.A1(KEYINPUT79), .A2(G97), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n476), .B1(new_n479), .B2(new_n380), .ZN(new_n480));
  INV_X1    g0280(.A(G116), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n260), .A2(new_n231), .B1(G20), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n474), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT79), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n217), .ZN(new_n486));
  NAND2_X1  g0286(.A1(KEYINPUT79), .A2(G97), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n486), .A2(new_n380), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n476), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(new_n473), .A3(new_n482), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n472), .B1(new_n484), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT84), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n305), .A2(G116), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n262), .B(new_n268), .C1(G1), .C2(new_n380), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(G116), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n492), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n472), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n490), .A2(new_n473), .A3(new_n482), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n473), .B1(new_n490), .B2(new_n482), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n496), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT84), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n470), .B1(new_n497), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT86), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT21), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n493), .B1(new_n492), .B2(new_n496), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n501), .A2(KEYINPUT84), .A3(new_n502), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n469), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT86), .B1(new_n510), .B2(KEYINPUT21), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n508), .A2(new_n509), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n467), .A2(KEYINPUT21), .A3(G169), .A4(new_n468), .ZN(new_n514));
  OR2_X1    g0314(.A1(new_n465), .A2(new_n337), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n513), .A2(new_n516), .A3(KEYINPUT85), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT85), .B1(new_n513), .B2(new_n516), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n513), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n467), .A2(new_n468), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G200), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n520), .B(new_n522), .C1(new_n289), .C2(new_n521), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n512), .A2(new_n519), .A3(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n268), .A2(G97), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n495), .A2(new_n217), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G107), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(new_n400), .B2(new_n402), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n479), .A2(KEYINPUT6), .A3(new_n529), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT6), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n217), .A2(new_n529), .ZN(new_n533));
  NOR2_X1   g0333(.A1(G97), .A2(G107), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n232), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n254), .A2(G77), .ZN(new_n537));
  XNOR2_X1  g0337(.A(new_n537), .B(KEYINPUT78), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n530), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n526), .B(new_n528), .C1(new_n539), .C2(new_n262), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT80), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n381), .A2(new_n384), .A3(G244), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT4), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n544), .A2(G1698), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n276), .A2(G244), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n547), .A3(new_n475), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n276), .A2(G250), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n354), .B1(new_n549), .B2(KEYINPUT4), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n542), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(KEYINPUT4), .B1(new_n409), .B2(new_n216), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G1698), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n543), .A2(new_n544), .B1(G33), .B2(G283), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n553), .A2(KEYINPUT80), .A3(new_n554), .A4(new_n547), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n551), .A2(new_n555), .A3(new_n281), .ZN(new_n556));
  INV_X1    g0356(.A(new_n460), .ZN(new_n557));
  INV_X1    g0357(.A(new_n231), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n457), .A2(new_n459), .B1(new_n558), .B2(new_n279), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n557), .B1(G257), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G200), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n556), .A2(G190), .A3(new_n560), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n541), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(new_n294), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n556), .A2(new_n337), .A3(new_n560), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n540), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n559), .A2(G264), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n216), .A2(new_n354), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n218), .A2(G1698), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n381), .A2(new_n570), .A3(new_n384), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G33), .A2(G294), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n281), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT89), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n569), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n280), .B1(new_n572), .B2(new_n573), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n460), .B1(new_n578), .B2(KEYINPUT89), .ZN(new_n579));
  OR2_X1    g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n281), .A2(new_n574), .B1(new_n559), .B2(G264), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n581), .A2(new_n460), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n580), .A2(G190), .B1(G200), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n305), .A2(KEYINPUT25), .A3(new_n529), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(KEYINPUT25), .B1(new_n305), .B2(new_n529), .ZN(new_n586));
  OAI22_X1  g0386(.A1(new_n495), .A2(new_n529), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT88), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n381), .A2(new_n384), .A3(new_n232), .A4(G87), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT22), .ZN(new_n591));
  OR2_X1    g0391(.A1(new_n591), .A2(KEYINPUT87), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n276), .A2(new_n232), .A3(new_n592), .A4(G87), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n232), .A2(G107), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n597), .B(KEYINPUT23), .ZN(new_n598));
  NAND2_X1  g0398(.A1(G33), .A2(G116), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(G20), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n596), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT24), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n600), .B1(new_n594), .B2(new_n595), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT24), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(new_n605), .A3(new_n598), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n589), .B1(new_n607), .B2(new_n261), .ZN(new_n608));
  AOI211_X1 g0408(.A(KEYINPUT88), .B(new_n262), .C1(new_n603), .C2(new_n606), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n583), .B(new_n588), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n215), .B(new_n529), .C1(new_n477), .C2(new_n478), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT19), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n232), .B1(new_n314), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n486), .A2(new_n487), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n612), .B1(new_n615), .B2(new_n256), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n276), .A2(new_n232), .A3(G68), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n618), .A2(new_n261), .B1(new_n305), .B2(new_n258), .ZN(new_n619));
  INV_X1    g0419(.A(new_n495), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n257), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n224), .A2(G1698), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n276), .B(new_n623), .C1(G238), .C2(G1698), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n280), .B1(new_n624), .B2(new_n599), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n459), .A2(new_n284), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n216), .B1(new_n458), .B2(G1), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(new_n280), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n337), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n294), .B1(new_n625), .B2(new_n629), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n622), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(G200), .B1(new_n625), .B2(new_n629), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n620), .A2(G87), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(new_n619), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT81), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n636), .A2(new_n637), .B1(G190), .B2(new_n630), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n634), .A2(new_n619), .A3(KEYINPUT81), .A4(new_n635), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n633), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n606), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n605), .B1(new_n604), .B2(new_n598), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n261), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT88), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n607), .A2(new_n589), .A3(new_n261), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n587), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n580), .A2(G169), .B1(G179), .B2(new_n582), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n610), .B(new_n640), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n524), .A2(new_n568), .A3(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n448), .A2(new_n649), .ZN(G372));
  OAI21_X1  g0450(.A(new_n588), .B1(new_n608), .B2(new_n609), .ZN(new_n651));
  INV_X1    g0451(.A(new_n647), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n513), .A2(new_n516), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n512), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n622), .A2(new_n631), .A3(new_n632), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n630), .A2(G190), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n657), .A2(new_n619), .A3(new_n634), .A4(new_n635), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n564), .A2(new_n660), .A3(new_n567), .ZN(new_n661));
  AOI21_X1  g0461(.A(G200), .B1(new_n581), .B2(new_n460), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n577), .A2(new_n579), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n662), .B1(new_n663), .B2(new_n289), .ZN(new_n664));
  AOI211_X1 g0464(.A(new_n587), .B(new_n664), .C1(new_n644), .C2(new_n645), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n655), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n567), .ZN(new_n668));
  XOR2_X1   g0468(.A(KEYINPUT90), .B(KEYINPUT26), .Z(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(new_n640), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n567), .A2(new_n659), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(KEYINPUT26), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n667), .A2(new_n656), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n448), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n438), .A2(new_n439), .ZN(new_n675));
  INV_X1    g0475(.A(new_n442), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT91), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n297), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n293), .A2(KEYINPUT91), .A3(new_n295), .A4(new_n296), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n331), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n675), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n419), .B(KEYINPUT18), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n373), .A2(new_n377), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n363), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n674), .A2(new_n685), .ZN(G369));
  NAND2_X1  g0486(.A1(new_n512), .A2(new_n654), .ZN(new_n687));
  INV_X1    g0487(.A(G13), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G20), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n263), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G213), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G343), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n520), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n687), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n524), .B2(new_n697), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G330), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n653), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(new_n665), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n646), .B2(new_n696), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n653), .B2(new_n696), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n695), .B1(new_n512), .B2(new_n519), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n703), .A2(new_n707), .B1(new_n702), .B2(new_n696), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(G399));
  INV_X1    g0509(.A(new_n211), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G41), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G1), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n611), .A2(G116), .ZN(new_n714));
  OAI22_X1  g0514(.A1(new_n713), .A2(new_n714), .B1(new_n234), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT29), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n512), .A2(new_n519), .A3(new_n653), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT92), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n512), .A2(new_n519), .A3(new_n653), .A4(KEYINPUT92), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(new_n666), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n671), .A2(KEYINPUT26), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n668), .A2(new_n640), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(new_n669), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n722), .A2(new_n656), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n717), .B1(new_n726), .B2(new_n696), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n673), .A2(new_n696), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(KEYINPUT29), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n515), .A2(new_n625), .A3(new_n629), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(new_n560), .A3(new_n556), .A4(new_n581), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT30), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n582), .A2(new_n630), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n561), .A2(new_n734), .A3(new_n337), .A4(new_n521), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT31), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n736), .A2(new_n737), .A3(new_n695), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n737), .B1(new_n649), .B2(new_n696), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n736), .A2(new_n695), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G330), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n730), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n716), .B1(new_n744), .B2(G1), .ZN(G364));
  NOR2_X1   g0545(.A1(G13), .A2(G33), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n699), .A2(new_n749), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n289), .A2(G179), .A3(G200), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n232), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n232), .A2(G179), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n754), .A2(new_n289), .A3(new_n329), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n753), .A2(G294), .B1(new_n756), .B2(G329), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n289), .A2(new_n329), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(new_n754), .ZN(new_n759));
  INV_X1    g0559(.A(G322), .ZN(new_n760));
  NAND2_X1  g0560(.A1(G20), .A2(G179), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n761), .A2(new_n289), .A3(G200), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n757), .B1(new_n449), .B2(new_n759), .C1(new_n760), .C2(new_n763), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n761), .A2(new_n329), .A3(G190), .ZN(new_n765));
  XNOR2_X1  g0565(.A(KEYINPUT33), .B(G317), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n761), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n758), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G326), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n754), .A2(new_n289), .A3(G200), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n772), .A2(KEYINPUT94), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(KEYINPUT94), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G283), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n761), .A2(G190), .A3(G200), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n276), .B1(G311), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n767), .A2(new_n771), .A3(new_n776), .A4(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n775), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n276), .B1(new_n780), .B2(new_n529), .ZN(new_n781));
  INV_X1    g0581(.A(new_n759), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n781), .B1(G87), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n765), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n752), .A2(new_n217), .B1(new_n784), .B2(new_n306), .ZN(new_n785));
  INV_X1    g0585(.A(G159), .ZN(new_n786));
  OAI21_X1  g0586(.A(KEYINPUT32), .B1(new_n755), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(new_n202), .B2(new_n769), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n785), .B(new_n788), .C1(G77), .C2(new_n777), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n756), .A2(G159), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n783), .B(new_n789), .C1(KEYINPUT32), .C2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n763), .A2(new_n226), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n779), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n231), .B1(G20), .B2(new_n294), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n276), .A2(G355), .A3(new_n211), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n248), .A2(G45), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT93), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n710), .A2(new_n276), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(G45), .B2(new_n234), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n796), .B1(G116), .B2(new_n211), .C1(new_n798), .C2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n748), .A2(new_n794), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n713), .B1(G45), .B2(new_n689), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n750), .A2(new_n795), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n699), .A2(G330), .ZN(new_n806));
  INV_X1    g0606(.A(new_n804), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n700), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n805), .B1(new_n806), .B2(new_n808), .ZN(G396));
  OAI21_X1  g0609(.A(new_n298), .B1(new_n275), .B2(new_n696), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n678), .A2(new_n293), .A3(new_n679), .A4(new_n695), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n728), .B(new_n812), .Z(new_n813));
  OR2_X1    g0613(.A1(new_n813), .A2(new_n743), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n743), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n814), .A2(new_n807), .A3(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n812), .A2(new_n747), .ZN(new_n817));
  INV_X1    g0617(.A(new_n794), .ZN(new_n818));
  INV_X1    g0618(.A(new_n777), .ZN(new_n819));
  INV_X1    g0619(.A(G283), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n819), .A2(new_n481), .B1(new_n784), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT96), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n823), .B(new_n824), .C1(new_n449), .C2(new_n769), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT97), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n409), .B1(new_n752), .B2(new_n217), .ZN(new_n827));
  INV_X1    g0627(.A(G311), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n755), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n780), .A2(new_n215), .ZN(new_n830));
  NOR4_X1   g0630(.A1(new_n826), .A2(new_n827), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G294), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n831), .B1(new_n529), .B2(new_n759), .C1(new_n832), .C2(new_n763), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n756), .A2(G132), .ZN(new_n834));
  XNOR2_X1  g0634(.A(KEYINPUT98), .B(G143), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n762), .A2(new_n835), .B1(new_n777), .B2(G159), .ZN(new_n836));
  INV_X1    g0636(.A(G137), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n836), .B1(new_n837), .B2(new_n769), .C1(new_n348), .C2(new_n784), .ZN(new_n838));
  XNOR2_X1  g0638(.A(KEYINPUT99), .B(KEYINPUT34), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n834), .B1(new_n202), .B2(new_n759), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(G58), .B2(new_n753), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n409), .B1(new_n838), .B2(new_n839), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n841), .B(new_n842), .C1(new_n306), .C2(new_n780), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n818), .B1(new_n833), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n817), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n794), .A2(new_n746), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT95), .Z(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n206), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n845), .A2(new_n804), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n816), .A2(new_n849), .ZN(G384));
  NAND2_X1  g0650(.A1(new_n531), .A2(new_n535), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n481), .B1(new_n851), .B2(KEYINPUT35), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n852), .B(new_n233), .C1(KEYINPUT35), .C2(new_n851), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT36), .ZN(new_n854));
  OAI21_X1  g0654(.A(G77), .B1(new_n226), .B2(new_n306), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n855), .A2(new_n234), .B1(G50), .B2(new_n306), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n856), .A2(G1), .A3(new_n688), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT100), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n434), .B1(new_n424), .B2(new_n395), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n424), .A2(new_n693), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT37), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n419), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n415), .A2(new_n418), .ZN(new_n864));
  INV_X1    g0664(.A(new_n693), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT37), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n863), .A2(new_n866), .A3(new_n867), .A4(new_n434), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n862), .A2(KEYINPUT101), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT101), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n870), .B(KEYINPUT37), .C1(new_n860), .C2(new_n861), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT76), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n424), .A2(new_n873), .A3(new_n432), .A4(new_n433), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n424), .A2(KEYINPUT75), .A3(new_n432), .A4(new_n433), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n435), .A2(new_n874), .B1(new_n875), .B2(KEYINPUT17), .ZN(new_n876));
  INV_X1    g0676(.A(new_n439), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n682), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n861), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT38), .B1(new_n872), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n423), .B1(KEYINPUT16), .B2(new_n422), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n881), .A2(new_n418), .ZN(new_n882));
  OR2_X1    g0682(.A1(new_n882), .A2(new_n693), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n419), .A2(KEYINPUT18), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT73), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n419), .A2(new_n427), .A3(KEYINPUT18), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n885), .A2(new_n420), .A3(new_n886), .A4(new_n425), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n883), .B1(new_n675), .B2(new_n887), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n392), .A2(new_n394), .A3(new_n865), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n434), .B1(new_n882), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n868), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n888), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT102), .B1(new_n880), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n866), .B1(new_n675), .B2(new_n682), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n869), .A2(new_n871), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT102), .ZN(new_n900));
  OAI211_X1 g0700(.A(KEYINPUT38), .B(new_n892), .C1(new_n440), .C2(new_n883), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n896), .A2(new_n902), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n512), .A2(new_n519), .A3(new_n523), .ZN(new_n904));
  INV_X1    g0704(.A(new_n568), .ZN(new_n905));
  INV_X1    g0705(.A(new_n648), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n904), .A2(new_n905), .A3(new_n906), .A4(new_n696), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(KEYINPUT31), .A3(new_n741), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n341), .A2(new_n695), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n333), .A2(new_n335), .A3(new_n338), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n443), .B(new_n909), .C1(new_n910), .C2(new_n310), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n340), .A2(new_n341), .A3(new_n695), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n908), .A2(new_n738), .A3(new_n812), .A4(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT40), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n894), .B1(new_n888), .B2(new_n893), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n901), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n742), .A2(new_n812), .A3(new_n918), .A4(new_n913), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n903), .A2(new_n916), .B1(new_n919), .B2(new_n915), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n920), .A2(new_n448), .A3(new_n742), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n917), .A2(new_n901), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n915), .B1(new_n914), .B2(new_n922), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n742), .A2(KEYINPUT40), .A3(new_n812), .A4(new_n913), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n896), .A2(new_n902), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n923), .B(G330), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n448), .A2(new_n742), .A3(G330), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n921), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n673), .A2(new_n696), .A3(new_n812), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n297), .A2(new_n695), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(new_n918), .A3(new_n913), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n682), .A2(new_n865), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  AND3_X1   g0736(.A1(new_n917), .A2(new_n901), .A3(KEYINPUT39), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT39), .B1(new_n899), .B2(new_n901), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n442), .A2(new_n695), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n937), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n936), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n929), .B(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n448), .B1(new_n727), .B2(new_n729), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n685), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n943), .B(new_n945), .Z(new_n946));
  NOR2_X1   g0746(.A1(new_n689), .A2(new_n263), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n859), .B1(new_n946), .B2(new_n947), .ZN(G367));
  OAI21_X1  g0748(.A(new_n905), .B1(new_n541), .B2(new_n696), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n668), .A2(new_n695), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n706), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n696), .B1(new_n619), .B2(new_n635), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT103), .Z(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n633), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n659), .B2(new_n955), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT104), .Z(new_n959));
  XNOR2_X1  g0759(.A(new_n953), .B(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n703), .A2(new_n707), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(new_n949), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT42), .Z(new_n964));
  OAI21_X1  g0764(.A(new_n567), .B1(new_n949), .B2(new_n653), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n965), .A2(new_n696), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n961), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n960), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n960), .A2(new_n967), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n689), .A2(G45), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(G1), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT107), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n708), .A2(new_n951), .ZN(new_n976));
  XOR2_X1   g0776(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n977));
  XNOR2_X1  g0777(.A(new_n976), .B(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n708), .A2(new_n951), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT45), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n706), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n962), .B1(new_n705), .B2(new_n707), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n982), .B1(new_n700), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n744), .A2(new_n981), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n744), .ZN(new_n986));
  XNOR2_X1  g0786(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n711), .B(new_n987), .Z(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n975), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n957), .A2(new_n749), .ZN(new_n991));
  INV_X1    g0791(.A(new_n799), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n802), .B1(new_n211), .B2(new_n258), .C1(new_n244), .C2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT108), .Z(new_n994));
  OAI22_X1  g0794(.A1(new_n819), .A2(new_n202), .B1(new_n763), .B2(new_n348), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n409), .B(new_n995), .C1(G68), .C2(new_n753), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n775), .A2(G77), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n770), .A2(new_n835), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n755), .A2(new_n837), .B1(new_n759), .B2(new_n226), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(G159), .B2(new_n765), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n996), .A2(new_n997), .A3(new_n998), .A4(new_n1000), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n763), .A2(new_n449), .B1(new_n769), .B2(new_n828), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT109), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n409), .B1(new_n752), .B2(new_n529), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT110), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n759), .B2(new_n481), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1004), .B1(KEYINPUT46), .B2(new_n1006), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1007), .B1(KEYINPUT46), .B2(new_n1006), .C1(new_n780), .C2(new_n615), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1003), .B(new_n1008), .C1(G317), .C2(new_n756), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n820), .B2(new_n819), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n784), .A2(new_n832), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1001), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT111), .Z(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT47), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n804), .B(new_n994), .C1(new_n1014), .C2(new_n818), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT112), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n971), .A2(new_n990), .B1(new_n991), .B2(new_n1017), .ZN(G387));
  NAND2_X1  g0818(.A1(new_n984), .A2(new_n975), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n819), .A2(new_n306), .B1(new_n769), .B2(new_n786), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n409), .B1(new_n782), .B2(G77), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n348), .B2(new_n755), .C1(new_n780), .C2(new_n217), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT113), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1020), .B(new_n1023), .C1(G50), .C2(new_n762), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n258), .B2(new_n752), .C1(new_n347), .C2(new_n784), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G303), .A2(new_n777), .B1(new_n765), .B2(G311), .ZN(new_n1026));
  INV_X1    g0826(.A(G317), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1026), .B1(new_n1027), .B2(new_n763), .C1(new_n760), .C2(new_n769), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT48), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n820), .B2(new_n752), .C1(new_n832), .C2(new_n759), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT49), .Z(new_n1031));
  AOI21_X1  g0831(.A(new_n276), .B1(new_n756), .B2(G326), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n780), .B2(new_n481), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1025), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n794), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n253), .A2(new_n202), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT50), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n306), .A2(new_n206), .ZN(new_n1038));
  NOR4_X1   g0838(.A1(new_n1037), .A2(G45), .A3(new_n1038), .A4(new_n714), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n799), .B1(new_n240), .B2(new_n458), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n714), .A2(new_n211), .A3(new_n276), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n211), .A2(G107), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n802), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n705), .A2(new_n749), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1035), .A2(new_n804), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n744), .A2(new_n984), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n711), .B1(new_n744), .B2(new_n984), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1019), .B(new_n1046), .C1(new_n1048), .C2(new_n1049), .ZN(G393));
  XNOR2_X1  g0850(.A(new_n981), .B(new_n982), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1051), .A2(new_n974), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n802), .B1(new_n211), .B2(new_n615), .C1(new_n251), .C2(new_n992), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n807), .B1(new_n952), .B2(new_n748), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n770), .A2(G150), .B1(G159), .B2(new_n762), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT51), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n752), .A2(new_n206), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n202), .A2(new_n784), .B1(new_n819), .B2(new_n347), .ZN(new_n1058));
  NOR4_X1   g0858(.A1(new_n830), .A2(new_n1056), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n756), .A2(new_n835), .B1(new_n782), .B2(G68), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT114), .Z(new_n1061));
  AND3_X1   g0861(.A1(new_n1059), .A2(new_n276), .A3(new_n1061), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n763), .A2(new_n828), .B1(new_n769), .B2(new_n1027), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT52), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n820), .B2(new_n759), .C1(new_n529), .C2(new_n780), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n752), .A2(new_n481), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n819), .A2(new_n832), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n409), .B1(new_n755), .B2(new_n760), .C1(new_n784), .C2(new_n449), .ZN(new_n1068));
  NOR4_X1   g0868(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n794), .B1(new_n1062), .B2(new_n1069), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n1054), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1052), .B1(new_n1053), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1051), .A2(new_n1047), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1073), .A2(new_n711), .A3(new_n985), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1074), .ZN(G390));
  AND2_X1   g0875(.A1(new_n911), .A2(new_n912), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n930), .B2(new_n931), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1077), .A2(new_n939), .B1(new_n937), .B2(new_n938), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n726), .A2(new_n696), .A3(new_n812), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1076), .B1(new_n1079), .B2(new_n931), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n896), .A2(new_n902), .A3(new_n940), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(G330), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n914), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT115), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1082), .B(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n975), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n746), .B1(new_n937), .B2(new_n938), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n847), .A2(new_n347), .ZN(new_n1090));
  XOR2_X1   g0890(.A(KEYINPUT54), .B(G143), .Z(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1092), .A2(new_n819), .ZN(new_n1093));
  INV_X1    g0893(.A(G132), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n276), .B1(new_n763), .B2(new_n1094), .C1(new_n837), .C2(new_n784), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1093), .B(new_n1095), .C1(G159), .C2(new_n753), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n775), .A2(G50), .B1(G125), .B2(new_n756), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n770), .A2(G128), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n759), .A2(new_n348), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT53), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n770), .A2(G283), .B1(new_n479), .B2(new_n777), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n529), .B2(new_n784), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1103), .A2(KEYINPUT116), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1057), .B1(new_n1103), .B2(KEYINPUT116), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n756), .A2(G294), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n775), .A2(G68), .B1(G116), .B2(new_n762), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n409), .B1(new_n759), .B2(new_n215), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT117), .Z(new_n1110));
  OAI21_X1  g0910(.A(new_n1101), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n794), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1089), .A2(new_n804), .A3(new_n1090), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1088), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n908), .A2(G330), .A3(new_n738), .A4(new_n812), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n1076), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n932), .B1(new_n1117), .B2(new_n1084), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n742), .A2(G330), .A3(new_n812), .A4(new_n913), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1119), .A2(new_n931), .A3(new_n1079), .A4(new_n1116), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n944), .A2(new_n685), .A3(new_n927), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  OR2_X1    g0925(.A1(new_n1125), .A2(new_n1087), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n712), .B1(new_n1125), .B2(new_n1087), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1114), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(G378));
  AOI22_X1  g0929(.A1(new_n753), .A2(G150), .B1(new_n770), .B2(G125), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1130), .B(KEYINPUT120), .Z(new_n1131));
  NOR2_X1   g0931(.A1(new_n1092), .A2(new_n759), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1133), .A2(KEYINPUT119), .B1(G128), .B2(new_n762), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1135), .B1(new_n1094), .B2(new_n784), .C1(new_n837), .C2(new_n819), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT119), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1136), .B1(new_n1137), .B2(new_n1132), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(G41), .B1(new_n1139), .B2(KEYINPUT59), .ZN(new_n1140));
  AOI21_X1  g0940(.A(G33), .B1(new_n756), .B2(G124), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1140), .B(new_n1141), .C1(new_n786), .C2(new_n780), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1139), .A2(KEYINPUT59), .ZN(new_n1143));
  AOI21_X1  g0943(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n1142), .A2(new_n1143), .B1(G50), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  AOI211_X1 g0946(.A(G41), .B(new_n276), .C1(new_n782), .C2(G77), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT118), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n775), .A2(G58), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n753), .A2(G68), .B1(new_n770), .B2(G116), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(new_n258), .C2(new_n819), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1148), .B(new_n1151), .C1(G97), .C2(new_n765), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1152), .B1(new_n529), .B2(new_n763), .C1(new_n820), .C2(new_n755), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT58), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n818), .B1(new_n1146), .B2(new_n1154), .ZN(new_n1155));
  XOR2_X1   g0955(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n378), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n378), .A2(new_n1157), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n353), .A2(new_n693), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1158), .A2(new_n1161), .A3(new_n1159), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1166), .A2(new_n747), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n846), .A2(new_n202), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NOR4_X1   g0969(.A1(new_n1155), .A2(new_n1167), .A3(new_n807), .A4(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1166), .B1(new_n936), .B2(new_n941), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n934), .B1(new_n1077), .B2(new_n918), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT39), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n880), .B2(new_n895), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n917), .A2(new_n901), .A3(KEYINPUT39), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1174), .A2(new_n939), .A3(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1172), .A2(new_n1176), .A3(new_n1165), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1171), .A2(new_n920), .A3(G330), .A4(new_n1177), .ZN(new_n1178));
  AND4_X1   g0978(.A1(new_n1176), .A2(new_n933), .A3(new_n935), .A4(new_n1165), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1165), .B1(new_n1172), .B2(new_n1176), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n926), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n1178), .A2(new_n1181), .A3(KEYINPUT121), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT121), .B1(new_n1178), .B2(new_n1181), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1170), .B1(new_n1184), .B2(new_n975), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1082), .A2(new_n1085), .A3(new_n1084), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1086), .B(new_n1078), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1186), .A2(new_n1121), .A3(new_n1187), .A4(new_n1123), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n1123), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT57), .B1(new_n1184), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1178), .A2(new_n1181), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1189), .A2(new_n1192), .A3(KEYINPUT57), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n711), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1185), .B1(new_n1190), .B2(new_n1194), .ZN(G375));
  NAND3_X1  g0995(.A1(new_n1118), .A2(new_n1122), .A3(new_n1120), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1124), .A2(new_n989), .A3(new_n1196), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1149), .B1(new_n1094), .B2(new_n769), .C1(new_n348), .C2(new_n819), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n765), .B2(new_n1091), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n782), .A2(G159), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n753), .A2(G50), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n409), .B1(G137), .B2(new_n762), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G128), .B2(new_n756), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n775), .A2(G77), .B1(G294), .B2(new_n770), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n755), .A2(new_n449), .B1(new_n759), .B2(new_n217), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT122), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1206), .A2(new_n1207), .B1(new_n257), .B2(new_n753), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1205), .B(new_n1208), .C1(new_n1207), .C2(new_n1206), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n819), .A2(new_n529), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n763), .A2(new_n820), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n409), .B1(new_n784), .B2(new_n481), .ZN(new_n1212));
  NOR4_X1   g1012(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n794), .B1(new_n1204), .B2(new_n1213), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n804), .B(new_n1214), .C1(new_n913), .C2(new_n747), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n306), .B2(new_n847), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n1121), .B2(new_n975), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1197), .A2(new_n1217), .ZN(G381));
  INV_X1    g1018(.A(G390), .ZN(new_n1219));
  INV_X1    g1019(.A(G387), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(G393), .A2(G396), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1222), .A2(G384), .A3(G381), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT121), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1177), .A2(new_n1171), .B1(new_n920), .B2(G330), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1179), .A2(new_n1180), .A3(new_n926), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1224), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1178), .A2(new_n1181), .A3(KEYINPUT121), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1227), .A2(new_n975), .A3(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1170), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1227), .A2(new_n1189), .A3(new_n1228), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT57), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1191), .B1(new_n1123), .B2(new_n1188), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n712), .B1(new_n1235), .B2(KEYINPUT57), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1231), .B1(new_n1234), .B2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1223), .A2(new_n1128), .A3(new_n1237), .ZN(G407));
  NOR2_X1   g1038(.A1(new_n1223), .A2(new_n694), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1237), .A2(new_n1128), .ZN(new_n1240));
  OAI21_X1  g1040(.A(G213), .B1(new_n1239), .B2(new_n1240), .ZN(G409));
  INV_X1    g1041(.A(KEYINPUT127), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT61), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT63), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n816), .A2(KEYINPUT124), .A3(new_n849), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1079), .A2(new_n931), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1117), .A2(new_n1084), .A3(new_n1246), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1119), .A2(new_n1116), .B1(new_n930), .B2(new_n931), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT123), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1249), .A2(new_n1250), .A3(KEYINPUT60), .A4(new_n1122), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT60), .ZN(new_n1252));
  OAI21_X1  g1052(.A(KEYINPUT123), .B1(new_n1196), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n712), .B1(new_n1196), .B2(new_n1252), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1124), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1217), .B(new_n1245), .C1(new_n1254), .C2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(KEYINPUT124), .B1(new_n816), .B2(new_n849), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1251), .A2(new_n1253), .A3(new_n1255), .A4(new_n1124), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1258), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1260), .A2(new_n1217), .A3(new_n1261), .A4(new_n1245), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n694), .A2(G213), .A3(G2897), .ZN(new_n1263));
  XOR2_X1   g1063(.A(new_n1263), .B(KEYINPUT125), .Z(new_n1264));
  AND3_X1   g1064(.A1(new_n1259), .A2(new_n1262), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1264), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n694), .A2(G213), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1184), .A2(new_n989), .A3(new_n1189), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1192), .A2(new_n975), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1128), .A2(new_n1269), .A3(new_n1230), .A4(new_n1270), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1268), .B(new_n1271), .C1(new_n1237), .C2(new_n1128), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1244), .B1(new_n1267), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1259), .A2(new_n1262), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1243), .B1(new_n1273), .B2(new_n1276), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(G393), .B(G396), .ZN(new_n1278));
  OR2_X1    g1078(.A1(new_n1278), .A2(G387), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(G387), .A3(KEYINPUT126), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1219), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1279), .A2(new_n1280), .A3(G390), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(G375), .A2(G378), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1285), .A2(new_n1268), .A3(new_n1271), .A4(new_n1274), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1284), .B1(new_n1244), .B2(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1277), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT62), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT61), .B1(new_n1276), .B2(new_n1289), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n1286), .A2(KEYINPUT62), .B1(new_n1272), .B2(new_n1267), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1284), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1242), .B1(new_n1288), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1294), .B1(new_n1276), .B2(KEYINPUT63), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1295), .B(new_n1243), .C1(new_n1276), .C2(new_n1273), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1267), .A2(new_n1272), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1297), .B1(new_n1276), .B2(new_n1289), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1243), .B1(new_n1286), .B2(KEYINPUT62), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1294), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1296), .A2(new_n1300), .A3(KEYINPUT127), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1293), .A2(new_n1301), .ZN(G405));
  NAND2_X1  g1102(.A1(new_n1285), .A2(new_n1240), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(new_n1303), .B(new_n1274), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(new_n1304), .B(new_n1284), .ZN(G402));
endmodule


