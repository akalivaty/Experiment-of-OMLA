//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n789, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003;
  AND2_X1   g000(.A1(KEYINPUT69), .A2(G134gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(KEYINPUT69), .A2(G134gat), .ZN(new_n203));
  OAI21_X1  g002(.A(G127gat), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G127gat), .B2(G134gat), .ZN(new_n205));
  INV_X1    g004(.A(G113gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(G120gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(G120gat), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT1), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT70), .B1(new_n205), .B2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(G127gat), .A2(G134gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT69), .B(G134gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n212), .B1(new_n213), .B2(G127gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT70), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n216));
  INV_X1    g015(.A(new_n209), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n216), .B1(new_n217), .B2(new_n207), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n214), .A2(new_n215), .A3(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n207), .B1(new_n217), .B2(KEYINPUT71), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(KEYINPUT71), .B2(new_n217), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT72), .B(KEYINPUT1), .ZN(new_n222));
  AND2_X1   g021(.A1(G127gat), .A2(G134gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n212), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n211), .A2(new_n219), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G183gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT27), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT27), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G183gat), .ZN(new_n230));
  INV_X1    g029(.A(G190gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n228), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n232), .A2(KEYINPUT28), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(KEYINPUT28), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n227), .A2(new_n231), .ZN(new_n235));
  NOR3_X1   g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT65), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT26), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(G169gat), .B2(G176gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n238), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT68), .ZN(new_n243));
  NAND2_X1  g042(.A1(G169gat), .A2(G176gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n238), .A2(new_n245), .A3(new_n241), .A4(new_n239), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n243), .A2(new_n244), .A3(new_n246), .A4(new_n249), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n236), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT25), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT64), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n227), .A2(new_n231), .ZN(new_n254));
  NAND3_X1  g053(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n253), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n257), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n259), .A2(new_n254), .A3(KEYINPUT64), .A4(new_n255), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n237), .A2(KEYINPUT23), .ZN(new_n261));
  INV_X1    g060(.A(new_n237), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n244), .A2(KEYINPUT23), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n258), .A2(new_n260), .A3(new_n261), .A4(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n257), .B(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n267), .A2(new_n254), .A3(new_n255), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n238), .A2(KEYINPUT23), .A3(new_n241), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n269), .A2(new_n264), .A3(KEYINPUT25), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n252), .A2(new_n265), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n226), .B1(new_n251), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G227gat), .A2(G233gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n265), .A2(new_n252), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n268), .A2(new_n270), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n221), .A2(new_n225), .ZN(new_n278));
  INV_X1    g077(.A(new_n219), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n215), .B1(new_n214), .B2(new_n218), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n236), .A2(new_n250), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n277), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n272), .A2(new_n274), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT33), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT73), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n284), .A2(new_n288), .A3(new_n285), .ZN(new_n289));
  XNOR2_X1  g088(.A(G15gat), .B(G43gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT74), .ZN(new_n291));
  XOR2_X1   g090(.A(G71gat), .B(G99gat), .Z(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n293), .B1(new_n284), .B2(KEYINPUT32), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n287), .A2(new_n289), .A3(new_n294), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n284), .B(KEYINPUT32), .C1(new_n285), .C2(new_n293), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n274), .B1(new_n272), .B2(new_n283), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT34), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT75), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n299), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n295), .A2(new_n296), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT77), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n295), .A2(new_n296), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n297), .A2(new_n301), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(new_n306), .A3(new_n299), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT77), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n295), .A2(new_n308), .A3(new_n296), .A4(new_n302), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n304), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G228gat), .ZN(new_n311));
  INV_X1    g110(.A(G233gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(G211gat), .B(G218gat), .Z(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G197gat), .B(G204gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT22), .ZN(new_n318));
  INV_X1    g117(.A(G211gat), .ZN(new_n319));
  INV_X1    g118(.A(G218gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n316), .A2(new_n317), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT86), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n317), .A2(new_n321), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n315), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n322), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n324), .A2(new_n315), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT29), .B1(new_n327), .B2(KEYINPUT86), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT3), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT80), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT80), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n332), .A2(G155gat), .A3(G162gat), .ZN(new_n333));
  INV_X1    g132(.A(G155gat), .ZN(new_n334));
  INV_X1    g133(.A(G162gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n331), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G141gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(G148gat), .ZN(new_n340));
  INV_X1    g139(.A(G148gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G141gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n332), .A2(KEYINPUT2), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n330), .B1(new_n336), .B2(KEYINPUT2), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT81), .B1(new_n341), .B2(G141gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT81), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(new_n339), .A3(G148gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n349), .A3(new_n342), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n338), .A2(new_n345), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n329), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n322), .A2(new_n325), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n353), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n314), .B1(new_n352), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n322), .A2(new_n325), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n354), .B1(new_n359), .B2(KEYINPUT29), .ZN(new_n360));
  INV_X1    g159(.A(new_n351), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n314), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n357), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT87), .B1(new_n358), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(G78gat), .B(G106gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT31), .B(G50gat), .ZN(new_n367));
  XOR2_X1   g166(.A(new_n366), .B(new_n367), .Z(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(G22gat), .B1(new_n365), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(G22gat), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n363), .B1(new_n351), .B2(new_n329), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n372), .A2(new_n314), .B1(new_n362), .B2(new_n363), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n371), .B(new_n368), .C1(new_n373), .C2(KEYINPUT87), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(KEYINPUT87), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n370), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n376), .B1(new_n370), .B2(new_n374), .ZN(new_n379));
  NOR3_X1   g178(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT35), .ZN(new_n380));
  XNOR2_X1  g179(.A(G1gat), .B(G29gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT0), .ZN(new_n382));
  XNOR2_X1  g181(.A(G57gat), .B(G85gat), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n382), .B(new_n383), .Z(new_n384));
  NAND2_X1  g183(.A1(new_n281), .A2(new_n361), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n351), .B(new_n278), .C1(new_n279), .C2(new_n280), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G225gat), .A2(G233gat), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n388), .B(KEYINPUT82), .Z(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n350), .A2(new_n346), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n337), .B1(new_n343), .B2(new_n344), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT3), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n281), .A2(new_n355), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT83), .B(KEYINPUT4), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n386), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n226), .A2(KEYINPUT4), .A3(new_n351), .ZN(new_n398));
  INV_X1    g197(.A(new_n389), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n395), .A2(new_n397), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT84), .B(KEYINPUT5), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n390), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n394), .A2(new_n355), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n399), .B(new_n401), .C1(new_n404), .C2(new_n226), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT85), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n386), .A2(new_n407), .A3(KEYINPUT4), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n226), .A2(new_n351), .A3(new_n396), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n407), .B1(new_n386), .B2(KEYINPUT4), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n406), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n384), .B1(new_n403), .B2(new_n412), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n413), .A2(KEYINPUT6), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n403), .A2(new_n412), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT88), .ZN(new_n416));
  INV_X1    g215(.A(new_n384), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT88), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n403), .A2(new_n412), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n416), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT6), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n421), .B1(new_n415), .B2(new_n417), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n414), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G8gat), .B(G36gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(G64gat), .B(G92gat), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n277), .A2(new_n282), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT79), .ZN(new_n431));
  NAND2_X1  g230(.A1(G226gat), .A2(G233gat), .ZN(new_n432));
  XOR2_X1   g231(.A(new_n432), .B(KEYINPUT78), .Z(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n275), .A2(new_n276), .B1(new_n236), .B2(new_n250), .ZN(new_n435));
  INV_X1    g234(.A(new_n433), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT79), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n436), .B1(new_n435), .B2(KEYINPUT29), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n353), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n430), .A2(new_n433), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(new_n441), .A3(new_n353), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n429), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n433), .B1(new_n430), .B2(new_n356), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n445), .B1(new_n437), .B2(new_n434), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n428), .B(new_n442), .C1(new_n446), .C2(new_n353), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n444), .A2(new_n447), .A3(KEYINPUT30), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n440), .A2(new_n443), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT30), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(new_n450), .A3(new_n428), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n310), .A2(new_n380), .A3(new_n425), .A4(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT76), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n302), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n306), .A2(KEYINPUT76), .A3(new_n299), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n305), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n370), .A2(new_n374), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n375), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n457), .A2(new_n459), .A3(new_n377), .A4(new_n303), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n413), .A2(KEYINPUT6), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n461), .B1(new_n422), .B2(new_n413), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n452), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT35), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n453), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n378), .A2(new_n379), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n395), .B1(new_n410), .B2(new_n411), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT39), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n468), .A3(new_n389), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n384), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT39), .B1(new_n387), .B2(new_n389), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n471), .B1(new_n467), .B2(new_n389), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT40), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n472), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT40), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n474), .A2(new_n475), .A3(new_n384), .A4(new_n469), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n420), .A2(new_n448), .A3(new_n451), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n466), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT38), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT89), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n438), .A2(new_n439), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n353), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n439), .A2(new_n441), .A3(new_n359), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n484), .A2(KEYINPUT37), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n481), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n359), .B1(new_n438), .B2(new_n439), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(KEYINPUT37), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT89), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n480), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n442), .B1(new_n446), .B2(new_n353), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n429), .B1(new_n491), .B2(KEYINPUT37), .ZN(new_n492));
  NOR3_X1   g291(.A1(new_n490), .A2(KEYINPUT90), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT90), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n483), .A2(new_n485), .A3(new_n481), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT89), .B1(new_n487), .B2(new_n488), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT38), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n492), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n493), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT37), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n449), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT38), .B1(new_n492), .B2(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n424), .A2(new_n503), .A3(new_n447), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n479), .B1(new_n500), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n459), .A2(new_n377), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n463), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n295), .A2(new_n296), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n455), .A2(new_n456), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n303), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT36), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT36), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n304), .A2(new_n307), .A3(new_n512), .A4(new_n309), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n507), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n465), .B1(new_n505), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT92), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n371), .A2(G15gat), .ZN(new_n517));
  INV_X1    g316(.A(G15gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(G22gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(G1gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(G8gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(KEYINPUT16), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n517), .A2(new_n519), .A3(new_n524), .ZN(new_n525));
  AND4_X1   g324(.A1(new_n516), .A2(new_n522), .A3(new_n523), .A4(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT92), .B1(new_n520), .B2(new_n521), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n523), .B1(new_n527), .B2(new_n525), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT93), .ZN(new_n530));
  AND2_X1   g329(.A1(G29gat), .A2(G36gat), .ZN(new_n531));
  NOR2_X1   g330(.A1(G29gat), .A2(G36gat), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n531), .B1(KEYINPUT14), .B2(new_n532), .ZN(new_n533));
  OR2_X1    g332(.A1(G43gat), .A2(G50gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT15), .ZN(new_n535));
  NAND2_X1  g334(.A1(G43gat), .A2(G50gat), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AND2_X1   g336(.A1(G43gat), .A2(G50gat), .ZN(new_n538));
  NOR2_X1   g337(.A1(G43gat), .A2(G50gat), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT15), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT14), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(G29gat), .B2(G36gat), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n533), .A2(new_n537), .A3(new_n540), .A4(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(G29gat), .ZN(new_n544));
  INV_X1    g343(.A(G36gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n545), .A3(KEYINPUT14), .ZN(new_n546));
  NAND2_X1  g345(.A1(G29gat), .A2(G36gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(new_n542), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n534), .A2(new_n536), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(KEYINPUT15), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n543), .A2(new_n550), .A3(KEYINPUT17), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n543), .A2(new_n550), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT17), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n529), .A2(new_n530), .A3(new_n551), .A4(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n522), .A2(new_n516), .A3(new_n525), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(G8gat), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n527), .A2(new_n523), .A3(new_n525), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n543), .A2(new_n550), .A3(KEYINPUT17), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT17), .B1(new_n543), .B2(new_n550), .ZN(new_n561));
  NOR3_X1   g360(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n552), .B1(new_n526), .B2(new_n528), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT93), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n555), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G229gat), .A2(G233gat), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(KEYINPUT18), .A3(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n559), .B(new_n552), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT94), .B(KEYINPUT13), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(new_n566), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT18), .B1(new_n565), .B2(new_n566), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT91), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G113gat), .B(G141gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(G197gat), .ZN(new_n576));
  XOR2_X1   g375(.A(KEYINPUT11), .B(G169gat), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT12), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g380(.A(KEYINPUT91), .B(new_n579), .C1(new_n572), .C2(new_n573), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n515), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G134gat), .B(G162gat), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G190gat), .B(G218gat), .Z(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT97), .B(G92gat), .ZN(new_n591));
  INV_X1    g390(.A(G85gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(G85gat), .A2(G92gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT7), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT7), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n595), .A2(G85gat), .A3(G92gat), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n591), .A2(new_n592), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G99gat), .B(G106gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(G99gat), .A2(G106gat), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT96), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(KEYINPUT96), .A2(G99gat), .A3(G106gat), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n601), .A2(KEYINPUT8), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n597), .A2(new_n598), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(G92gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT97), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT97), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(G92gat), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n608), .A3(new_n592), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n596), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n603), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n598), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n552), .A2(new_n604), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AND4_X1   g415(.A1(new_n598), .A2(new_n603), .A3(new_n609), .A4(new_n610), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n598), .B1(new_n597), .B2(new_n603), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n554), .B(new_n551), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n590), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n616), .A2(new_n619), .A3(new_n590), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n588), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n622), .ZN(new_n624));
  INV_X1    g423(.A(new_n588), .ZN(new_n625));
  NOR3_X1   g424(.A1(new_n624), .A2(new_n625), .A3(new_n620), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(G71gat), .A2(G78gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(G71gat), .A2(G78gat), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G57gat), .B(G64gat), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(G57gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(G64gat), .ZN(new_n635));
  INV_X1    g434(.A(G64gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(G57gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G71gat), .B(G78gat), .ZN(new_n639));
  INV_X1    g438(.A(new_n632), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n633), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n642), .B1(new_n618), .B2(new_n617), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n633), .A2(new_n641), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n644), .A2(new_n604), .A3(new_n613), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT98), .B(KEYINPUT10), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n643), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n644), .A2(new_n604), .A3(new_n613), .A4(KEYINPUT10), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G230gat), .A2(G233gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n643), .A2(new_n645), .ZN(new_n652));
  INV_X1    g451(.A(new_n650), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n656), .B(new_n657), .Z(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n655), .A2(new_n659), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT95), .B(KEYINPUT21), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n642), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(G231gat), .A2(G233gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G127gat), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n559), .B1(KEYINPUT21), .B2(new_n644), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(new_n334), .ZN(new_n672));
  XNOR2_X1  g471(.A(G183gat), .B(G211gat), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n672), .B(new_n673), .Z(new_n674));
  OR2_X1    g473(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n670), .A2(new_n674), .ZN(new_n676));
  AOI211_X1 g475(.A(new_n627), .B(new_n663), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n585), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(new_n462), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(new_n521), .ZN(G1324gat));
  NOR2_X1   g479(.A1(new_n678), .A2(new_n452), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(new_n523), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT16), .B(G8gat), .Z(new_n683));
  AND2_X1   g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n682), .B1(new_n684), .B2(KEYINPUT42), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n681), .A2(new_n683), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT99), .B(KEYINPUT42), .Z(new_n687));
  AND3_X1   g486(.A1(new_n686), .A2(KEYINPUT100), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(KEYINPUT100), .B1(new_n686), .B2(new_n687), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n685), .B1(new_n688), .B2(new_n689), .ZN(G1325gat));
  INV_X1    g489(.A(new_n310), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n518), .B1(new_n678), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT101), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n511), .A2(new_n513), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT102), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n511), .A2(new_n513), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n678), .A2(new_n518), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n693), .A2(new_n699), .ZN(G1326gat));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n678), .B2(new_n466), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n585), .A2(KEYINPUT103), .A3(new_n506), .A4(new_n677), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT43), .B(G22gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  INV_X1    g505(.A(new_n663), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n675), .A2(new_n676), .ZN(new_n708));
  INV_X1    g507(.A(new_n627), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n515), .A2(new_n584), .A3(new_n707), .A4(new_n710), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n711), .A2(G29gat), .A3(new_n462), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT45), .Z(new_n713));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(new_n515), .B2(new_n627), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n627), .A2(KEYINPUT104), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n623), .B2(new_n626), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(KEYINPUT44), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n420), .A2(new_n448), .A3(new_n451), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n473), .A2(new_n476), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n506), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(KEYINPUT90), .B1(new_n490), .B2(new_n492), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n498), .A2(new_n497), .A3(new_n494), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n424), .A2(new_n503), .A3(new_n447), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n725), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n511), .A2(new_n513), .A3(new_n696), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n696), .B1(new_n511), .B2(new_n513), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n730), .B(new_n507), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n722), .B1(new_n733), .B2(new_n465), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n715), .A2(new_n734), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n708), .A2(new_n583), .A3(new_n663), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n735), .A2(new_n462), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n713), .B1(new_n544), .B2(new_n738), .ZN(G1328gat));
  INV_X1    g538(.A(new_n452), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n740), .B(new_n736), .C1(new_n715), .C2(new_n734), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G36gat), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n545), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT46), .B1(new_n711), .B2(new_n743), .ZN(new_n744));
  OR3_X1    g543(.A1(new_n711), .A2(KEYINPUT46), .A3(new_n743), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n742), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT105), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1329gat));
  NOR2_X1   g547(.A1(new_n691), .A2(G43gat), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  OR3_X1    g549(.A1(new_n711), .A2(KEYINPUT107), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(KEYINPUT107), .B1(new_n711), .B2(new_n750), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n731), .A2(new_n732), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n754), .B(new_n736), .C1(new_n715), .C2(new_n734), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G43gat), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT47), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT106), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n753), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n755), .A2(KEYINPUT106), .A3(G43gat), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n756), .B(new_n758), .C1(new_n711), .C2(new_n750), .ZN(new_n761));
  AOI22_X1  g560(.A1(new_n759), .A2(new_n760), .B1(new_n761), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g561(.A1(new_n711), .A2(G50gat), .A3(new_n466), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n763), .A2(KEYINPUT109), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n506), .B(new_n736), .C1(new_n715), .C2(new_n734), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G50gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n763), .A2(KEYINPUT109), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n764), .A2(KEYINPUT48), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n765), .A2(new_n769), .A3(G50gat), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n769), .B1(new_n765), .B2(G50gat), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n770), .A2(new_n771), .A3(new_n763), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n768), .B1(new_n772), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g572(.A1(new_n733), .A2(new_n465), .ZN(new_n774));
  INV_X1    g573(.A(new_n708), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n583), .A2(new_n663), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n775), .A2(new_n776), .A3(new_n627), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(new_n462), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(new_n634), .ZN(G1332gat));
  NOR2_X1   g579(.A1(new_n778), .A2(new_n452), .ZN(new_n781));
  NOR2_X1   g580(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n782));
  AND2_X1   g581(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n781), .B2(new_n782), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT110), .ZN(G1333gat));
  OR3_X1    g585(.A1(new_n778), .A2(G71gat), .A3(new_n691), .ZN(new_n787));
  OAI21_X1  g586(.A(G71gat), .B1(new_n778), .B2(new_n698), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n789), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g589(.A1(new_n778), .A2(new_n466), .ZN(new_n791));
  XOR2_X1   g590(.A(new_n791), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n708), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n715), .B2(new_n734), .ZN(new_n794));
  OAI21_X1  g593(.A(G85gat), .B1(new_n794), .B2(new_n462), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n796));
  INV_X1    g595(.A(new_n507), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n503), .A2(new_n447), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n798), .A2(new_n424), .A3(new_n726), .A4(new_n727), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n797), .B1(new_n799), .B2(new_n725), .ZN(new_n800));
  AOI22_X1  g599(.A1(new_n800), .A2(new_n698), .B1(new_n464), .B2(new_n453), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n710), .A2(new_n583), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n796), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n802), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n774), .A2(KEYINPUT51), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT111), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n707), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n807), .B2(new_n806), .ZN(new_n809));
  INV_X1    g608(.A(new_n462), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n592), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n795), .B1(new_n809), .B2(new_n811), .ZN(G1336gat));
  NAND3_X1  g611(.A1(new_n803), .A2(KEYINPUT112), .A3(new_n805), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n814), .B(new_n796), .C1(new_n801), .C2(new_n802), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n452), .A2(G92gat), .A3(new_n707), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n813), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n591), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n794), .B2(new_n452), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT52), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT52), .B1(new_n806), .B2(new_n816), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n819), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(G1337gat));
  OAI21_X1  g623(.A(G99gat), .B1(new_n794), .B2(new_n698), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n691), .A2(G99gat), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n809), .B2(new_n826), .ZN(G1338gat));
  NOR3_X1   g626(.A1(new_n466), .A2(G106gat), .A3(new_n707), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n815), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(G106gat), .B1(new_n794), .B2(new_n466), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT53), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT53), .B1(new_n806), .B2(new_n828), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n833), .A2(new_n834), .A3(new_n830), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n834), .B1(new_n833), .B2(new_n830), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n832), .B1(new_n835), .B2(new_n836), .ZN(G1339gat));
  AOI211_X1 g636(.A(KEYINPUT54), .B(new_n653), .C1(new_n647), .C2(new_n648), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n838), .A2(new_n839), .A3(new_n658), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n649), .A2(new_n841), .A3(new_n650), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT115), .B1(new_n842), .B2(new_n659), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n643), .A2(new_n645), .A3(new_n646), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n648), .A2(new_n653), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT54), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n653), .B1(new_n647), .B2(new_n648), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n846), .A2(KEYINPUT114), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n648), .A2(new_n653), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n841), .B1(new_n850), .B2(new_n647), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n849), .B1(new_n651), .B2(new_n851), .ZN(new_n852));
  OAI22_X1  g651(.A1(new_n840), .A2(new_n843), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT55), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT114), .B1(new_n846), .B2(new_n847), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n651), .A2(new_n851), .A3(new_n849), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n854), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n839), .B1(new_n838), .B2(new_n658), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n842), .A2(KEYINPUT115), .A3(new_n659), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n660), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n855), .A2(new_n862), .A3(new_n581), .A4(new_n582), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n565), .A2(new_n566), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT18), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n866), .A2(new_n571), .A3(new_n567), .A4(new_n579), .ZN(new_n867));
  OAI22_X1  g666(.A1(new_n565), .A2(new_n566), .B1(new_n568), .B2(new_n570), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(KEYINPUT116), .A3(new_n578), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n578), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n663), .A2(new_n867), .A3(new_n869), .A4(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n719), .B1(new_n863), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n872), .A2(new_n867), .A3(new_n869), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n719), .A2(new_n875), .A3(new_n855), .A4(new_n862), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n775), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n677), .A2(new_n583), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n462), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n460), .A2(new_n740), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(G113gat), .B1(new_n882), .B2(new_n584), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n506), .B1(new_n878), .B2(new_n879), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n740), .A2(new_n462), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n884), .A2(new_n310), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n583), .A2(new_n206), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(G1340gat));
  AOI21_X1  g687(.A(G120gat), .B1(new_n882), .B2(new_n663), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n663), .A2(G120gat), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n886), .B2(new_n890), .ZN(G1341gat));
  NAND3_X1  g690(.A1(new_n886), .A2(G127gat), .A3(new_n708), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n892), .A2(KEYINPUT117), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(KEYINPUT117), .ZN(new_n894));
  AOI21_X1  g693(.A(G127gat), .B1(new_n882), .B2(new_n708), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(G1342gat));
  NOR2_X1   g695(.A1(new_n709), .A2(new_n213), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n898), .A2(KEYINPUT56), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n886), .A2(new_n627), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(G134gat), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT118), .B1(new_n898), .B2(KEYINPUT56), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n898), .A2(KEYINPUT118), .A3(KEYINPUT56), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n901), .B(KEYINPUT119), .C1(new_n902), .C2(new_n903), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1343gat));
  NAND2_X1  g707(.A1(new_n698), .A2(new_n885), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n627), .B1(new_n863), .B2(new_n873), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n775), .B1(new_n910), .B2(new_n877), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n911), .A2(KEYINPUT120), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n879), .B1(new_n911), .B2(KEYINPUT120), .ZN(new_n913));
  OAI211_X1 g712(.A(KEYINPUT57), .B(new_n506), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n466), .B1(new_n878), .B2(new_n879), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n915), .A2(KEYINPUT57), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n909), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n584), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G141gat), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT121), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n754), .A2(new_n466), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n921), .A2(new_n880), .A3(new_n452), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n339), .A3(new_n584), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n920), .A2(new_n924), .A3(KEYINPUT58), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT58), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n919), .B(new_n923), .C1(KEYINPUT121), .C2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1344gat));
  NAND3_X1  g727(.A1(new_n922), .A2(new_n341), .A3(new_n663), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n341), .B1(new_n917), .B2(new_n663), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT122), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n506), .A2(KEYINPUT57), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n932), .B1(new_n878), .B2(new_n879), .ZN(new_n933));
  AND4_X1   g732(.A1(new_n627), .A2(new_n875), .A3(new_n855), .A4(new_n862), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n775), .B1(new_n910), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n466), .B1(new_n935), .B2(new_n879), .ZN(new_n936));
  OAI22_X1  g735(.A1(new_n931), .A2(new_n933), .B1(new_n936), .B2(KEYINPUT57), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n933), .A2(new_n931), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AND4_X1   g738(.A1(new_n663), .A2(new_n939), .A3(new_n698), .A4(new_n885), .ZN(new_n940));
  NAND2_X1  g739(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n941));
  OAI221_X1 g740(.A(new_n929), .B1(KEYINPUT59), .B2(new_n930), .C1(new_n940), .C2(new_n941), .ZN(G1345gat));
  INV_X1    g741(.A(new_n917), .ZN(new_n943));
  OAI21_X1  g742(.A(G155gat), .B1(new_n943), .B2(new_n775), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n922), .A2(new_n334), .A3(new_n708), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1346gat));
  OAI21_X1  g745(.A(G162gat), .B1(new_n943), .B2(new_n720), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n922), .A2(new_n335), .A3(new_n627), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(G1347gat));
  NOR2_X1   g748(.A1(new_n810), .A2(new_n452), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT123), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n951), .A2(new_n310), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(new_n884), .ZN(new_n953));
  INV_X1    g752(.A(G169gat), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n953), .A2(new_n954), .A3(new_n583), .ZN(new_n955));
  AOI211_X1 g754(.A(new_n810), .B(new_n452), .C1(new_n878), .C2(new_n879), .ZN(new_n956));
  INV_X1    g755(.A(new_n460), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(new_n584), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n955), .B1(new_n954), .B2(new_n960), .ZN(G1348gat));
  OAI21_X1  g760(.A(G176gat), .B1(new_n953), .B2(new_n707), .ZN(new_n962));
  OR2_X1    g761(.A1(new_n707), .A2(G176gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n958), .B2(new_n963), .ZN(G1349gat));
  NAND4_X1  g763(.A1(new_n959), .A2(new_n228), .A3(new_n230), .A4(new_n708), .ZN(new_n965));
  OAI21_X1  g764(.A(G183gat), .B1(new_n953), .B2(new_n775), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT60), .ZN(new_n967));
  AOI22_X1  g766(.A1(new_n965), .A2(new_n966), .B1(KEYINPUT124), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n967), .A2(KEYINPUT124), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n968), .B(new_n969), .ZN(G1350gat));
  NAND3_X1  g769(.A1(new_n959), .A2(new_n231), .A3(new_n719), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n952), .A2(new_n627), .A3(new_n884), .ZN(new_n972));
  XNOR2_X1  g771(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n972), .A2(G190gat), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n973), .B1(new_n972), .B2(G190gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n971), .B1(new_n974), .B2(new_n975), .ZN(G1351gat));
  AND2_X1   g775(.A1(new_n921), .A2(new_n956), .ZN(new_n977));
  AOI21_X1  g776(.A(G197gat), .B1(new_n977), .B2(new_n584), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n698), .A2(new_n951), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n939), .A2(new_n979), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n584), .A2(G197gat), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(G1352gat));
  NAND3_X1  g781(.A1(new_n939), .A2(new_n663), .A3(new_n979), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(G204gat), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n707), .A2(G204gat), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n921), .A2(new_n956), .A3(new_n985), .ZN(new_n986));
  XOR2_X1   g785(.A(new_n986), .B(KEYINPUT62), .Z(new_n987));
  NAND2_X1  g786(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT126), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n984), .A2(KEYINPUT126), .A3(new_n987), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(G1353gat));
  NAND3_X1  g791(.A1(new_n977), .A2(new_n319), .A3(new_n708), .ZN(new_n993));
  OAI211_X1 g792(.A(new_n708), .B(new_n979), .C1(new_n937), .C2(new_n938), .ZN(new_n994));
  AND3_X1   g793(.A1(new_n994), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n995));
  AOI21_X1  g794(.A(KEYINPUT63), .B1(new_n994), .B2(G211gat), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n993), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI211_X1 g798(.A(KEYINPUT127), .B(new_n993), .C1(new_n995), .C2(new_n996), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(G1354gat));
  AOI21_X1  g800(.A(new_n320), .B1(new_n980), .B2(new_n627), .ZN(new_n1002));
  AND3_X1   g801(.A1(new_n977), .A2(new_n320), .A3(new_n719), .ZN(new_n1003));
  OR2_X1    g802(.A1(new_n1002), .A2(new_n1003), .ZN(G1355gat));
endmodule


