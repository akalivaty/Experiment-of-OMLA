//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1231,
    new_n1232, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n207), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT1), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n207), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT0), .Z(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(new_n201), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n215), .B(new_n218), .C1(new_n221), .C2(new_n224), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT65), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n230), .B(new_n233), .Z(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XNOR2_X1  g0035(.A(G107), .B(G116), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n202), .A2(G68), .ZN(new_n238));
  INV_X1    g0038(.A(G68), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n239), .A2(G50), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n237), .B(new_n243), .ZN(G351));
  NAND2_X1  g0044(.A1(G33), .A2(G41), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n245), .A2(G1), .A3(G13), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n247), .A2(G222), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n247), .A2(G223), .A3(G1698), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G77), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n249), .A2(new_n250), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n246), .B1(new_n257), .B2(KEYINPUT66), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(KEYINPUT66), .B2(new_n257), .ZN(new_n259));
  INV_X1    g0059(.A(new_n246), .ZN(new_n260));
  INV_X1    g0060(.A(G274), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(G41), .B2(G45), .ZN(new_n263));
  NOR3_X1   g0063(.A1(new_n260), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n246), .A2(new_n263), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n264), .B1(G226), .B2(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G190), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n203), .A2(G20), .ZN(new_n269));
  INV_X1    g0069(.A(G150), .ZN(new_n270));
  NOR2_X1   g0070(.A1(G20), .A2(G33), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n269), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n220), .A2(G33), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT68), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n220), .A2(KEYINPUT68), .A3(G33), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT8), .B(G58), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n273), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n219), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT67), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n282), .A2(KEYINPUT67), .A3(new_n219), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n262), .A2(G13), .A3(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n288), .B1(new_n202), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n286), .ZN(new_n292));
  AOI21_X1  g0092(.A(KEYINPUT67), .B1(new_n282), .B2(new_n219), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(new_n290), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n262), .A2(G20), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(G50), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n291), .A2(new_n297), .A3(KEYINPUT9), .ZN(new_n298));
  OAI221_X1 g0098(.A(new_n297), .B1(G50), .B2(new_n289), .C1(new_n287), .C2(new_n281), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT9), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n268), .A2(new_n298), .A3(new_n301), .A4(KEYINPUT70), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n268), .A2(new_n298), .A3(new_n301), .ZN(new_n305));
  INV_X1    g0105(.A(G200), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n267), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n302), .B(new_n303), .C1(new_n305), .C2(new_n307), .ZN(new_n310));
  INV_X1    g0110(.A(G179), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n267), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n299), .B1(new_n267), .B2(G169), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n309), .A2(new_n310), .A3(new_n315), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n252), .A2(new_n254), .A3(G232), .A4(G1698), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n252), .A2(new_n254), .A3(G226), .A4(new_n248), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G97), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n260), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT13), .ZN(new_n322));
  INV_X1    g0122(.A(new_n263), .ZN(new_n323));
  INV_X1    g0123(.A(new_n219), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n261), .B1(new_n324), .B2(new_n245), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n265), .A2(G238), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n321), .A2(new_n322), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n322), .B1(new_n321), .B2(new_n326), .ZN(new_n328));
  OAI21_X1  g0128(.A(G169), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT14), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g0131(.A(KEYINPUT14), .B(G169), .C1(new_n327), .C2(new_n328), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n321), .A2(new_n322), .A3(new_n326), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT72), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT72), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n321), .A2(new_n326), .A3(new_n336), .A4(new_n322), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n328), .A2(new_n311), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n333), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n276), .A2(G77), .A3(new_n277), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n271), .A2(G50), .B1(G20), .B2(new_n239), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n294), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT73), .B(KEYINPUT11), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n344), .A2(new_n294), .A3(new_n346), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OR3_X1    g0150(.A1(new_n289), .A2(KEYINPUT74), .A3(G68), .ZN(new_n351));
  OAI21_X1  g0151(.A(KEYINPUT74), .B1(new_n289), .B2(G68), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(KEYINPUT12), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n239), .B1(new_n262), .B2(G20), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n289), .B(new_n354), .C1(new_n292), .C2(new_n293), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT12), .ZN(new_n356));
  OAI211_X1 g0156(.A(KEYINPUT74), .B(new_n356), .C1(new_n289), .C2(G68), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n353), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT75), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n353), .A2(new_n355), .A3(KEYINPUT75), .A4(new_n357), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n350), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n341), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n280), .B1(KEYINPUT69), .B2(new_n271), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(KEYINPUT69), .B2(new_n271), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT15), .B(G87), .ZN(new_n366));
  INV_X1    g0166(.A(G77), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n366), .A2(new_n274), .B1(new_n220), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n294), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n295), .A2(G77), .A3(new_n296), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n369), .B(new_n370), .C1(G77), .C2(new_n289), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n247), .A2(G232), .A3(new_n248), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n247), .A2(G238), .A3(G1698), .ZN(new_n373));
  INV_X1    g0173(.A(G107), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n372), .B(new_n373), .C1(new_n374), .C2(new_n247), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n260), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n264), .B1(G244), .B2(new_n265), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(new_n377), .A3(new_n311), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n377), .ZN(new_n379));
  INV_X1    g0179(.A(G169), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n371), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n371), .B1(G200), .B2(new_n379), .ZN(new_n383));
  INV_X1    g0183(.A(G190), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n383), .B1(new_n384), .B2(new_n379), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n328), .A2(new_n384), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n362), .B1(new_n338), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(G200), .B1(new_n327), .B2(new_n328), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT71), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g0190(.A(KEYINPUT71), .B(G200), .C1(new_n327), .C2(new_n328), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n363), .A2(new_n382), .A3(new_n385), .A4(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n316), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT7), .B1(new_n255), .B2(new_n220), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  AOI211_X1 g0197(.A(new_n397), .B(G20), .C1(new_n252), .C2(new_n254), .ZN(new_n398));
  OAI21_X1  g0198(.A(G68), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n271), .A2(G159), .ZN(new_n400));
  INV_X1    g0200(.A(G58), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n401), .A2(new_n239), .ZN(new_n402));
  OAI21_X1  g0202(.A(G20), .B1(new_n402), .B2(new_n201), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n399), .A2(KEYINPUT16), .A3(new_n400), .A4(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT16), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n397), .B1(new_n247), .B2(G20), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n255), .A2(KEYINPUT7), .A3(new_n220), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n239), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n403), .A2(new_n400), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n405), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n404), .A2(new_n410), .A3(new_n294), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n279), .B1(new_n262), .B2(G20), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n295), .A2(new_n412), .B1(new_n279), .B2(new_n290), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n252), .A2(new_n254), .A3(G226), .A4(G1698), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n252), .A2(new_n254), .A3(G223), .A4(new_n248), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G33), .A2(G87), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n260), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n265), .A2(G232), .B1(new_n323), .B2(new_n325), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n418), .A2(G190), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n419), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G200), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n411), .A2(new_n413), .A3(new_n420), .A4(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT17), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n423), .B(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n418), .A2(new_n311), .A3(new_n419), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT76), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT76), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n418), .A2(new_n419), .A3(new_n428), .A4(new_n311), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n421), .A2(new_n380), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n427), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n411), .A2(new_n413), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(new_n432), .A3(KEYINPUT18), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT77), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n431), .A2(new_n432), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT18), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n436), .A2(new_n434), .A3(new_n437), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n425), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n395), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT78), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT6), .ZN(new_n444));
  AND2_X1   g0244(.A1(G97), .A2(G107), .ZN(new_n445));
  NOR2_X1   g0245(.A1(G97), .A2(G107), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(KEYINPUT6), .A2(G97), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(G107), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n220), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n272), .A2(new_n367), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n443), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(G107), .B1(new_n396), .B2(new_n398), .ZN(new_n454));
  INV_X1    g0254(.A(new_n452), .ZN(new_n455));
  XNOR2_X1  g0255(.A(G97), .B(G107), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n449), .B1(new_n456), .B2(new_n444), .ZN(new_n457));
  OAI211_X1 g0257(.A(KEYINPUT78), .B(new_n455), .C1(new_n457), .C2(new_n220), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n453), .A2(new_n454), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n294), .ZN(new_n460));
  INV_X1    g0260(.A(G97), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n290), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n262), .A2(G33), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n287), .A2(new_n289), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n462), .B1(new_n464), .B2(new_n461), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n460), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G45), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(G1), .ZN(new_n469));
  AND2_X1   g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  NOR2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n472), .A2(new_n260), .A3(new_n261), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n472), .A2(G257), .A3(new_n246), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n252), .A2(new_n254), .A3(G244), .A4(new_n248), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT4), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n247), .A2(KEYINPUT4), .A3(G244), .A4(new_n248), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G283), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n247), .A2(G250), .A3(G1698), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n477), .A2(new_n478), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  AOI211_X1 g0281(.A(new_n473), .B(new_n474), .C1(new_n481), .C2(new_n260), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n311), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n260), .ZN(new_n484));
  XNOR2_X1  g0284(.A(KEYINPUT5), .B(G41), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n325), .A2(new_n469), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n474), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n380), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n467), .A2(new_n483), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(G200), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n465), .B1(new_n459), .B2(new_n294), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n474), .B1(new_n481), .B2(new_n260), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(G190), .A3(new_n486), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n287), .A2(G87), .A3(new_n289), .A4(new_n463), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT19), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n220), .B1(new_n319), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(G87), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n446), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n252), .A2(new_n254), .A3(new_n220), .A4(G68), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n497), .B1(new_n274), .B2(new_n461), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n294), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n366), .A2(new_n290), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n496), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n246), .A2(G274), .A3(new_n469), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n262), .A2(G45), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n246), .A2(G250), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n252), .A2(new_n254), .A3(G244), .A4(G1698), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n252), .A2(new_n254), .A3(G238), .A4(new_n248), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G116), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n511), .B1(new_n260), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G190), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n507), .B(new_n517), .C1(new_n306), .C2(new_n516), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n515), .A2(new_n260), .ZN(new_n519));
  INV_X1    g0319(.A(new_n511), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(G179), .A3(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n380), .B2(new_n516), .ZN(new_n522));
  INV_X1    g0322(.A(new_n366), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n287), .A2(new_n289), .A3(new_n523), .A4(new_n463), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n524), .A2(new_n505), .A3(new_n506), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT79), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT79), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n524), .A2(new_n505), .A3(new_n527), .A4(new_n506), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n522), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  AND4_X1   g0329(.A1(new_n490), .A2(new_n495), .A3(new_n518), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n255), .A2(G303), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n252), .A2(new_n254), .A3(G257), .A4(new_n248), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n252), .A2(new_n254), .A3(G264), .A4(G1698), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT80), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT80), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n531), .A2(new_n536), .A3(new_n532), .A4(new_n533), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n260), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n472), .A2(new_n246), .ZN(new_n539));
  INV_X1    g0339(.A(G270), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n486), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n538), .A2(G190), .A3(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n479), .B(new_n220), .C1(G33), .C2(new_n461), .ZN(new_n544));
  INV_X1    g0344(.A(G116), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G20), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n283), .A3(new_n546), .ZN(new_n547));
  OR2_X1    g0347(.A1(KEYINPUT81), .A2(KEYINPUT20), .ZN(new_n548));
  OR2_X1    g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  XOR2_X1   g0349(.A(KEYINPUT81), .B(KEYINPUT20), .Z(new_n550));
  AOI22_X1  g0350(.A1(new_n547), .A2(new_n550), .B1(new_n545), .B2(new_n290), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n549), .B(new_n551), .C1(new_n464), .C2(new_n545), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n246), .B1(new_n534), .B2(KEYINPUT80), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n541), .B1(new_n554), .B2(new_n537), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n543), .B(new_n553), .C1(new_n306), .C2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT21), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n552), .A2(G169), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n557), .B1(new_n558), .B2(new_n555), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n555), .A2(G179), .A3(new_n552), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n538), .A2(new_n542), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n561), .A2(KEYINPUT21), .A3(G169), .A4(new_n552), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n556), .A2(new_n559), .A3(new_n560), .A4(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n464), .A2(new_n374), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n290), .A2(new_n374), .ZN(new_n566));
  XNOR2_X1  g0366(.A(new_n566), .B(KEYINPUT25), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g0368(.A(KEYINPUT82), .B(KEYINPUT22), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n247), .A2(new_n569), .A3(new_n220), .A4(G87), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n252), .A2(new_n254), .A3(new_n220), .A4(G87), .ZN(new_n571));
  XOR2_X1   g0371(.A(KEYINPUT82), .B(KEYINPUT22), .Z(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n514), .A2(G20), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT23), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n220), .B2(G107), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n374), .A2(KEYINPUT23), .A3(G20), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n570), .A2(new_n573), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT24), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT24), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n570), .A2(new_n573), .A3(new_n581), .A4(new_n578), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(KEYINPUT83), .B1(new_n583), .B2(new_n294), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT83), .ZN(new_n585));
  AOI211_X1 g0385(.A(new_n585), .B(new_n287), .C1(new_n580), .C2(new_n582), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n568), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(G264), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n486), .B1(new_n539), .B2(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n252), .A2(new_n254), .A3(G257), .A4(G1698), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT84), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n247), .A2(KEYINPUT84), .A3(G257), .A4(G1698), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n252), .A2(new_n254), .A3(G250), .A4(new_n248), .ZN(new_n595));
  NAND2_X1  g0395(.A1(G33), .A2(G294), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n589), .B1(new_n599), .B2(new_n260), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(G179), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n472), .A2(new_n246), .ZN(new_n602));
  INV_X1    g0402(.A(new_n472), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n602), .A2(G264), .B1(new_n603), .B2(new_n325), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n597), .B1(new_n592), .B2(new_n593), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n604), .B1(new_n605), .B2(new_n246), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G169), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n601), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n587), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n604), .B(new_n384), .C1(new_n605), .C2(new_n246), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n600), .B2(G200), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n611), .B(new_n568), .C1(new_n584), .C2(new_n586), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n530), .A2(new_n564), .A3(new_n609), .A4(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n442), .A2(new_n613), .ZN(G372));
  INV_X1    g0414(.A(new_n433), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT18), .B1(new_n431), .B2(new_n432), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n386), .A2(new_n335), .A3(new_n337), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n350), .A2(new_n360), .A3(new_n361), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n620), .B1(new_n390), .B2(new_n391), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n363), .B1(new_n382), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n425), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n617), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n309), .A2(new_n310), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n315), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  XOR2_X1   g0426(.A(new_n626), .B(KEYINPUT86), .Z(new_n627));
  INV_X1    g0427(.A(new_n442), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n529), .A2(new_n518), .ZN(new_n629));
  OAI21_X1  g0429(.A(KEYINPUT26), .B1(new_n490), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n522), .A2(new_n525), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n306), .B1(new_n519), .B2(new_n520), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(G190), .B2(new_n516), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n633), .A2(new_n507), .B1(new_n525), .B2(new_n522), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n460), .A2(new_n466), .B1(new_n482), .B2(new_n311), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT26), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n634), .A2(new_n635), .A3(new_n636), .A4(new_n489), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n630), .A2(new_n631), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT85), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n612), .A2(new_n490), .A3(new_n495), .A4(new_n634), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n562), .A2(new_n560), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n609), .A2(new_n559), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n630), .A2(new_n637), .A3(KEYINPUT85), .A4(new_n631), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n640), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n628), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n627), .A2(new_n648), .ZN(G369));
  NAND3_X1  g0449(.A1(new_n262), .A2(new_n220), .A3(G13), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n553), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n563), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n559), .A2(new_n562), .A3(new_n560), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(new_n657), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G330), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT87), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n609), .A2(new_n656), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n664), .A2(KEYINPUT88), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(KEYINPUT88), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n568), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n220), .A2(G33), .A3(G116), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n374), .A2(KEYINPUT23), .A3(G20), .ZN(new_n670));
  AOI21_X1  g0470(.A(KEYINPUT23), .B1(new_n374), .B2(G20), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n672), .B1(new_n571), .B2(new_n572), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n581), .B1(new_n673), .B2(new_n570), .ZN(new_n674));
  INV_X1    g0474(.A(new_n582), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n294), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n585), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n583), .A2(KEYINPUT83), .A3(new_n294), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n668), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n608), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n612), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n587), .A2(new_n655), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n667), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n663), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n609), .A2(new_n655), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n659), .A2(new_n656), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n687), .B1(new_n685), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n686), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n216), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n500), .A2(G116), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n693), .A2(new_n262), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n224), .B2(new_n693), .ZN(new_n697));
  XOR2_X1   g0497(.A(new_n697), .B(KEYINPUT28), .Z(new_n698));
  INV_X1    g0498(.A(KEYINPUT30), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n600), .A2(new_n493), .A3(new_n516), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n555), .A2(G179), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n516), .B(new_n604), .C1(new_n246), .C2(new_n605), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  AOI211_X1 g0504(.A(new_n311), .B(new_n541), .C1(new_n554), .C2(new_n537), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n704), .A2(new_n705), .A3(KEYINPUT30), .A4(new_n493), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n600), .A2(G179), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n519), .A2(KEYINPUT89), .A3(new_n520), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT89), .B1(new_n519), .B2(new_n520), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n707), .A2(new_n710), .A3(new_n561), .A4(new_n488), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n702), .A2(new_n706), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n655), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT31), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT90), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n712), .A2(KEYINPUT31), .A3(new_n655), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n613), .B2(new_n655), .ZN(new_n718));
  OAI21_X1  g0518(.A(G330), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n638), .A2(new_n639), .B1(new_n642), .B2(new_n644), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n655), .B1(new_n721), .B2(new_n646), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT91), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n647), .A2(new_n656), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT91), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT29), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n723), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n659), .B1(new_n608), .B2(new_n587), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n641), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n467), .A2(new_n489), .A3(new_n483), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(new_n636), .A3(new_n518), .A4(new_n529), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n518), .A2(new_n631), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT26), .B1(new_n490), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n732), .A2(new_n631), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n656), .B1(new_n730), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(KEYINPUT92), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT92), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n738), .B(new_n656), .C1(new_n730), .C2(new_n735), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT29), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n720), .B1(new_n728), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n698), .B1(new_n742), .B2(G1), .ZN(G364));
  INV_X1    g0543(.A(new_n693), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n220), .A2(G13), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n262), .B1(new_n745), .B2(G45), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT93), .Z(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n219), .B1(G20), .B2(new_n380), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(G20), .A2(G179), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT95), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n754), .A2(new_n384), .A3(G200), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n755), .A2(KEYINPUT97), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(KEYINPUT97), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G68), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n220), .A2(G179), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n761), .A2(new_n384), .A3(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G190), .A2(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n754), .A2(new_n763), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n247), .B1(new_n374), .B2(new_n762), .C1(new_n764), .C2(new_n367), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n384), .A2(G200), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n754), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n765), .B1(G58), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n754), .A2(G190), .A3(G200), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G50), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n766), .A2(new_n311), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n461), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n761), .A2(new_n763), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  XOR2_X1   g0577(.A(KEYINPUT96), .B(KEYINPUT32), .Z(new_n778));
  AND3_X1   g0578(.A1(new_n777), .A2(G159), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n778), .B1(new_n777), .B2(G159), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n761), .A2(G190), .A3(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n499), .ZN(new_n782));
  NOR4_X1   g0582(.A1(new_n775), .A2(new_n779), .A3(new_n780), .A4(new_n782), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n760), .A2(new_n768), .A3(new_n771), .A4(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n767), .ZN(new_n785));
  INV_X1    g0585(.A(G322), .ZN(new_n786));
  INV_X1    g0586(.A(G311), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n785), .A2(new_n786), .B1(new_n787), .B2(new_n764), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n247), .B1(new_n777), .B2(G329), .ZN(new_n789));
  INV_X1    g0589(.A(G283), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n789), .B1(new_n790), .B2(new_n762), .ZN(new_n791));
  INV_X1    g0591(.A(G294), .ZN(new_n792));
  INV_X1    g0592(.A(G303), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n774), .A2(new_n792), .B1(new_n781), .B2(new_n793), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n788), .A2(new_n791), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n770), .A2(G326), .ZN(new_n796));
  XOR2_X1   g0596(.A(KEYINPUT33), .B(G317), .Z(new_n797));
  OAI211_X1 g0597(.A(new_n795), .B(new_n796), .C1(new_n758), .C2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n751), .B1(new_n784), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G13), .A2(G33), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G20), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n750), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT94), .Z(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n216), .A2(G355), .A3(new_n247), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n692), .A2(new_n247), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(G45), .B2(new_n223), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n243), .A2(new_n468), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n806), .B1(G116), .B2(new_n216), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n749), .B(new_n799), .C1(new_n805), .C2(new_n810), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT98), .Z(new_n812));
  INV_X1    g0612(.A(new_n661), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n802), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT87), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n662), .B(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n747), .ZN(new_n817));
  INV_X1    g0617(.A(G330), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(new_n813), .B2(new_n818), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n812), .A2(new_n814), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G396));
  NAND2_X1  g0621(.A1(new_n371), .A2(new_n655), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n385), .A2(new_n382), .A3(new_n822), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n371), .A2(new_n378), .A3(new_n381), .A4(new_n655), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT101), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n723), .A2(new_n726), .A3(KEYINPUT103), .A4(new_n827), .ZN(new_n828));
  AND3_X1   g0628(.A1(new_n723), .A2(new_n726), .A3(new_n827), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n647), .A2(new_n656), .A3(new_n826), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT103), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n828), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n720), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n828), .B(new_n719), .C1(new_n829), .C2(new_n832), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n834), .A2(new_n747), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n751), .A2(new_n801), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n748), .B1(G77), .B2(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT99), .Z(new_n839));
  OAI22_X1  g0639(.A1(new_n785), .A2(new_n792), .B1(new_n545), .B2(new_n764), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n255), .B1(new_n776), .B2(new_n787), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n499), .A2(new_n762), .B1(new_n781), .B2(new_n374), .ZN(new_n842));
  NOR4_X1   g0642(.A1(new_n840), .A2(new_n775), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n793), .B2(new_n769), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(G283), .B2(new_n759), .ZN(new_n845));
  INV_X1    g0645(.A(new_n764), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(G159), .ZN(new_n847));
  INV_X1    g0647(.A(G137), .ZN(new_n848));
  XNOR2_X1  g0648(.A(KEYINPUT100), .B(G143), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n847), .B1(new_n848), .B2(new_n769), .C1(new_n785), .C2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G150), .B2(new_n759), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT34), .Z(new_n852));
  INV_X1    g0652(.A(G132), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n247), .B1(new_n776), .B2(new_n853), .C1(new_n774), .C2(new_n401), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n202), .A2(new_n781), .B1(new_n762), .B2(new_n239), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n845), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n839), .B1(new_n801), .B2(new_n826), .C1(new_n857), .C2(new_n751), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT102), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n836), .A2(new_n859), .ZN(G384));
  INV_X1    g0660(.A(new_n457), .ZN(new_n861));
  OR2_X1    g0661(.A1(new_n861), .A2(KEYINPUT35), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(KEYINPUT35), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n862), .A2(new_n863), .A3(G116), .A4(new_n221), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n864), .B(KEYINPUT36), .Z(new_n865));
  OR3_X1    g0665(.A1(new_n223), .A2(new_n367), .A3(new_n402), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n262), .B(G13), .C1(new_n866), .C2(new_n238), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n436), .A2(new_n423), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n653), .B1(new_n411), .B2(new_n413), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT37), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n653), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n432), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT105), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT105), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n874), .A2(new_n423), .A3(new_n436), .A4(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n871), .B1(new_n877), .B2(KEYINPUT37), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n441), .B2(new_n873), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT40), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n878), .B(KEYINPUT38), .C1(new_n441), .C2(new_n873), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n619), .A2(new_n656), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n621), .B2(new_n341), .ZN(new_n886));
  INV_X1    g0686(.A(new_n885), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n331), .A2(new_n332), .B1(new_n338), .B2(new_n339), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n393), .B(new_n887), .C1(new_n619), .C2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n886), .A2(new_n889), .A3(KEYINPUT104), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT104), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n363), .A2(new_n891), .A3(new_n393), .A4(new_n887), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n890), .A2(new_n826), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n715), .A2(new_n717), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n490), .A2(new_n495), .A3(new_n518), .A4(new_n529), .ZN(new_n895));
  NOR4_X1   g0695(.A1(new_n681), .A2(new_n895), .A3(new_n563), .A4(new_n655), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g0697(.A1(KEYINPUT106), .A2(KEYINPUT40), .ZN(new_n898));
  NOR3_X1   g0698(.A1(new_n893), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n884), .A2(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n717), .B(new_n715), .C1(new_n613), .C2(new_n655), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n901), .A2(new_n826), .A3(new_n890), .A4(new_n892), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n870), .A2(new_n875), .ZN(new_n903));
  AOI211_X1 g0703(.A(KEYINPUT105), .B(new_n653), .C1(new_n411), .C2(new_n413), .ZN(new_n904));
  OAI22_X1  g0704(.A1(new_n617), .A2(new_n425), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n877), .A2(KEYINPUT37), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n903), .A2(new_n904), .ZN(new_n908));
  INV_X1    g0708(.A(new_n869), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n905), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n880), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n902), .A2(KEYINPUT106), .B1(new_n912), .B2(new_n883), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n900), .B1(new_n913), .B2(new_n882), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT107), .ZN(new_n915));
  OR3_X1    g0715(.A1(new_n915), .A2(new_n442), .A3(new_n897), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n915), .B1(new_n442), .B2(new_n897), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n916), .A2(G330), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n728), .A2(new_n628), .A3(new_n741), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n627), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n912), .A2(new_n883), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT39), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n363), .A2(new_n655), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n881), .A2(KEYINPUT39), .A3(new_n883), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n890), .A2(new_n892), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n382), .A2(new_n655), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n927), .B1(new_n830), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n881), .A2(new_n883), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n930), .A2(new_n931), .B1(new_n617), .B2(new_n653), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n926), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n920), .B(new_n933), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n918), .A2(new_n934), .B1(new_n262), .B2(new_n745), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT108), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n918), .A2(new_n934), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n935), .A2(KEYINPUT108), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n868), .B1(new_n938), .B2(new_n939), .ZN(G367));
  OAI21_X1  g0740(.A(new_n803), .B1(new_n216), .B2(new_n366), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n807), .B2(new_n233), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n749), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n802), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n634), .B1(new_n507), .B2(new_n656), .ZN(new_n945));
  OR3_X1    g0745(.A1(new_n631), .A2(new_n507), .A3(new_n656), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n785), .A2(new_n270), .B1(new_n202), .B2(new_n764), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n774), .A2(new_n239), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n247), .B1(new_n776), .B2(new_n848), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n401), .A2(new_n781), .B1(new_n762), .B2(new_n367), .ZN(new_n951));
  NOR4_X1   g0751(.A1(new_n948), .A2(new_n949), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(G159), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n952), .B1(new_n769), .B2(new_n849), .C1(new_n953), .C2(new_n758), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n762), .A2(new_n461), .ZN(new_n955));
  INV_X1    g0755(.A(G317), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n255), .B1(new_n776), .B2(new_n956), .C1(new_n774), .C2(new_n374), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n955), .B(new_n957), .C1(new_n770), .C2(G311), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n781), .A2(new_n545), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n959), .A2(KEYINPUT46), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n764), .A2(new_n790), .B1(new_n959), .B2(KEYINPUT46), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n960), .B(new_n961), .C1(G303), .C2(new_n767), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n958), .B(new_n962), .C1(new_n792), .C2(new_n758), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n954), .A2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT47), .Z(new_n965));
  OAI221_X1 g0765(.A(new_n943), .B1(new_n944), .B2(new_n947), .C1(new_n965), .C2(new_n751), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n665), .A2(new_n666), .B1(new_n682), .B2(new_n683), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(new_n688), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n490), .B(new_n495), .C1(new_n492), .C2(new_n656), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n731), .A2(new_n655), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n972), .A2(KEYINPUT42), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n490), .B1(new_n969), .B2(new_n609), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n972), .A2(KEYINPUT42), .B1(new_n656), .B2(new_n974), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n973), .A2(new_n975), .B1(KEYINPUT43), .B2(new_n947), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n976), .B(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n686), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n971), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n978), .B(new_n980), .Z(new_n981));
  XOR2_X1   g0781(.A(new_n746), .B(KEYINPUT109), .Z(new_n982));
  NAND2_X1  g0782(.A1(new_n690), .A2(new_n971), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT45), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n690), .A2(KEYINPUT45), .A3(new_n971), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT44), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n690), .B2(new_n971), .ZN(new_n989));
  INV_X1    g0789(.A(new_n971), .ZN(new_n990));
  OAI211_X1 g0790(.A(KEYINPUT44), .B(new_n990), .C1(new_n968), .C2(new_n687), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n987), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n979), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n685), .A2(new_n689), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n967), .A2(new_n688), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(new_n663), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n742), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n987), .A2(new_n686), .A3(new_n992), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n994), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n742), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n693), .B(KEYINPUT41), .Z(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n982), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n966), .B1(new_n981), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT110), .ZN(G387));
  NAND2_X1  g0808(.A1(new_n967), .A2(new_n802), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n807), .B1(new_n230), .B2(new_n468), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n216), .A2(new_n247), .A3(new_n695), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OR3_X1    g0812(.A1(new_n279), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1013));
  OAI21_X1  g0813(.A(KEYINPUT50), .B1(new_n279), .B2(G50), .ZN(new_n1014));
  AOI21_X1  g0814(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1013), .A2(new_n694), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1012), .A2(new_n1016), .B1(new_n374), .B2(new_n692), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n748), .B1(new_n1017), .B2(new_n804), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n758), .A2(new_n279), .B1(new_n239), .B2(new_n764), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT112), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n247), .B1(new_n762), .B2(new_n461), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n774), .A2(new_n366), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(G50), .C2(new_n767), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n781), .A2(new_n367), .B1(new_n776), .B2(new_n270), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1024), .A2(KEYINPUT111), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n770), .A2(G159), .B1(KEYINPUT111), .B2(new_n1024), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1020), .A2(new_n1023), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT113), .Z(new_n1028));
  AOI21_X1  g0828(.A(new_n247), .B1(new_n777), .B2(G326), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G303), .A2(new_n846), .B1(new_n767), .B2(G317), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n786), .B2(new_n769), .C1(new_n758), .C2(new_n787), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT48), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n781), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G294), .A2(new_n1035), .B1(new_n773), .B2(G283), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1033), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT114), .Z(new_n1038));
  INV_X1    g0838(.A(KEYINPUT49), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1029), .B1(new_n545), .B2(new_n762), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1028), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1018), .B1(new_n1042), .B2(new_n750), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1009), .A2(new_n1043), .B1(new_n998), .B2(new_n982), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n999), .A2(new_n693), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n998), .A2(new_n742), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(G393));
  AND3_X1   g0847(.A1(new_n987), .A2(new_n686), .A3(new_n992), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n686), .B1(new_n987), .B2(new_n992), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n990), .A2(new_n802), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n237), .A2(new_n692), .A3(new_n247), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n803), .B1(new_n216), .B2(new_n461), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n748), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n785), .A2(new_n787), .B1(new_n956), .B2(new_n769), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT52), .Z(new_n1056));
  OAI221_X1 g0856(.A(new_n255), .B1(new_n776), .B2(new_n786), .C1(new_n374), .C2(new_n762), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n774), .A2(new_n545), .B1(new_n781), .B2(new_n790), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(G294), .C2(new_n846), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n758), .B2(new_n793), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n785), .A2(new_n953), .B1(new_n270), .B2(new_n769), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT51), .Z(new_n1062));
  OAI221_X1 g0862(.A(new_n247), .B1(new_n776), .B2(new_n849), .C1(new_n499), .C2(new_n762), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n774), .A2(new_n367), .B1(new_n781), .B2(new_n239), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(new_n280), .C2(new_n846), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n758), .B2(new_n202), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n1056), .A2(new_n1060), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1054), .B1(new_n1067), .B2(new_n750), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1050), .A2(new_n982), .B1(new_n1051), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n999), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1070), .A2(new_n1002), .A3(new_n693), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(KEYINPUT115), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT115), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1069), .A2(new_n1071), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1075), .ZN(G390));
  INV_X1    g0876(.A(new_n927), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n827), .B1(new_n737), .B2(new_n739), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1077), .B1(new_n1078), .B2(new_n928), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n924), .B1(new_n912), .B2(new_n883), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AND3_X1   g0881(.A1(new_n881), .A2(KEYINPUT39), .A3(new_n883), .ZN(new_n1082));
  AOI21_X1  g0882(.A(KEYINPUT39), .B1(new_n912), .B2(new_n883), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n1082), .A2(new_n1083), .B1(new_n930), .B2(new_n924), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n720), .A2(new_n826), .A3(new_n1077), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1081), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n923), .A2(new_n925), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n928), .B1(new_n722), .B2(new_n826), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n1088), .A2(new_n927), .B1(new_n363), .B2(new_n655), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1087), .A2(new_n1089), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n897), .A2(new_n818), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1091), .A2(new_n826), .A3(new_n1077), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1086), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n982), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1087), .A2(new_n800), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n748), .B1(new_n280), .B2(new_n837), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(KEYINPUT54), .B(G143), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n785), .A2(new_n853), .B1(new_n764), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n255), .B1(new_n777), .B2(G125), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n202), .B2(new_n762), .C1(new_n953), .C2(new_n774), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n781), .A2(new_n270), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT53), .ZN(new_n1104));
  INV_X1    g0904(.A(G128), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1102), .B(new_n1104), .C1(new_n1105), .C2(new_n769), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n758), .A2(new_n848), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n758), .A2(new_n374), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n247), .B(new_n782), .C1(G294), .C2(new_n777), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(G97), .A2(new_n846), .B1(new_n767), .B2(G116), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n770), .A2(G283), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n762), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G68), .A2(new_n1112), .B1(new_n773), .B2(G77), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .A4(new_n1113), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n1106), .A2(new_n1107), .B1(new_n1108), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1097), .B1(new_n1115), .B2(new_n750), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1095), .B1(new_n1096), .B2(new_n1116), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n628), .A2(new_n1091), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n627), .A2(new_n919), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1091), .A2(new_n826), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n927), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1078), .A2(new_n928), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n1085), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n927), .B1(new_n719), .B2(new_n827), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n1092), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1088), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1126), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1118), .A2(new_n1086), .A3(new_n1121), .A4(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1125), .A2(new_n1085), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1093), .B1(new_n1120), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1132), .A2(new_n693), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1117), .A2(new_n1135), .ZN(G378));
  OAI21_X1  g0936(.A(KEYINPUT106), .B1(new_n893), .B2(new_n897), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n921), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1138), .A2(KEYINPUT40), .B1(new_n884), .B2(new_n899), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n299), .A2(new_n872), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n316), .A2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n309), .A2(new_n310), .A3(new_n315), .A4(new_n1140), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1144), .B(new_n1145), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n1139), .A2(new_n1146), .A3(new_n818), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1145), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1144), .B(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n914), .B2(G330), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n933), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1146), .B1(new_n1139), .B2(new_n818), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n914), .A2(G330), .A3(new_n1149), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1152), .A2(new_n1153), .A3(new_n926), .A4(new_n932), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1121), .B1(new_n1093), .B2(new_n1133), .ZN(new_n1156));
  AOI21_X1  g0956(.A(KEYINPUT57), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n1157), .A2(KEYINPUT120), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT120), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1159), .B(KEYINPUT57), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1155), .A2(new_n1156), .A3(KEYINPUT57), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1158), .A2(new_n1161), .A3(new_n693), .A4(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n767), .A2(G107), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT116), .Z(new_n1165));
  INV_X1    g0965(.A(G41), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1166), .B(new_n255), .C1(new_n776), .C2(new_n790), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n949), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n762), .A2(new_n401), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G77), .B2(new_n1035), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1168), .B(new_n1170), .C1(new_n545), .C2(new_n769), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1165), .A2(new_n1171), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n759), .A2(G97), .B1(new_n523), .B2(new_n846), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(KEYINPUT117), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1174), .A2(KEYINPUT117), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1172), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  XOR2_X1   g0978(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(G33), .A2(G41), .ZN(new_n1181));
  AOI211_X1 g0981(.A(G50), .B(new_n1181), .C1(new_n255), .C2(new_n1166), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1098), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1035), .A2(new_n1183), .B1(new_n773), .B2(G150), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n848), .B2(new_n764), .C1(new_n785), .C2(new_n1105), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G125), .B2(new_n770), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n853), .B2(new_n758), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1188));
  INV_X1    g0988(.A(G124), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1181), .B1(new_n776), .B2(new_n1189), .C1(new_n953), .C2(new_n762), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n1187), .B2(KEYINPUT59), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1182), .B1(new_n1188), .B2(new_n1191), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1180), .A2(new_n1192), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n751), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n817), .B1(G50), .B2(new_n837), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(new_n1146), .C2(new_n800), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT119), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n982), .B2(new_n1155), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1163), .A2(new_n1199), .ZN(G375));
  OAI21_X1  g1000(.A(new_n748), .B1(G68), .B2(new_n837), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n758), .A2(new_n545), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1022), .B1(G97), .B2(new_n1035), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n770), .A2(G294), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n255), .B1(new_n776), .B2(new_n793), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G77), .B2(new_n1112), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G107), .A2(new_n846), .B1(new_n767), .B2(G283), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1203), .A2(new_n1204), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n758), .A2(new_n1098), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n255), .B(new_n1169), .C1(G128), .C2(new_n777), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G150), .A2(new_n846), .B1(new_n767), .B2(G137), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n770), .A2(G132), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G159), .A2(new_n1035), .B1(new_n773), .B2(G50), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n1202), .A2(new_n1208), .B1(new_n1209), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1201), .B1(new_n1215), .B2(new_n750), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n1077), .B2(new_n801), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n1133), .B2(new_n1094), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1005), .B1(new_n1133), .B2(new_n1120), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1133), .A2(new_n1120), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1219), .B1(new_n1220), .B2(new_n1222), .ZN(G381));
  OR2_X1    g1023(.A1(G393), .A2(G396), .ZN(new_n1224));
  OR4_X1    g1024(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT121), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(G378), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1117), .A2(new_n1135), .A3(KEYINPUT121), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  OR4_X1    g1029(.A1(G387), .A2(new_n1225), .A3(G375), .A4(new_n1229), .ZN(G407));
  NAND2_X1  g1030(.A1(new_n654), .A2(G213), .ZN(new_n1231));
  OR3_X1    g1031(.A1(G375), .A2(new_n1229), .A3(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(G407), .A2(G213), .A3(new_n1232), .ZN(G409));
  INV_X1    g1033(.A(KEYINPUT61), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(G393), .A2(G396), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1224), .A2(new_n1235), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1073), .A2(KEYINPUT110), .A3(new_n1075), .A4(new_n1236), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n1224), .A2(new_n1235), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1069), .A2(new_n1071), .A3(new_n1074), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1074), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1238), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1237), .A2(new_n1241), .A3(new_n1007), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1007), .B1(new_n1237), .B2(new_n1241), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1234), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT122), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n836), .A2(new_n1245), .A3(new_n859), .ZN(new_n1246));
  OAI21_X1  g1046(.A(KEYINPUT60), .B1(new_n1133), .B2(new_n1120), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1247), .A2(new_n1221), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1133), .A2(new_n1120), .A3(KEYINPUT60), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n693), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1219), .B(new_n1246), .C1(new_n1248), .C2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1250), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1247), .A2(new_n1221), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1218), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(G384), .B(new_n1245), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1251), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1231), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1256), .A2(G2897), .A3(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT124), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(G2897), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1251), .B(new_n1260), .C1(new_n1254), .C2(new_n1255), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1258), .A2(new_n1259), .A3(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1259), .B1(new_n1258), .B2(new_n1261), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n693), .B(new_n1162), .C1(new_n1157), .C2(KEYINPUT120), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G378), .B(new_n1199), .C1(new_n1265), .C2(new_n1160), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1197), .B1(new_n1155), .B2(new_n982), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1155), .A2(new_n1156), .A3(new_n1005), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1227), .A2(new_n1228), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1266), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1231), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1244), .B1(new_n1264), .B2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1257), .B1(new_n1266), .B2(new_n1270), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1256), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(KEYINPUT63), .A3(new_n1275), .ZN(new_n1276));
  AOI211_X1 g1076(.A(KEYINPUT123), .B(KEYINPUT63), .C1(new_n1274), .C2(new_n1275), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT123), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1271), .A2(new_n1231), .A3(new_n1275), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT63), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1278), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1273), .B(new_n1276), .C1(new_n1277), .C2(new_n1281), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1234), .B1(new_n1274), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1279), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1274), .A2(KEYINPUT62), .A3(new_n1275), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1285), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1283), .B1(new_n1289), .B2(KEYINPUT125), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1284), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT61), .B1(new_n1272), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1288), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT62), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1294));
  OAI211_X1 g1094(.A(KEYINPUT125), .B(new_n1292), .C1(new_n1293), .C2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1282), .B1(new_n1290), .B2(new_n1296), .ZN(G405));
  INV_X1    g1097(.A(KEYINPUT126), .ZN(new_n1298));
  INV_X1    g1098(.A(G375), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1298), .B(new_n1266), .C1(new_n1299), .C2(new_n1229), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1229), .B1(new_n1163), .B2(new_n1199), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1266), .ZN(new_n1302));
  OAI21_X1  g1102(.A(KEYINPUT126), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1300), .A2(new_n1303), .A3(new_n1275), .ZN(new_n1304));
  OAI211_X1 g1104(.A(KEYINPUT126), .B(new_n1256), .C1(new_n1301), .C2(new_n1302), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1304), .A2(KEYINPUT127), .A3(new_n1283), .A4(new_n1305), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1283), .B(KEYINPUT127), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1306), .B1(new_n1307), .B2(new_n1308), .ZN(G402));
endmodule


