//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G58), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n206), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT64), .B(G77), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G107), .A2(G264), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n203), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n215), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT66), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n234), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT67), .ZN(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XOR2_X1   g0044(.A(G50), .B(G58), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  INV_X1    g0047(.A(KEYINPUT18), .ZN(new_n248));
  AND2_X1   g0048(.A1(G1), .A2(G13), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G226), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G1698), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n254), .B1(G223), .B2(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  INV_X1    g0059(.A(G87), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n252), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT72), .B(G179), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OR2_X1    g0064(.A1(KEYINPUT69), .A2(G1), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT69), .A2(G1), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G41), .A2(G45), .ZN(new_n268));
  OAI211_X1 g0068(.A(G232), .B(new_n251), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT68), .B(G45), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n270), .B(G274), .C1(new_n271), .C2(G41), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n262), .A2(new_n264), .A3(new_n269), .A4(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G223), .A2(G1698), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n274), .B1(new_n253), .B2(G1698), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n259), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n261), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n269), .B(new_n272), .C1(new_n280), .C2(new_n251), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G169), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT16), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n277), .A2(new_n208), .A3(new_n278), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT7), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n277), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n278), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n211), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G58), .A2(G68), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT77), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT77), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G58), .A3(G68), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(new_n292), .A3(new_n212), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G20), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G20), .A2(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G159), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n283), .B1(new_n288), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n255), .A2(new_n256), .ZN(new_n299));
  AOI21_X1  g0099(.A(KEYINPUT7), .B1(new_n299), .B2(new_n208), .ZN(new_n300));
  INV_X1    g0100(.A(new_n287), .ZN(new_n301));
  OAI21_X1  g0101(.A(G68), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n293), .A2(G20), .B1(G159), .B2(new_n295), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n302), .A2(KEYINPUT16), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n207), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n298), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  AND2_X1   g0107(.A1(KEYINPUT69), .A2(G1), .ZN(new_n308));
  NOR2_X1   g0108(.A1(KEYINPUT69), .A2(G1), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n308), .A2(new_n309), .A3(new_n208), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(new_n306), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(KEYINPUT71), .A2(G58), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT8), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n314), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n265), .A2(G13), .A3(G20), .A4(new_n266), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  AOI221_X4 g0119(.A(new_n248), .B1(new_n273), .B2(new_n282), .C1(new_n307), .C2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n307), .A2(new_n319), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n273), .A2(new_n282), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT18), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT78), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n307), .A2(new_n319), .B1(new_n273), .B2(new_n282), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT78), .B1(new_n326), .B2(KEYINPUT18), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n320), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G190), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n281), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n281), .A2(G200), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n307), .A2(new_n330), .A3(new_n319), .A4(new_n331), .ZN(new_n332));
  XOR2_X1   g0132(.A(new_n332), .B(KEYINPUT17), .Z(new_n333));
  OR2_X1    g0133(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n259), .A2(G20), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n314), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G50), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(new_n210), .A3(new_n211), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n338), .A2(G20), .B1(G150), .B2(new_n295), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n306), .ZN(new_n341));
  INV_X1    g0141(.A(new_n317), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n337), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n311), .A2(G50), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n345), .A2(KEYINPUT9), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(KEYINPUT9), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n346), .A2(new_n347), .B1(KEYINPUT74), .B2(KEYINPUT10), .ZN(new_n348));
  INV_X1    g0148(.A(new_n272), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n308), .A2(new_n309), .ZN(new_n350));
  INV_X1    g0150(.A(new_n268), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n252), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n349), .B1(G226), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G1698), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(new_n277), .B2(new_n278), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(G223), .B1(new_n299), .B2(new_n216), .ZN(new_n356));
  AOI21_X1  g0156(.A(G1698), .B1(new_n277), .B2(new_n278), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G222), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n252), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n353), .A2(new_n360), .A3(KEYINPUT70), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT70), .B1(new_n353), .B2(new_n360), .ZN(new_n363));
  OAI21_X1  g0163(.A(G190), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n363), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n365), .A2(G200), .A3(new_n361), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n348), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(KEYINPUT74), .A2(KEYINPUT10), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n368), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n348), .A2(new_n364), .A3(new_n370), .A4(new_n366), .ZN(new_n371));
  INV_X1    g0171(.A(G169), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n365), .A2(new_n372), .A3(new_n361), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n263), .B1(new_n362), .B2(new_n363), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n374), .A3(new_n345), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n369), .A2(new_n371), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G77), .ZN(new_n377));
  OAI22_X1  g0177(.A1(new_n312), .A2(new_n377), .B1(new_n216), .B2(new_n317), .ZN(new_n378));
  INV_X1    g0178(.A(new_n306), .ZN(new_n379));
  XOR2_X1   g0179(.A(KEYINPUT15), .B(G87), .Z(new_n380));
  AOI22_X1  g0180(.A1(new_n380), .A2(new_n335), .B1(new_n216), .B2(G20), .ZN(new_n381));
  XNOR2_X1  g0181(.A(KEYINPUT8), .B(G58), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n295), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n379), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n378), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n352), .A2(G244), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n272), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n357), .A2(G232), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT73), .ZN(new_n391));
  XNOR2_X1  g0191(.A(new_n390), .B(new_n391), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n355), .A2(G238), .B1(new_n299), .B2(G107), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n389), .B1(new_n394), .B2(new_n251), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n386), .B1(new_n395), .B2(new_n329), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n251), .B1(new_n392), .B2(new_n393), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n397), .A2(new_n388), .ZN(new_n398));
  INV_X1    g0198(.A(G200), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OR2_X1    g0200(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT12), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n342), .A2(new_n402), .A3(new_n211), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT12), .B1(new_n317), .B2(G68), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n403), .A2(new_n404), .B1(new_n311), .B2(G68), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT75), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n208), .A2(new_n259), .A3(G50), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n208), .A2(G33), .A3(G77), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n211), .A2(G20), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n410), .A2(KEYINPUT11), .A3(new_n306), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT11), .B1(new_n410), .B2(new_n306), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n406), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n410), .A2(new_n306), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT11), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n410), .A2(KEYINPUT11), .A3(new_n306), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(KEYINPUT75), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n405), .A2(new_n413), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT76), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n405), .A2(new_n413), .A3(new_n418), .A4(KEYINPUT76), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT14), .ZN(new_n424));
  OAI211_X1 g0224(.A(G226), .B(new_n354), .C1(new_n255), .C2(new_n256), .ZN(new_n425));
  OAI211_X1 g0225(.A(G232), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G97), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n428), .A2(new_n252), .ZN(new_n429));
  OAI211_X1 g0229(.A(G238), .B(new_n251), .C1(new_n267), .C2(new_n268), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n272), .ZN(new_n431));
  NOR3_X1   g0231(.A1(new_n429), .A2(KEYINPUT13), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT13), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n430), .A2(new_n272), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n428), .A2(new_n252), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n424), .B(G169), .C1(new_n432), .C2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT13), .B1(new_n429), .B2(new_n431), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n434), .A2(new_n433), .A3(new_n435), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(G179), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n439), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n424), .B1(new_n442), .B2(G169), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n423), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n421), .A2(new_n422), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n442), .A2(G200), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n445), .B(new_n446), .C1(new_n329), .C2(new_n442), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n263), .B(new_n389), .C1(new_n394), .C2(new_n251), .ZN(new_n448));
  INV_X1    g0248(.A(new_n386), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n372), .B1(new_n397), .B2(new_n388), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n401), .A2(new_n444), .A3(new_n447), .A4(new_n451), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n334), .A2(new_n376), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT88), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT25), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(G107), .B1(new_n454), .B2(new_n455), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n456), .B1(new_n342), .B2(new_n457), .ZN(new_n458));
  NOR4_X1   g0258(.A1(new_n317), .A2(new_n454), .A3(new_n455), .A4(G107), .ZN(new_n459));
  INV_X1    g0259(.A(G107), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n265), .A2(G33), .A3(new_n266), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n317), .A2(new_n379), .A3(new_n461), .ZN(new_n462));
  OAI22_X1  g0262(.A1(new_n458), .A2(new_n459), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT87), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(new_n208), .B2(G107), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT23), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT23), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n464), .B(new_n467), .C1(new_n208), .C2(G107), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n466), .A2(new_n468), .B1(G116), .B2(new_n335), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n208), .B(G87), .C1(new_n255), .C2(new_n256), .ZN(new_n470));
  AND2_X1   g0270(.A1(KEYINPUT86), .A2(KEYINPUT22), .ZN(new_n471));
  NOR2_X1   g0271(.A1(KEYINPUT86), .A2(KEYINPUT22), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(G20), .B1(new_n277), .B2(new_n278), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(G87), .A3(new_n471), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n469), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT24), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT24), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n469), .A2(new_n476), .A3(new_n479), .A4(new_n474), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n463), .B1(new_n481), .B2(new_n306), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n265), .A2(G45), .A3(new_n266), .ZN(new_n483));
  AND2_X1   g0283(.A1(KEYINPUT5), .A2(G41), .ZN(new_n484));
  NOR2_X1   g0284(.A1(KEYINPUT5), .A2(G41), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(G264), .B(new_n251), .C1(new_n483), .C2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(G257), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT89), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT89), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n279), .A2(new_n491), .A3(G257), .A4(G1698), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n279), .A2(G250), .A3(new_n354), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G294), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n490), .A2(new_n492), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n488), .B1(new_n495), .B2(new_n252), .ZN(new_n496));
  INV_X1    g0296(.A(G274), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n497), .B1(new_n249), .B2(new_n250), .ZN(new_n498));
  XNOR2_X1  g0298(.A(KEYINPUT5), .B(G41), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n498), .A2(new_n350), .A3(new_n499), .A4(G45), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT81), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G45), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n308), .A2(new_n309), .A3(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n504), .A2(KEYINPUT81), .A3(new_n498), .A4(new_n499), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n496), .A2(new_n329), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(G200), .B1(new_n496), .B2(new_n506), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n482), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(G97), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n342), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n510), .B2(new_n462), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n208), .A2(new_n259), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT79), .B1(new_n513), .B2(new_n377), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT79), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n295), .A2(new_n515), .A3(G77), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT6), .ZN(new_n518));
  AND2_X1   g0318(.A1(G97), .A2(G107), .ZN(new_n519));
  NOR2_X1   g0319(.A1(G97), .A2(G107), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n460), .A2(KEYINPUT6), .A3(G97), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n517), .B(KEYINPUT80), .C1(new_n523), .C2(new_n208), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT80), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n208), .B1(new_n521), .B2(new_n522), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n514), .A2(new_n516), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n460), .B1(new_n286), .B2(new_n287), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n524), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n512), .B1(new_n531), .B2(new_n306), .ZN(new_n532));
  AND2_X1   g0332(.A1(KEYINPUT4), .A2(G244), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n354), .B(new_n533), .C1(new_n255), .C2(new_n256), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G283), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n218), .B1(new_n277), .B2(new_n278), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n534), .B(new_n535), .C1(new_n536), .C2(KEYINPUT4), .ZN(new_n537));
  OAI21_X1  g0337(.A(G250), .B1(new_n255), .B2(new_n256), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n354), .B1(new_n538), .B2(KEYINPUT4), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n252), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n252), .B1(new_n504), .B2(new_n499), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G257), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n506), .A3(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n543), .A2(G190), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n502), .A2(new_n505), .B1(new_n541), .B2(G257), .ZN(new_n545));
  AOI21_X1  g0345(.A(G200), .B1(new_n545), .B2(new_n540), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n532), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n543), .A2(new_n372), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n545), .A2(new_n263), .A3(new_n540), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n526), .A2(new_n527), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n529), .B1(new_n550), .B2(KEYINPUT80), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n379), .B1(new_n551), .B2(new_n528), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n548), .B(new_n549), .C1(new_n552), .C2(new_n512), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n509), .A2(new_n547), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(G116), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n305), .A2(new_n207), .B1(G20), .B2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n535), .B(new_n208), .C1(G33), .C2(new_n510), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT20), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n556), .A2(KEYINPUT20), .A3(new_n557), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n560), .A2(new_n561), .B1(new_n555), .B2(new_n342), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n317), .A2(new_n379), .A3(new_n461), .A4(G116), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n563), .A2(KEYINPUT85), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n563), .A2(KEYINPUT85), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(G257), .B(new_n354), .C1(new_n255), .C2(new_n256), .ZN(new_n567));
  OAI211_X1 g0367(.A(G264), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n568));
  INV_X1    g0368(.A(G303), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n567), .B(new_n568), .C1(new_n569), .C2(new_n279), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n252), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n541), .A2(G270), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n506), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n566), .A2(new_n573), .A3(G169), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT21), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n573), .A2(G200), .ZN(new_n577));
  INV_X1    g0377(.A(new_n561), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT20), .B1(new_n556), .B2(new_n557), .ZN(new_n579));
  OAI22_X1  g0379(.A1(new_n578), .A2(new_n579), .B1(G116), .B2(new_n317), .ZN(new_n580));
  INV_X1    g0380(.A(new_n565), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n563), .A2(KEYINPUT85), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n506), .A2(G190), .A3(new_n571), .A4(new_n572), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n577), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n506), .A2(G179), .A3(new_n571), .A4(new_n572), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n566), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n566), .A2(new_n573), .A3(KEYINPUT21), .A4(G169), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n576), .A2(new_n585), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n208), .B(G68), .C1(new_n255), .C2(new_n256), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT19), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n260), .A2(new_n510), .A3(new_n460), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n427), .A2(new_n208), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR4_X1   g0395(.A1(new_n259), .A2(new_n510), .A3(KEYINPUT19), .A4(G20), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n591), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT83), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(KEYINPUT83), .B(new_n591), .C1(new_n595), .C2(new_n596), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n306), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n380), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n342), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT84), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n462), .B2(new_n602), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n306), .B1(new_n350), .B2(G33), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n606), .A2(KEYINPUT84), .A3(new_n317), .A4(new_n380), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n601), .A2(new_n603), .A3(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(G244), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n610));
  OAI211_X1 g0410(.A(G238), .B(new_n354), .C1(new_n255), .C2(new_n256), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n610), .B(new_n611), .C1(new_n259), .C2(new_n555), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n252), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n504), .A2(new_n498), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n483), .A2(G250), .A3(new_n251), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n613), .A2(new_n616), .A3(new_n263), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT82), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n609), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n613), .A2(new_n616), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n372), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n618), .B1(new_n622), .B2(new_n617), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n606), .A2(G87), .A3(new_n317), .ZN(new_n624));
  NOR3_X1   g0424(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n625));
  AOI21_X1  g0425(.A(G20), .B1(G33), .B2(G97), .ZN(new_n626));
  OAI21_X1  g0426(.A(KEYINPUT19), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n335), .A2(new_n592), .A3(G97), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n627), .A2(new_n628), .B1(new_n475), .B2(G68), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n306), .B1(new_n629), .B2(KEYINPUT83), .ZN(new_n630));
  INV_X1    g0430(.A(new_n600), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n624), .B(new_n603), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n621), .A2(G200), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n613), .A2(new_n616), .A3(G190), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI22_X1  g0435(.A1(new_n620), .A2(new_n623), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(G179), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n496), .A2(new_n637), .A3(new_n506), .ZN(new_n638));
  AOI21_X1  g0438(.A(G169), .B1(new_n496), .B2(new_n506), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n482), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NOR4_X1   g0440(.A1(new_n554), .A2(new_n590), .A3(new_n636), .A4(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n453), .A2(new_n641), .ZN(G372));
  INV_X1    g0442(.A(new_n375), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n369), .A2(new_n371), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT93), .B1(new_n320), .B2(new_n323), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n315), .A2(new_n318), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n288), .A2(new_n297), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n379), .B1(new_n647), .B2(KEYINPUT16), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n646), .B1(new_n648), .B2(new_n298), .ZN(new_n649));
  INV_X1    g0449(.A(new_n322), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n248), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT93), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n321), .A2(KEYINPUT18), .A3(new_n322), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n645), .A2(new_n654), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n441), .A2(new_n443), .ZN(new_n656));
  INV_X1    g0456(.A(new_n451), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n656), .A2(new_n423), .B1(new_n657), .B2(new_n447), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n655), .B1(new_n658), .B2(new_n333), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n644), .B1(new_n659), .B2(KEYINPUT94), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT94), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n661), .B(new_n655), .C1(new_n658), .C2(new_n333), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n643), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n453), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n632), .A2(KEYINPUT90), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT90), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n601), .A2(new_n666), .A3(new_n624), .A4(new_n603), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n635), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n609), .A2(new_n617), .A3(new_n622), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n668), .A2(new_n553), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT92), .B1(new_n670), .B2(KEYINPUT26), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n665), .A2(new_n667), .ZN(new_n672));
  INV_X1    g0472(.A(new_n635), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n553), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n609), .A2(new_n617), .A3(new_n622), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT92), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT26), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n636), .A2(new_n553), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(KEYINPUT26), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n671), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n676), .B(KEYINPUT91), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n554), .A2(new_n668), .A3(new_n669), .ZN(new_n685));
  INV_X1    g0485(.A(new_n639), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n496), .A2(new_n637), .A3(new_n506), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n379), .B1(new_n478), .B2(new_n480), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n686), .B(new_n687), .C1(new_n688), .C2(new_n463), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n574), .A2(new_n575), .B1(new_n587), .B2(new_n566), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(new_n690), .A3(new_n589), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n684), .B1(new_n685), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n683), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n663), .B1(new_n664), .B2(new_n694), .ZN(G369));
  NAND2_X1  g0495(.A1(new_n690), .A2(new_n589), .ZN(new_n696));
  INV_X1    g0496(.A(G213), .ZN(new_n697));
  INV_X1    g0497(.A(G13), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G20), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n350), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT95), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT95), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n700), .A2(new_n704), .A3(KEYINPUT27), .ZN(new_n705));
  AOI211_X1 g0505(.A(new_n697), .B(new_n701), .C1(new_n703), .C2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G343), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(new_n583), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n696), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n590), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n703), .A2(new_n705), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n701), .A2(new_n697), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n713), .A2(G343), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n688), .B2(new_n463), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n640), .B1(new_n509), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n689), .A2(new_n715), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n712), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n696), .A2(new_n707), .ZN(new_n721));
  OAI22_X1  g0521(.A1(new_n717), .A2(new_n721), .B1(new_n689), .B2(new_n715), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n720), .A2(new_n723), .ZN(G399));
  INV_X1    g0524(.A(new_n204), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G41), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n593), .A2(G116), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(G1), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n213), .B2(new_n727), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT28), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT29), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n509), .A2(new_n553), .A3(new_n547), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n668), .A2(new_n669), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(new_n691), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n677), .A2(KEYINPUT26), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n681), .A2(new_n679), .ZN(new_n737));
  INV_X1    g0537(.A(new_n684), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n735), .A2(new_n736), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n732), .B1(new_n739), .B2(new_n707), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n715), .B1(new_n683), .B2(new_n692), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n740), .B1(new_n732), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n614), .A2(new_n615), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n743), .B1(new_n252), .B2(new_n612), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n496), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(KEYINPUT96), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n586), .A2(new_n543), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT96), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n496), .A2(new_n744), .A3(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n746), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT30), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n746), .A2(new_n747), .A3(KEYINPUT30), .A4(new_n749), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n496), .A2(new_n506), .ZN(new_n754));
  AND3_X1   g0554(.A1(new_n754), .A2(new_n263), .A3(new_n543), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT97), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n744), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n621), .A2(KEYINPUT97), .ZN(new_n758));
  AND3_X1   g0558(.A1(new_n757), .A2(new_n758), .A3(new_n573), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n752), .A2(new_n753), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n715), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT31), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n750), .A2(new_n751), .B1(new_n755), .B2(new_n759), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n707), .B1(new_n765), .B2(new_n753), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(KEYINPUT31), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n636), .A2(new_n640), .ZN(new_n768));
  INV_X1    g0568(.A(new_n590), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n768), .A2(new_n733), .A3(new_n769), .A4(new_n707), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n764), .A2(new_n767), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G330), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n742), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n731), .B1(new_n773), .B2(G1), .ZN(G364));
  AOI21_X1  g0574(.A(new_n270), .B1(new_n699), .B2(G45), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n726), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n712), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(G330), .B2(new_n710), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n777), .B(KEYINPUT98), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n279), .A2(new_n204), .ZN(new_n781));
  INV_X1    g0581(.A(G355), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n781), .A2(new_n782), .B1(G116), .B2(new_n204), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n246), .A2(G45), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n725), .A2(new_n279), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  XOR2_X1   g0586(.A(KEYINPUT68), .B(G45), .Z(new_n787));
  AOI21_X1  g0587(.A(new_n786), .B1(new_n214), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n783), .B1(new_n784), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n207), .B1(G20), .B2(new_n372), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n780), .B1(new_n789), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n263), .A2(new_n208), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n329), .A2(G200), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G322), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n399), .A2(G190), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(KEYINPUT33), .B(G317), .Z(new_n804));
  OAI22_X1  g0604(.A1(new_n800), .A2(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G190), .A2(G200), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n797), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n805), .B1(G311), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n329), .A2(new_n399), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n208), .A2(G179), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n299), .B1(new_n812), .B2(new_n569), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n811), .A2(new_n802), .ZN(new_n814));
  INV_X1    g0614(.A(G283), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n811), .A2(new_n806), .ZN(new_n816));
  INV_X1    g0616(.A(G329), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n814), .A2(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n798), .A2(new_n637), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(G20), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n813), .B(new_n818), .C1(G294), .C2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G326), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n797), .A2(new_n810), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT101), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n809), .B(new_n821), .C1(new_n822), .C2(new_n824), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n825), .A2(KEYINPUT102), .ZN(new_n826));
  INV_X1    g0626(.A(new_n820), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n510), .ZN(new_n828));
  INV_X1    g0628(.A(new_n803), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n828), .B1(G68), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT100), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n279), .B1(new_n814), .B2(new_n460), .C1(new_n260), .C2(new_n812), .ZN(new_n832));
  INV_X1    g0632(.A(new_n823), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(G50), .B2(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n216), .A2(new_n808), .B1(new_n799), .B2(G58), .ZN(new_n835));
  INV_X1    g0635(.A(new_n816), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(G159), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT99), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT32), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n831), .A2(new_n834), .A3(new_n835), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n825), .A2(KEYINPUT102), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n826), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n796), .B1(new_n842), .B2(new_n793), .ZN(new_n843));
  INV_X1    g0643(.A(new_n792), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n710), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n779), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(G396));
  INV_X1    g0647(.A(KEYINPUT105), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n707), .B2(new_n386), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n449), .A2(KEYINPUT105), .A3(new_n715), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n401), .A2(new_n451), .A3(new_n707), .A4(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(new_n683), .B2(new_n692), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n451), .A2(new_n715), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n849), .B(new_n850), .C1(new_n396), .C2(new_n400), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n855), .B1(new_n856), .B2(new_n451), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n854), .B1(new_n741), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n777), .B1(new_n858), .B2(new_n772), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n772), .B2(new_n858), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n555), .A2(new_n807), .B1(new_n803), .B2(new_n815), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT103), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n861), .A2(new_n862), .B1(new_n569), .B2(new_n823), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n862), .B2(new_n861), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT104), .ZN(new_n865));
  INV_X1    g0665(.A(G294), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n800), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n814), .A2(new_n260), .ZN(new_n868));
  INV_X1    g0668(.A(new_n812), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n868), .B1(G107), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(G311), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n870), .B(new_n299), .C1(new_n871), .C2(new_n816), .ZN(new_n872));
  NOR4_X1   g0672(.A1(new_n865), .A2(new_n828), .A3(new_n867), .A4(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(G132), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n279), .B1(new_n816), .B2(new_n874), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n812), .A2(new_n337), .B1(new_n814), .B2(new_n211), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n875), .B(new_n876), .C1(G58), .C2(new_n820), .ZN(new_n877));
  AOI22_X1  g0677(.A1(G137), .A2(new_n833), .B1(new_n799), .B2(G143), .ZN(new_n878));
  INV_X1    g0678(.A(G150), .ZN(new_n879));
  INV_X1    g0679(.A(G159), .ZN(new_n880));
  OAI221_X1 g0680(.A(new_n878), .B1(new_n879), .B2(new_n803), .C1(new_n880), .C2(new_n807), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT34), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n877), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n882), .B2(new_n881), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n793), .B1(new_n873), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n780), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n793), .A2(new_n790), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n886), .B1(new_n377), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n885), .B(new_n888), .C1(new_n791), .C2(new_n857), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n860), .A2(new_n889), .ZN(G384));
  INV_X1    g0690(.A(new_n523), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n891), .A2(KEYINPUT35), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(KEYINPUT35), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n892), .A2(G116), .A3(new_n209), .A4(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT36), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n217), .A2(new_n293), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n896), .A2(new_n337), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n267), .B(new_n698), .C1(G50), .C2(G68), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n321), .A2(new_n706), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n332), .B(KEYINPUT17), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n900), .B1(new_n655), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n322), .A2(new_n706), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n332), .B1(new_n903), .B2(new_n649), .ZN(new_n904));
  INV_X1    g0704(.A(new_n903), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT108), .B1(new_n905), .B2(new_n321), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n905), .A2(new_n321), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n909), .A2(KEYINPUT108), .A3(KEYINPUT37), .A4(new_n332), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n899), .B1(new_n902), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n647), .A2(KEYINPUT107), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT107), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n288), .B2(new_n297), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n913), .A2(new_n283), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n646), .B1(new_n916), .B2(new_n648), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n713), .A2(new_n714), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n328), .B2(new_n333), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n332), .B1(new_n917), .B2(new_n903), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT37), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(KEYINPUT37), .B2(new_n904), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n920), .A2(KEYINPUT38), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n912), .A2(new_n924), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n421), .A2(new_n715), .A3(new_n422), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n444), .A2(new_n447), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n926), .B1(new_n441), .B2(new_n443), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT106), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT106), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n926), .B(new_n931), .C1(new_n441), .C2(new_n443), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n928), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n857), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n641), .A2(new_n707), .B1(new_n762), .B2(new_n763), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n934), .B1(new_n935), .B2(new_n767), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n925), .A2(new_n936), .A3(KEYINPUT40), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT109), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT40), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n912), .B2(new_n924), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(KEYINPUT109), .A3(new_n936), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n920), .A2(new_n923), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n899), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n924), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n936), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n940), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n943), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n453), .A2(new_n771), .ZN(new_n951));
  OAI21_X1  g0751(.A(G330), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n951), .B2(new_n950), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT39), .B1(new_n912), .B2(new_n924), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n656), .A2(new_n423), .A3(new_n707), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n945), .A2(KEYINPUT39), .A3(new_n924), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n955), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n855), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n854), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n961), .A2(new_n946), .A3(new_n933), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n645), .A2(new_n654), .A3(new_n918), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n959), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n663), .B1(new_n742), .B2(new_n664), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n964), .B(new_n965), .Z(new_n966));
  NAND2_X1  g0766(.A1(new_n953), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n953), .A2(new_n966), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT110), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n967), .B1(new_n350), .B2(new_n699), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n968), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(KEYINPUT110), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n895), .B1(new_n897), .B2(new_n898), .C1(new_n970), .C2(new_n972), .ZN(G367));
  NOR2_X1   g0773(.A1(new_n234), .A2(new_n786), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n794), .B1(new_n204), .B2(new_n602), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n780), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI22_X1  g0776(.A1(G283), .A2(new_n808), .B1(new_n829), .B2(G294), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n869), .A2(G116), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT46), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n977), .B(new_n979), .C1(new_n569), .C2(new_n800), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n824), .A2(new_n871), .ZN(new_n981));
  INV_X1    g0781(.A(new_n814), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n279), .B1(new_n982), .B2(G97), .ZN(new_n983));
  INV_X1    g0783(.A(G317), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n983), .B1(new_n984), .B2(new_n816), .C1(new_n460), .C2(new_n827), .ZN(new_n985));
  NOR3_X1   g0785(.A1(new_n980), .A2(new_n981), .A3(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT114), .Z(new_n987));
  INV_X1    g0787(.A(G143), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n824), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n820), .A2(G68), .ZN(new_n990));
  INV_X1    g0790(.A(G137), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n990), .B1(new_n210), .B2(new_n812), .C1(new_n991), .C2(new_n816), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G150), .B2(new_n799), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n279), .B1(new_n217), .B2(new_n814), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT115), .ZN(new_n995));
  AOI22_X1  g0795(.A1(G50), .A2(new_n808), .B1(new_n829), .B2(G159), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n987), .B1(new_n989), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT47), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n976), .B1(new_n999), .B2(new_n793), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n665), .A2(new_n667), .A3(new_n715), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n734), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n738), .B2(new_n1001), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1000), .B1(new_n844), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n721), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n675), .A2(new_n715), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n547), .B(new_n553), .C1(new_n532), .C2(new_n707), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n719), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(KEYINPUT42), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT42), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n719), .A2(new_n1011), .A3(new_n1005), .A4(new_n1008), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n553), .B1(new_n1007), .B2(new_n689), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n707), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1010), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT112), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1015), .A2(new_n1016), .B1(KEYINPUT43), .B2(new_n1003), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n1016), .B2(new_n1015), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1003), .A2(KEYINPUT43), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT111), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(KEYINPUT113), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1008), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n720), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1018), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1024), .B1(new_n1018), .B2(new_n1022), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n1026), .A2(new_n1027), .B1(KEYINPUT113), .B2(new_n1021), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1027), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1021), .A2(KEYINPUT113), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1029), .A2(new_n1030), .A3(new_n1025), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n723), .A2(new_n1008), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT45), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1033), .B(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n722), .A2(new_n1023), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT44), .Z(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1038), .A2(new_n712), .A3(new_n719), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1035), .A2(new_n1037), .A3(new_n720), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n719), .B(new_n721), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(new_n711), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n773), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n773), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n726), .B(KEYINPUT41), .Z(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n776), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1004), .B1(new_n1032), .B2(new_n1048), .ZN(G387));
  NAND2_X1  g0849(.A1(new_n1043), .A2(new_n776), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n382), .A2(G50), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT50), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n503), .B1(new_n211), .B2(new_n377), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n728), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1053), .B1(new_n1054), .B2(KEYINPUT116), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1052), .B(new_n1055), .C1(KEYINPUT116), .C2(new_n1054), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1056), .B(new_n785), .C1(new_n238), .C2(new_n787), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(G107), .B2(new_n204), .C1(new_n728), .C2(new_n781), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n886), .B1(new_n1058), .B2(new_n794), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n800), .A2(new_n337), .B1(new_n211), .B2(new_n807), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n299), .B1(new_n982), .B2(G97), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n820), .A2(new_n380), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n869), .A2(new_n216), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n836), .A2(G150), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n880), .A2(new_n823), .B1(new_n803), .B2(new_n316), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n1060), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G303), .A2(new_n808), .B1(new_n829), .B2(G311), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n984), .B2(new_n800), .C1(new_n824), .C2(new_n801), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT48), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n827), .A2(new_n815), .B1(new_n812), .B2(new_n866), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1074), .A2(KEYINPUT49), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n299), .B1(new_n816), .B2(new_n822), .C1(new_n555), .C2(new_n814), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n1074), .B2(KEYINPUT49), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1067), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n793), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1059), .B1(new_n719), .B2(new_n844), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1044), .A2(new_n726), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n773), .A2(new_n1043), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1050), .B(new_n1080), .C1(new_n1081), .C2(new_n1082), .ZN(G393));
  NAND2_X1  g0883(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT118), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1041), .A2(new_n1044), .A3(KEYINPUT118), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1089), .A2(new_n727), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1023), .A2(new_n792), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n243), .A2(new_n786), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n794), .B1(new_n510), .B2(new_n204), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n780), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n800), .A2(new_n871), .B1(new_n984), .B2(new_n823), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT52), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n299), .B1(new_n814), .B2(new_n460), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n812), .A2(new_n815), .B1(new_n816), .B2(new_n801), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1098), .B(new_n1099), .C1(G116), .C2(new_n820), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G294), .A2(new_n808), .B1(new_n829), .B2(G303), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1097), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G150), .A2(new_n833), .B1(new_n799), .B2(G159), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(KEYINPUT117), .B(KEYINPUT51), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n827), .A2(new_n377), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n812), .A2(new_n211), .B1(new_n816), .B2(new_n988), .ZN(new_n1108));
  NOR4_X1   g0908(.A1(new_n1107), .A2(new_n299), .A3(new_n868), .A4(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(G50), .A2(new_n829), .B1(new_n808), .B2(new_n383), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1106), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1102), .B1(new_n1105), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1095), .B1(new_n1112), .B2(new_n793), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1092), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n1041), .B2(new_n775), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1091), .A2(new_n1116), .ZN(G390));
  OAI21_X1  g0917(.A(new_n770), .B1(KEYINPUT31), .B2(new_n766), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n762), .A2(new_n763), .ZN(new_n1119));
  OAI211_X1 g0919(.A(G330), .B(new_n857), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n933), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n771), .A2(G330), .A3(new_n857), .A4(new_n933), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n961), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n739), .A2(new_n707), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n855), .B1(new_n1126), .B2(new_n857), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1127), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n453), .A2(G330), .A3(new_n771), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n663), .B(new_n1130), .C1(new_n742), .C2(new_n664), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1123), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n925), .A2(new_n956), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n739), .A2(new_n707), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n857), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n960), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1135), .B1(new_n933), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n933), .B1(new_n853), .B2(new_n855), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n956), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1141), .A2(KEYINPUT119), .B1(new_n955), .B2(new_n958), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT119), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1140), .A2(new_n1143), .A3(new_n956), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1134), .B(new_n1139), .C1(new_n1142), .C2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1141), .A2(KEYINPUT119), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n955), .A2(new_n958), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1146), .A2(new_n1147), .A3(new_n1144), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1139), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1123), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1133), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1144), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1143), .B1(new_n1140), .B2(new_n956), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n924), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT38), .B1(new_n920), .B2(new_n923), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n954), .B1(KEYINPUT39), .B2(new_n1156), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n1152), .A2(new_n1153), .A3(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1134), .B1(new_n1158), .B2(new_n1139), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1148), .A2(new_n1123), .A3(new_n1149), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1133), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1151), .A2(new_n1162), .A3(new_n726), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n887), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(G97), .A2(new_n808), .B1(new_n799), .B2(G116), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n460), .B2(new_n803), .C1(new_n815), .C2(new_n823), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n299), .B1(new_n812), .B2(new_n260), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n814), .A2(new_n211), .B1(new_n816), .B2(new_n866), .ZN(new_n1168));
  NOR4_X1   g0968(.A1(new_n1166), .A2(new_n1107), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G128), .A2(new_n833), .B1(new_n799), .B2(G132), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n1170), .B(KEYINPUT120), .Z(new_n1171));
  OAI21_X1  g0971(.A(new_n279), .B1(new_n814), .B2(new_n337), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G125), .B2(new_n836), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT54), .B(G143), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1173), .B1(new_n991), .B2(new_n803), .C1(new_n807), .C2(new_n1174), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n812), .A2(KEYINPUT53), .A3(new_n879), .ZN(new_n1176));
  OAI21_X1  g0976(.A(KEYINPUT53), .B1(new_n812), .B2(new_n879), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n827), .B2(new_n880), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1175), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1169), .B1(new_n1171), .B2(new_n1179), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n780), .B1(new_n314), .B2(new_n1164), .C1(new_n1180), .C2(new_n1079), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n1147), .B2(new_n790), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1145), .A2(new_n1150), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1182), .B1(new_n1183), .B2(new_n776), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1163), .A2(new_n1184), .ZN(G378));
  AOI211_X1 g0985(.A(new_n776), .B(new_n726), .C1(new_n337), .C2(new_n887), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n827), .A2(new_n879), .B1(new_n812), .B2(new_n1174), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G132), .A2(new_n829), .B1(new_n799), .B2(G128), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n991), .B2(new_n807), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1187), .B(new_n1189), .C1(G125), .C2(new_n833), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n982), .A2(G159), .ZN(new_n1193));
  AOI211_X1 g0993(.A(G33), .B(G41), .C1(new_n836), .C2(G124), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT59), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1195), .B1(new_n1196), .B2(new_n1190), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n279), .A2(G41), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n337), .B1(G33), .B2(G41), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n990), .B1(new_n823), .B2(new_n555), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT121), .Z(new_n1202));
  AOI22_X1  g1002(.A1(G58), .A2(new_n982), .B1(new_n836), .B2(G283), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1203), .A2(new_n1063), .A3(new_n1198), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G97), .B2(new_n829), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n380), .A2(new_n808), .B1(new_n799), .B2(G107), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1202), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT58), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1200), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1209), .B(KEYINPUT122), .Z(new_n1210));
  NOR2_X1   g1010(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n1197), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  XOR2_X1   g1012(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1213));
  XNOR2_X1  g1013(.A(new_n376), .B(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n706), .A2(new_n345), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT123), .Z(new_n1216));
  XOR2_X1   g1016(.A(new_n1214), .B(new_n1216), .Z(new_n1217));
  OAI221_X1 g1017(.A(new_n1186), .B1(new_n1079), .B2(new_n1212), .C1(new_n1217), .C2(new_n791), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  AND4_X1   g1019(.A1(KEYINPUT109), .A2(new_n925), .A3(new_n936), .A4(KEYINPUT40), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT109), .B1(new_n941), .B2(new_n936), .ZN(new_n1221));
  OAI211_X1 g1021(.A(G330), .B(new_n948), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1217), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n943), .A2(G330), .A3(new_n948), .A4(new_n1217), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n964), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n964), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1224), .A2(new_n1225), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1219), .B1(new_n1230), .B2(new_n776), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1131), .B1(new_n1183), .B2(new_n1129), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1224), .A2(new_n1228), .A3(new_n1225), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1228), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1234));
  OAI21_X1  g1034(.A(KEYINPUT57), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n726), .B1(new_n1232), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1162), .A2(new_n1132), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT57), .B1(new_n1237), .B2(new_n1230), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1231), .B1(new_n1236), .B2(new_n1238), .ZN(G375));
  NAND2_X1  g1039(.A1(new_n1121), .A2(new_n790), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n780), .B1(G68), .B2(new_n1164), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(G97), .A2(new_n869), .B1(new_n836), .B2(G303), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n279), .B1(new_n982), .B2(G77), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1242), .A2(new_n1062), .A3(new_n1243), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(G107), .A2(new_n808), .B1(new_n799), .B2(G283), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n1245), .B1(new_n555), .B2(new_n803), .C1(new_n866), .C2(new_n823), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(G150), .A2(new_n808), .B1(new_n799), .B2(G137), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n1247), .B1(new_n874), .B2(new_n823), .C1(new_n803), .C2(new_n1174), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(G159), .A2(new_n869), .B1(new_n836), .B2(G128), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n299), .B1(new_n982), .B2(G58), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1249), .B(new_n1250), .C1(new_n337), .C2(new_n827), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n1244), .A2(new_n1246), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1241), .B1(new_n1252), .B2(new_n793), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1129), .A2(new_n776), .B1(new_n1240), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1133), .A2(new_n1047), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1254), .B1(new_n1255), .B2(new_n1256), .ZN(G381));
  INV_X1    g1057(.A(G375), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n1163), .A2(new_n1184), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1031), .B(new_n1028), .C1(new_n1260), .C2(new_n776), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1115), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(new_n1004), .A3(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NOR4_X1   g1064(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1258), .A2(new_n1259), .A3(new_n1264), .A4(new_n1265), .ZN(G407));
  NOR2_X1   g1066(.A1(new_n697), .A2(G343), .ZN(new_n1267));
  XOR2_X1   g1067(.A(new_n1267), .B(KEYINPUT124), .Z(new_n1268));
  NAND3_X1  g1068(.A1(new_n1258), .A2(new_n1259), .A3(new_n1268), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1269), .B(KEYINPUT125), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1270), .A2(G213), .A3(G407), .ZN(G409));
  OAI211_X1 g1071(.A(G378), .B(new_n1231), .C1(new_n1236), .C2(new_n1238), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1237), .A2(new_n1230), .A3(new_n1047), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1218), .B1(new_n1274), .B2(new_n775), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1259), .B1(new_n1273), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1272), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1267), .ZN(new_n1278));
  INV_X1    g1078(.A(G384), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1131), .A2(new_n1125), .A3(KEYINPUT60), .A4(new_n1128), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n726), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1256), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1127), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n1122), .A2(new_n1123), .B1(new_n960), .B2(new_n854), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(KEYINPUT60), .B1(new_n1285), .B2(new_n1131), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1281), .B1(new_n1282), .B2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1254), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1279), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1256), .B1(new_n1133), .B2(KEYINPUT60), .ZN(new_n1290));
  OAI211_X1 g1090(.A(G384), .B(new_n1254), .C1(new_n1290), .C2(new_n1281), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1277), .A2(new_n1278), .A3(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT63), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1267), .A2(G2897), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1289), .A2(new_n1291), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(KEYINPUT126), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT126), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1289), .A2(new_n1291), .A3(new_n1300), .A4(new_n1297), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1292), .A2(G2897), .A3(new_n1268), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(G390), .A2(G387), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(G393), .B(new_n846), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1263), .A2(new_n1308), .A3(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1310), .B1(new_n1263), .B2(new_n1308), .ZN(new_n1312));
  NOR3_X1   g1112(.A1(new_n1311), .A2(new_n1312), .A3(KEYINPUT61), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1268), .B1(new_n1272), .B2(new_n1276), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1314), .A2(KEYINPUT63), .A3(new_n1293), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1296), .A2(new_n1307), .A3(new_n1313), .A4(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT61), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1317), .B1(new_n1314), .B2(new_n1304), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT62), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1294), .A2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1314), .A2(KEYINPUT62), .A3(new_n1293), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1318), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1316), .B1(new_n1322), .B2(new_n1323), .ZN(G405));
  NOR2_X1   g1124(.A1(new_n1293), .A2(KEYINPUT127), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1325), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1263), .A2(new_n1308), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1309), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1263), .A2(new_n1308), .A3(new_n1310), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1325), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1328), .A2(new_n1329), .A3(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1326), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT127), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1272), .B1(new_n1333), .B2(new_n1292), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1334), .B1(new_n1259), .B2(G375), .ZN(new_n1335));
  XNOR2_X1  g1135(.A(new_n1332), .B(new_n1335), .ZN(G402));
endmodule


