//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n812, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n986, new_n987,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1049, new_n1050,
    new_n1051;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G1gat), .B2(new_n202), .ZN(new_n206));
  OR2_X1    g005(.A1(new_n206), .A2(G8gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(G8gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT21), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT9), .ZN(new_n212));
  NOR3_X1   g011(.A1(new_n212), .A2(G71gat), .A3(G78gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(G71gat), .A2(G78gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G64gat), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n216), .A2(G57gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(G57gat), .ZN(new_n218));
  OAI22_X1  g017(.A1(new_n213), .A2(new_n215), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G57gat), .B(G64gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n214), .B1(new_n220), .B2(new_n212), .ZN(new_n221));
  NOR2_X1   g020(.A1(G71gat), .A2(G78gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT93), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n222), .B(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n219), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n210), .B1(new_n211), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(G183gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(G231gat), .A2(G233gat), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT94), .B(KEYINPUT20), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n222), .B(KEYINPUT93), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT9), .B1(new_n217), .B2(new_n218), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(new_n233), .A3(new_n214), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT21), .B1(new_n234), .B2(new_n219), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(KEYINPUT96), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(G211gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(G127gat), .B(G155gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n231), .B(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  XOR2_X1   g042(.A(G190gat), .B(G218gat), .Z(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(KEYINPUT98), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G29gat), .A2(G36gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT90), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT14), .ZN(new_n251));
  INV_X1    g050(.A(G29gat), .ZN(new_n252));
  INV_X1    g051(.A(G36gat), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT89), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  OR2_X1    g056(.A1(new_n256), .A2(new_n255), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n250), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G43gat), .B(G50gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(KEYINPUT15), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT91), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT15), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT15), .ZN(new_n264));
  INV_X1    g063(.A(G50gat), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n265), .A2(G43gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(G43gat), .ZN(new_n267));
  OAI211_X1 g066(.A(KEYINPUT91), .B(new_n264), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n254), .A2(new_n256), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n263), .A2(new_n268), .A3(new_n250), .A4(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n261), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G99gat), .A2(G106gat), .ZN(new_n272));
  INV_X1    g071(.A(G85gat), .ZN(new_n273));
  INV_X1    g072(.A(G92gat), .ZN(new_n274));
  AOI22_X1  g073(.A1(KEYINPUT8), .A2(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G99gat), .B(G106gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(G85gat), .A2(G92gat), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT7), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n275), .A2(new_n276), .A3(new_n279), .A4(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n272), .A2(KEYINPUT8), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n273), .A2(new_n274), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n282), .A2(new_n279), .A3(new_n283), .A4(new_n280), .ZN(new_n284));
  INV_X1    g083(.A(new_n276), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n271), .A2(new_n281), .A3(new_n286), .ZN(new_n287));
  AND2_X1   g086(.A1(G232gat), .A2(G233gat), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n245), .A2(KEYINPUT98), .B1(KEYINPUT41), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT97), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n271), .A2(KEYINPUT17), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT17), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n261), .A2(new_n292), .A3(new_n270), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n286), .A2(new_n281), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n290), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n261), .A2(new_n292), .A3(new_n270), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n292), .B1(new_n261), .B2(new_n270), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n290), .B(new_n295), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n287), .B(new_n289), .C1(new_n296), .C2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n288), .A2(KEYINPUT41), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n295), .B1(new_n297), .B2(new_n298), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT97), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(new_n299), .ZN(new_n306));
  INV_X1    g105(.A(new_n302), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n306), .A2(new_n307), .A3(new_n287), .A4(new_n289), .ZN(new_n308));
  XOR2_X1   g107(.A(G134gat), .B(G162gat), .Z(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n303), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n310), .B1(new_n303), .B2(new_n308), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n247), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n303), .A2(new_n308), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(new_n309), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n303), .A2(new_n308), .A3(new_n310), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n315), .A2(new_n246), .A3(new_n316), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n243), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT38), .ZN(new_n320));
  XNOR2_X1  g119(.A(G8gat), .B(G36gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(G64gat), .B(G92gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT77), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT69), .ZN(new_n325));
  INV_X1    g124(.A(G183gat), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n325), .B1(new_n326), .B2(KEYINPUT27), .ZN(new_n327));
  AOI21_X1  g126(.A(G190gat), .B1(new_n326), .B2(KEYINPUT27), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT27), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n329), .A2(KEYINPUT69), .A3(G183gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n327), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT70), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT28), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n327), .A2(new_n328), .A3(KEYINPUT70), .A4(new_n330), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n329), .A2(G183gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n328), .A2(KEYINPUT28), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT71), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n340), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n341), .A2(new_n343), .A3(KEYINPUT71), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT26), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT65), .ZN(new_n349));
  NOR3_X1   g148(.A1(new_n349), .A2(G169gat), .A3(G176gat), .ZN(new_n350));
  INV_X1    g149(.A(G169gat), .ZN(new_n351));
  INV_X1    g150(.A(G176gat), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT65), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n348), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  AOI22_X1  g153(.A1(new_n347), .A2(new_n354), .B1(G183gat), .B2(G190gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT72), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT72), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n339), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT68), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT23), .B1(new_n351), .B2(new_n352), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n344), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n343), .A2(KEYINPUT23), .ZN(new_n363));
  NAND2_X1  g162(.A1(G183gat), .A2(G190gat), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT24), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(G183gat), .A2(G190gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n368), .B2(KEYINPUT64), .ZN(new_n369));
  NAND3_X1  g168(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT64), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n370), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n362), .B(new_n363), .C1(new_n369), .C2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT25), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT23), .B1(new_n350), .B2(new_n353), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n374), .B1(new_n361), .B2(new_n344), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT66), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n370), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g177(.A1(KEYINPUT66), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n378), .A2(new_n368), .A3(new_n366), .A4(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n375), .A2(new_n376), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT67), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n375), .A2(new_n376), .A3(new_n380), .A4(KEYINPUT67), .ZN(new_n384));
  AOI221_X4 g183(.A(new_n360), .B1(new_n373), .B2(new_n374), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n384), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n373), .A2(new_n374), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT68), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n357), .B(new_n359), .C1(new_n385), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G226gat), .A2(G233gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n391), .A2(KEYINPUT29), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  XOR2_X1   g192(.A(G197gat), .B(G204gat), .Z(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT76), .B(G211gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(G218gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT22), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G211gat), .B(G218gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n399), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT22), .B1(new_n395), .B2(G218gat), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n401), .B1(new_n402), .B2(new_n394), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT23), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n406), .B1(G169gat), .B2(G176gat), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT25), .B1(new_n407), .B2(new_n343), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT65), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n349), .B1(G169gat), .B2(G176gat), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n406), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT67), .B1(new_n412), .B2(new_n380), .ZN(new_n413));
  INV_X1    g212(.A(new_n384), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n387), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(new_n356), .A3(new_n391), .ZN(new_n416));
  AND4_X1   g215(.A1(new_n324), .A2(new_n393), .A3(new_n405), .A4(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n393), .A2(new_n405), .A3(new_n416), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n415), .A2(new_n360), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n386), .A2(KEYINPUT68), .A3(new_n387), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n339), .A2(new_n355), .A3(new_n358), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n358), .B1(new_n339), .B2(new_n355), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n421), .A2(new_n424), .A3(new_n391), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n415), .A2(new_n356), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n392), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n405), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(new_n324), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n417), .B1(new_n418), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n323), .B1(new_n430), .B2(KEYINPUT37), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n425), .A2(new_n427), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n405), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n393), .A2(new_n404), .A3(new_n416), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n433), .A2(KEYINPUT37), .A3(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n320), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n432), .A2(new_n404), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n437), .A2(KEYINPUT77), .A3(new_n418), .ZN(new_n438));
  INV_X1    g237(.A(new_n416), .ZN(new_n439));
  AOI211_X1 g238(.A(new_n404), .B(new_n439), .C1(new_n389), .C2(new_n392), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n324), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT37), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT38), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n436), .B1(new_n431), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G141gat), .B(G148gat), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n446), .A2(KEYINPUT2), .ZN(new_n447));
  XNOR2_X1  g246(.A(G155gat), .B(G162gat), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT79), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(G141gat), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n452), .A2(G148gat), .ZN(new_n453));
  INV_X1    g252(.A(G148gat), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n454), .A2(G141gat), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT79), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(G155gat), .A2(G162gat), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n451), .A2(new_n456), .B1(KEYINPUT2), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n448), .B(KEYINPUT80), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n449), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT4), .ZN(new_n461));
  XNOR2_X1  g260(.A(G113gat), .B(G120gat), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n462), .A2(KEYINPUT1), .ZN(new_n463));
  XNOR2_X1  g262(.A(G127gat), .B(G134gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n464), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n466), .B1(KEYINPUT1), .B2(new_n462), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n460), .A2(new_n461), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n461), .B1(new_n460), .B2(new_n469), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT81), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OR2_X1    g272(.A1(new_n447), .A2(new_n448), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n457), .A2(KEYINPUT2), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n446), .A2(new_n450), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n454), .A2(G141gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n452), .A2(G148gat), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n477), .A2(new_n478), .A3(new_n450), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n475), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT80), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n448), .B(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n474), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n483), .A2(new_n468), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(KEYINPUT81), .A3(new_n461), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n473), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(G225gat), .A2(G233gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n483), .A2(KEYINPUT3), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT3), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n460), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n490), .A3(new_n468), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n486), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n487), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n460), .A2(new_n469), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n493), .B1(new_n484), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT5), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(G1gat), .B(G29gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(new_n273), .ZN(new_n500));
  XNOR2_X1  g299(.A(KEYINPUT0), .B(G57gat), .ZN(new_n501));
  XOR2_X1   g300(.A(new_n500), .B(new_n501), .Z(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n484), .B(new_n461), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n493), .A2(KEYINPUT5), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n491), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n498), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n493), .B1(new_n473), .B2(new_n485), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n496), .B1(new_n508), .B2(new_n491), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n504), .A2(new_n491), .A3(new_n505), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n502), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT6), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n507), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n506), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n514), .A2(KEYINPUT82), .A3(KEYINPUT6), .A4(new_n502), .ZN(new_n515));
  OAI211_X1 g314(.A(KEYINPUT6), .B(new_n502), .C1(new_n509), .C2(new_n510), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT82), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n513), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n323), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n519), .B1(new_n442), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n445), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(G228gat), .ZN(new_n523));
  INV_X1    g322(.A(G233gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT29), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n490), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n405), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT29), .B1(new_n400), .B2(new_n403), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n483), .B1(new_n530), .B2(KEYINPUT3), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n526), .B1(new_n532), .B2(KEYINPUT84), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT84), .ZN(new_n534));
  AOI211_X1 g333(.A(new_n534), .B(new_n525), .C1(new_n529), .C2(new_n531), .ZN(new_n535));
  OAI21_X1  g334(.A(G22gat), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n532), .A2(KEYINPUT84), .A3(new_n526), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n404), .A2(new_n527), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n460), .B1(new_n538), .B2(new_n489), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n404), .B1(new_n490), .B2(new_n527), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT84), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n525), .ZN(new_n542));
  INV_X1    g341(.A(G22gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n537), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n536), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G78gat), .B(G106gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT83), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT31), .B(G50gat), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n547), .B(new_n548), .Z(new_n549));
  NAND2_X1  g348(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT86), .ZN(new_n551));
  INV_X1    g350(.A(new_n549), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT85), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n537), .A2(new_n542), .A3(new_n553), .A4(new_n543), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n536), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n544), .A2(KEYINPUT85), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n551), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n536), .A2(new_n554), .A3(new_n552), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n544), .A2(KEYINPUT85), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n558), .A2(new_n559), .A3(KEYINPUT86), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n550), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT87), .ZN(new_n562));
  NOR3_X1   g361(.A1(new_n440), .A2(new_n428), .A3(new_n324), .ZN(new_n563));
  OAI211_X1 g362(.A(KEYINPUT30), .B(new_n520), .C1(new_n563), .C2(new_n417), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n438), .A2(new_n441), .A3(new_n323), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT30), .B1(new_n442), .B2(new_n520), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n562), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT30), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(new_n430), .B2(new_n323), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n570), .A2(KEYINPUT87), .A3(new_n565), .A4(new_n564), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n504), .A2(new_n491), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n493), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n484), .A2(new_n494), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n575), .B(KEYINPUT39), .C1(new_n493), .C2(new_n576), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n577), .B(new_n503), .C1(KEYINPUT39), .C2(new_n575), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT40), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n579), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(new_n511), .A3(new_n581), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n522), .B(new_n561), .C1(new_n573), .C2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT78), .ZN(new_n584));
  AOI211_X1 g383(.A(new_n569), .B(new_n323), .C1(new_n438), .C2(new_n441), .ZN(new_n585));
  INV_X1    g384(.A(new_n565), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n564), .A2(KEYINPUT78), .A3(new_n565), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n587), .A2(new_n588), .A3(new_n519), .A4(new_n570), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n555), .A2(new_n551), .A3(new_n556), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT86), .B1(new_n558), .B2(new_n559), .ZN(new_n591));
  AOI22_X1  g390(.A1(new_n590), .A2(new_n591), .B1(new_n545), .B2(new_n549), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n385), .A2(new_n388), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n357), .A2(new_n359), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT73), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT73), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n421), .A2(new_n424), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n596), .A2(new_n468), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(G227gat), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n600), .A2(new_n524), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n389), .A2(KEYINPUT73), .A3(new_n469), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT32), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT33), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G15gat), .B(G43gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT74), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(G71gat), .ZN(new_n609));
  INV_X1    g408(.A(G99gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n604), .A2(new_n606), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n611), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n603), .B(KEYINPUT32), .C1(new_n605), .C2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT75), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT34), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n599), .A2(new_n602), .ZN(new_n618));
  INV_X1    g417(.A(new_n601), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI211_X1 g419(.A(KEYINPUT34), .B(new_n601), .C1(new_n599), .C2(new_n602), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n615), .A2(new_n616), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n618), .A2(new_n619), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT34), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n618), .A2(new_n617), .A3(new_n619), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n625), .A2(new_n616), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(KEYINPUT75), .B1(new_n620), .B2(new_n621), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n627), .A2(new_n628), .A3(new_n614), .A4(new_n612), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT36), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n623), .A2(new_n629), .A3(KEYINPUT36), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n583), .A2(new_n593), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT35), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n519), .A2(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n568), .A2(new_n571), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT88), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n630), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n623), .A2(new_n629), .A3(KEYINPUT88), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n638), .A2(new_n640), .A3(new_n561), .A4(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n630), .A2(new_n561), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT35), .B1(new_n643), .B2(new_n589), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n319), .B1(new_n635), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G229gat), .A2(G233gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT13), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n209), .A2(new_n271), .ZN(new_n650));
  AOI22_X1  g449(.A1(new_n207), .A2(new_n208), .B1(new_n270), .B2(new_n261), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT92), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g453(.A(KEYINPUT92), .B(new_n649), .C1(new_n650), .C2(new_n651), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n294), .A2(new_n210), .ZN(new_n657));
  INV_X1    g456(.A(new_n651), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(new_n647), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT18), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n657), .A2(KEYINPUT18), .A3(new_n647), .A4(new_n658), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n656), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G113gat), .B(G141gat), .ZN(new_n664));
  INV_X1    g463(.A(G197gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT11), .B(G169gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT12), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n656), .A2(new_n661), .A3(new_n662), .A4(new_n669), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n225), .A2(new_n295), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n234), .A2(new_n281), .A3(new_n286), .A4(new_n219), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(G230gat), .A2(G233gat), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT101), .B(G120gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(G148gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(G176gat), .B(G204gat), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n682), .B(new_n683), .Z(new_n684));
  INV_X1    g483(.A(KEYINPUT10), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n675), .A2(new_n676), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT99), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n676), .A2(new_n685), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n675), .A2(new_n676), .A3(KEYINPUT99), .A4(new_n685), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n691), .A2(KEYINPUT100), .A3(new_n678), .ZN(new_n692));
  AOI21_X1  g491(.A(KEYINPUT100), .B1(new_n691), .B2(new_n678), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n680), .B(new_n684), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n691), .A2(new_n678), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n680), .ZN(new_n696));
  INV_X1    g495(.A(new_n684), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n674), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n646), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n519), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g503(.A1(new_n701), .A2(new_n572), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT16), .B(G8gat), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT42), .Z(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(G8gat), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(G1325gat));
  INV_X1    g509(.A(new_n641), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT88), .B1(new_n623), .B2(new_n629), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(G15gat), .B1(new_n701), .B2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n634), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n701), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n714), .B1(new_n716), .B2(G15gat), .ZN(G1326gat));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n592), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT43), .B(G22gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1327gat));
  AOI21_X1  g519(.A(new_n318), .B1(new_n635), .B2(new_n645), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n242), .A2(new_n700), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n724), .A2(new_n252), .A3(new_n702), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT45), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n721), .A2(KEYINPUT44), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n568), .A2(new_n561), .A3(new_n571), .A4(new_n637), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n711), .A2(new_n728), .A3(new_n712), .ZN(new_n729));
  INV_X1    g528(.A(new_n589), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n592), .B1(new_n623), .B2(new_n629), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n636), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(KEYINPUT102), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT102), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n642), .A2(new_n644), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n318), .B1(new_n736), .B2(new_n635), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n723), .B(new_n727), .C1(new_n737), .C2(KEYINPUT44), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT103), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n593), .A2(new_n632), .A3(new_n633), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n582), .B1(new_n568), .B2(new_n571), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n592), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n741), .B1(new_n522), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n744), .B1(new_n733), .B2(new_n735), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n740), .B1(new_n745), .B2(new_n318), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT103), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n746), .A2(new_n747), .A3(new_n723), .A4(new_n727), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n519), .B1(new_n739), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n726), .B1(new_n749), .B2(new_n252), .ZN(G1328gat));
  NAND3_X1  g549(.A1(new_n724), .A2(new_n253), .A3(new_n572), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT46), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n573), .B1(new_n739), .B2(new_n748), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n753), .B1(new_n754), .B2(new_n253), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT104), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n753), .B(KEYINPUT104), .C1(new_n754), .C2(new_n253), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(G1329gat));
  INV_X1    g558(.A(new_n724), .ZN(new_n760));
  INV_X1    g559(.A(new_n713), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n760), .A2(G43gat), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(G43gat), .B1(new_n738), .B2(new_n634), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n763), .A2(KEYINPUT47), .A3(new_n764), .ZN(new_n765));
  AOI211_X1 g564(.A(new_n740), .B(new_n318), .C1(new_n635), .C2(new_n645), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n729), .A2(new_n732), .A3(KEYINPUT102), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n734), .B1(new_n642), .B2(new_n644), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n635), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n313), .A2(new_n317), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n766), .B1(new_n771), .B2(new_n740), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n747), .B1(new_n772), .B2(new_n723), .ZN(new_n773));
  INV_X1    g572(.A(new_n748), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n715), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n762), .B1(new_n775), .B2(G43gat), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n765), .B1(new_n776), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g576(.A1(new_n760), .A2(G50gat), .A3(new_n561), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(G50gat), .B1(new_n738), .B2(new_n561), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n779), .A2(KEYINPUT48), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n592), .B1(new_n773), .B2(new_n774), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n778), .B1(new_n782), .B2(G50gat), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n783), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g583(.A1(new_n745), .A2(new_n673), .ZN(new_n785));
  INV_X1    g584(.A(new_n699), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n319), .A2(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n519), .B(KEYINPUT105), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(G57gat), .ZN(G1332gat));
  INV_X1    g590(.A(KEYINPUT49), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n572), .B1(new_n792), .B2(new_n216), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT106), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n788), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n792), .A2(new_n216), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n795), .B(new_n796), .ZN(G1333gat));
  XOR2_X1   g596(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n785), .A2(new_n713), .A3(new_n787), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT107), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n785), .A2(KEYINPUT107), .A3(new_n713), .A4(new_n787), .ZN(new_n803));
  AOI21_X1  g602(.A(G71gat), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(G71gat), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n788), .B2(new_n715), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n799), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n804), .A2(new_n798), .A3(new_n807), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(G1334gat));
  NAND2_X1  g610(.A1(new_n788), .A2(new_n592), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g612(.A1(new_n243), .A2(new_n673), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n769), .A2(new_n770), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n737), .A2(KEYINPUT51), .A3(new_n814), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT109), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n817), .A2(new_n818), .A3(KEYINPUT109), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n821), .A2(new_n273), .A3(new_n699), .A4(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n814), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(new_n786), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n772), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n826), .A2(new_n702), .ZN(new_n827));
  OAI22_X1  g626(.A1(new_n823), .A2(new_n519), .B1(new_n827), .B2(new_n273), .ZN(G1336gat));
  NAND3_X1  g627(.A1(new_n772), .A2(new_n572), .A3(new_n825), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(G92gat), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n819), .A2(new_n274), .A3(new_n699), .A4(new_n572), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT52), .ZN(G1337gat));
  NAND4_X1  g632(.A1(new_n821), .A2(new_n610), .A3(new_n699), .A4(new_n822), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n826), .A2(new_n715), .ZN(new_n835));
  OAI22_X1  g634(.A1(new_n834), .A2(new_n761), .B1(new_n835), .B2(new_n610), .ZN(G1338gat));
  NOR2_X1   g635(.A1(new_n561), .A2(G106gat), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT51), .B1(new_n737), .B2(new_n814), .ZN(new_n838));
  NOR4_X1   g637(.A1(new_n745), .A2(new_n816), .A3(new_n318), .A4(new_n824), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n699), .B(new_n837), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT111), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n819), .A2(KEYINPUT111), .A3(new_n699), .A4(new_n837), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n746), .A2(new_n592), .A3(new_n727), .A4(new_n825), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(G106gat), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n842), .A2(new_n843), .A3(new_n844), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n840), .A2(new_n846), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT110), .B1(new_n848), .B2(KEYINPUT53), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT110), .ZN(new_n850));
  AOI211_X1 g649(.A(new_n850), .B(new_n843), .C1(new_n840), .C2(new_n846), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n847), .B1(new_n849), .B2(new_n851), .ZN(G1339gat));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n688), .A2(new_n679), .A3(new_n689), .A4(new_n690), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n854), .A2(KEYINPUT54), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n855), .B1(new_n692), .B2(new_n693), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n691), .A2(new_n857), .A3(new_n678), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n858), .A2(new_n697), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n856), .A2(KEYINPUT55), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n694), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n860), .A2(KEYINPUT112), .A3(new_n694), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n856), .A2(new_n859), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT55), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n863), .A2(new_n673), .A3(new_n864), .A4(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n672), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n647), .B1(new_n657), .B2(new_n658), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n870), .A2(KEYINPUT113), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n650), .A2(new_n651), .A3(new_n649), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT114), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n870), .A2(KEYINPUT113), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n869), .B1(new_n668), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n699), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n770), .B1(new_n868), .B2(new_n877), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n863), .A2(new_n876), .A3(new_n864), .A4(new_n867), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(new_n318), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n853), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n860), .A2(KEYINPUT112), .A3(new_n694), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT112), .B1(new_n860), .B2(new_n694), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n884), .A2(new_n770), .A3(new_n876), .A4(new_n867), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n673), .A2(new_n867), .ZN(new_n886));
  AOI22_X1  g685(.A1(new_n884), .A2(new_n886), .B1(new_n699), .B2(new_n876), .ZN(new_n887));
  OAI211_X1 g686(.A(KEYINPUT115), .B(new_n885), .C1(new_n887), .C2(new_n770), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n881), .A2(new_n888), .A3(new_n242), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n243), .A2(new_n674), .A3(new_n786), .A4(new_n318), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n889), .A2(KEYINPUT116), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT116), .B1(new_n889), .B2(new_n890), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(KEYINPUT117), .A3(new_n561), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n889), .A2(new_n890), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT116), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n889), .A2(KEYINPUT116), .A3(new_n890), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n897), .A2(new_n561), .A3(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT117), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n894), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n572), .A2(new_n519), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n713), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G113gat), .B1(new_n904), .B2(new_n674), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n893), .A2(new_n573), .A3(new_n789), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(new_n643), .ZN(new_n907));
  INV_X1    g706(.A(G113gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n907), .A2(new_n908), .A3(new_n673), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n905), .A2(new_n909), .ZN(G1340gat));
  OAI21_X1  g709(.A(G120gat), .B1(new_n904), .B2(new_n786), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n786), .A2(G120gat), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT118), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n907), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n911), .A2(new_n914), .ZN(G1341gat));
  INV_X1    g714(.A(G127gat), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n904), .A2(new_n916), .A3(new_n242), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n906), .A2(new_n643), .A3(new_n242), .ZN(new_n918));
  XOR2_X1   g717(.A(new_n918), .B(KEYINPUT119), .Z(new_n919));
  AOI21_X1  g718(.A(new_n917), .B1(new_n919), .B2(new_n916), .ZN(G1342gat));
  NOR4_X1   g719(.A1(new_n906), .A2(G134gat), .A3(new_n643), .A4(new_n318), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT56), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(G134gat), .B1(new_n904), .B2(new_n318), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n921), .A2(new_n922), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(G1343gat));
  NAND2_X1  g725(.A1(new_n897), .A2(new_n898), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n927), .A2(KEYINPUT57), .A3(new_n561), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n634), .A2(new_n903), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n865), .A2(KEYINPUT120), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT55), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n865), .A2(KEYINPUT120), .A3(new_n866), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n931), .A2(new_n673), .A3(new_n694), .A4(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n933), .A2(new_n934), .A3(new_n877), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n934), .B1(new_n933), .B2(new_n877), .ZN(new_n937));
  OAI211_X1 g736(.A(KEYINPUT122), .B(new_n318), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(new_n885), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n933), .A2(new_n877), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT121), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n935), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT122), .B1(new_n942), .B2(new_n318), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n242), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n561), .B1(new_n944), .B2(new_n890), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT57), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n929), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(KEYINPUT123), .B1(new_n928), .B2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(new_n890), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n942), .A2(new_n318), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT122), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n952), .A2(new_n885), .A3(new_n938), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n949), .B1(new_n953), .B2(new_n242), .ZN(new_n954));
  OAI21_X1  g753(.A(KEYINPUT57), .B1(new_n954), .B2(new_n561), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n893), .A2(new_n946), .A3(new_n592), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT123), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n955), .A2(new_n956), .A3(new_n957), .A4(new_n929), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n948), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n452), .B1(new_n959), .B2(new_n673), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n715), .A2(new_n561), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n906), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n963), .A2(new_n452), .A3(new_n673), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(KEYINPUT58), .B1(new_n960), .B2(new_n965), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n955), .A2(new_n956), .A3(new_n673), .A4(new_n929), .ZN(new_n967));
  AOI21_X1  g766(.A(KEYINPUT58), .B1(new_n967), .B2(G141gat), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(new_n964), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(KEYINPUT124), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT124), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n968), .A2(new_n971), .A3(new_n964), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n966), .A2(new_n970), .A3(new_n972), .ZN(G1344gat));
  OAI21_X1  g772(.A(KEYINPUT57), .B1(new_n927), .B2(new_n561), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n243), .B1(new_n950), .B2(new_n885), .ZN(new_n975));
  OAI211_X1 g774(.A(new_n946), .B(new_n592), .C1(new_n975), .C2(new_n949), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n977), .A2(KEYINPUT59), .A3(new_n699), .A4(new_n929), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n786), .B1(new_n948), .B2(new_n958), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n978), .B1(new_n979), .B2(KEYINPUT59), .ZN(new_n980));
  AOI21_X1  g779(.A(G148gat), .B1(new_n963), .B2(new_n699), .ZN(new_n981));
  AOI22_X1  g780(.A1(new_n980), .A2(G148gat), .B1(KEYINPUT59), .B2(new_n981), .ZN(G1345gat));
  AOI21_X1  g781(.A(G155gat), .B1(new_n963), .B2(new_n243), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n242), .B1(new_n948), .B2(new_n958), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n983), .B1(new_n984), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g784(.A(G162gat), .B1(new_n963), .B2(new_n770), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n318), .B1(new_n948), .B2(new_n958), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n986), .B1(new_n987), .B2(G162gat), .ZN(G1347gat));
  NAND3_X1  g787(.A1(new_n893), .A2(new_n519), .A3(new_n572), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n989), .A2(new_n643), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n990), .A2(new_n351), .A3(new_n673), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n573), .A2(new_n789), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n713), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n993), .B1(new_n894), .B2(new_n901), .ZN(new_n994));
  AND2_X1   g793(.A1(new_n994), .A2(new_n673), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n991), .B1(new_n995), .B2(new_n351), .ZN(G1348gat));
  AOI21_X1  g795(.A(G176gat), .B1(new_n990), .B2(new_n699), .ZN(new_n997));
  AND2_X1   g796(.A1(new_n994), .A2(new_n699), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n997), .B1(new_n998), .B2(G176gat), .ZN(G1349gat));
  INV_X1    g798(.A(new_n993), .ZN(new_n1000));
  AOI21_X1  g799(.A(KEYINPUT117), .B1(new_n893), .B2(new_n561), .ZN(new_n1001));
  NOR4_X1   g800(.A1(new_n891), .A2(new_n892), .A3(new_n900), .A4(new_n592), .ZN(new_n1002));
  OAI211_X1 g801(.A(new_n243), .B(new_n1000), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(KEYINPUT125), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT125), .ZN(new_n1005));
  NAND4_X1  g804(.A1(new_n902), .A2(new_n1005), .A3(new_n243), .A4(new_n1000), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n1004), .A2(G183gat), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n326), .A2(KEYINPUT27), .ZN(new_n1008));
  NAND4_X1  g807(.A1(new_n990), .A2(new_n1008), .A3(new_n337), .A4(new_n243), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1010), .A2(KEYINPUT60), .ZN(new_n1011));
  INV_X1    g810(.A(KEYINPUT60), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n1007), .A2(new_n1012), .A3(new_n1009), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1011), .A2(new_n1013), .ZN(G1350gat));
  AOI211_X1 g813(.A(new_n318), .B(new_n993), .C1(new_n894), .C2(new_n901), .ZN(new_n1015));
  INV_X1    g814(.A(G190gat), .ZN(new_n1016));
  OAI21_X1  g815(.A(KEYINPUT126), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n994), .A2(new_n770), .ZN(new_n1018));
  INV_X1    g817(.A(KEYINPUT126), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n1018), .A2(new_n1019), .A3(G190gat), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g820(.A(KEYINPUT61), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g822(.A1(new_n990), .A2(new_n1016), .A3(new_n770), .ZN(new_n1024));
  NAND3_X1  g823(.A1(new_n1017), .A2(new_n1020), .A3(KEYINPUT61), .ZN(new_n1025));
  NAND3_X1  g824(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(G1351gat));
  NOR2_X1   g825(.A1(new_n989), .A2(new_n962), .ZN(new_n1027));
  OR2_X1    g826(.A1(new_n1027), .A2(KEYINPUT127), .ZN(new_n1028));
  NAND2_X1  g827(.A1(new_n1027), .A2(KEYINPUT127), .ZN(new_n1029));
  NAND4_X1  g828(.A1(new_n1028), .A2(new_n665), .A3(new_n673), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g829(.A1(new_n634), .A2(new_n992), .ZN(new_n1031));
  INV_X1    g830(.A(new_n1031), .ZN(new_n1032));
  AND2_X1   g831(.A1(new_n977), .A2(new_n1032), .ZN(new_n1033));
  AND2_X1   g832(.A1(new_n1033), .A2(new_n673), .ZN(new_n1034));
  OAI21_X1  g833(.A(new_n1030), .B1(new_n1034), .B2(new_n665), .ZN(G1352gat));
  NAND3_X1  g834(.A1(new_n977), .A2(new_n699), .A3(new_n1032), .ZN(new_n1036));
  NAND2_X1  g835(.A1(new_n1036), .A2(G204gat), .ZN(new_n1037));
  NOR4_X1   g836(.A1(new_n989), .A2(G204gat), .A3(new_n786), .A4(new_n962), .ZN(new_n1038));
  INV_X1    g837(.A(KEYINPUT62), .ZN(new_n1039));
  OR2_X1    g838(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  NAND3_X1  g840(.A1(new_n1037), .A2(new_n1040), .A3(new_n1041), .ZN(G1353gat));
  INV_X1    g841(.A(new_n395), .ZN(new_n1043));
  NAND4_X1  g842(.A1(new_n1028), .A2(new_n1043), .A3(new_n243), .A4(new_n1029), .ZN(new_n1044));
  NAND3_X1  g843(.A1(new_n977), .A2(new_n243), .A3(new_n1032), .ZN(new_n1045));
  AND3_X1   g844(.A1(new_n1045), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1046));
  AOI21_X1  g845(.A(KEYINPUT63), .B1(new_n1045), .B2(G211gat), .ZN(new_n1047));
  OAI21_X1  g846(.A(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(G1354gat));
  NAND3_X1  g847(.A1(new_n1028), .A2(new_n770), .A3(new_n1029), .ZN(new_n1049));
  INV_X1    g848(.A(G218gat), .ZN(new_n1050));
  NOR2_X1   g849(.A1(new_n318), .A2(new_n1050), .ZN(new_n1051));
  AOI22_X1  g850(.A1(new_n1049), .A2(new_n1050), .B1(new_n1033), .B2(new_n1051), .ZN(G1355gat));
endmodule


