//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1253, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n208), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT65), .B(G77), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G58), .A2(G232), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n223), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n210), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n213), .B(new_n218), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT66), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n235), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT67), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NOR2_X1   g0048(.A1(G58), .A2(G68), .ZN(new_n249));
  INV_X1    g0049(.A(G50), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n208), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT71), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT69), .ZN(new_n254));
  XOR2_X1   g0054(.A(KEYINPUT8), .B(G58), .Z(new_n255));
  NAND2_X1  g0055(.A1(new_n208), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n254), .A2(G150), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT70), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n252), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(new_n259), .B2(new_n258), .ZN(new_n261));
  NAND3_X1  g0061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n216), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(G50), .B1(new_n208), .B2(G1), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT72), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(new_n263), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n266), .A2(new_n269), .B1(new_n250), .B2(new_n268), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g0071(.A(new_n271), .B(KEYINPUT9), .Z(new_n272));
  INV_X1    g0072(.A(KEYINPUT74), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT10), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(KEYINPUT3), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G222), .A2(G1698), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G223), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n280), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n284), .B(new_n285), .C1(new_n219), .C2(new_n280), .ZN(new_n286));
  INV_X1    g0086(.A(G274), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n288));
  NOR3_X1   g0088(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n288), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n289), .B1(G226), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n286), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT68), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n293), .B(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G200), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(G190), .B2(new_n295), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n271), .B(KEYINPUT9), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT74), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n274), .A2(new_n275), .A3(new_n298), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n298), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT75), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT75), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n302), .A2(new_n305), .A3(KEYINPUT10), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n301), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n295), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n309), .B(new_n271), .C1(G169), .C2(new_n295), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G87), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n278), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT76), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n276), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT77), .ZN(new_n316));
  NAND2_X1  g0116(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n315), .A2(new_n316), .A3(G33), .A4(new_n317), .ZN(new_n318));
  AND2_X1   g0118(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n319));
  NOR2_X1   g0119(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n319), .A2(new_n320), .A3(new_n278), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT77), .B1(new_n276), .B2(G33), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n318), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(G223), .A2(G1698), .ZN(new_n324));
  INV_X1    g0124(.A(G226), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n324), .B1(new_n325), .B2(G1698), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n313), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT79), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n326), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n315), .A2(G33), .A3(new_n317), .ZN(new_n331));
  INV_X1    g0131(.A(new_n322), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n330), .B1(new_n333), .B2(new_n318), .ZN(new_n334));
  OAI21_X1  g0134(.A(KEYINPUT79), .B1(new_n334), .B2(new_n313), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n329), .A2(new_n285), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n289), .B1(G232), .B2(new_n291), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G169), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n336), .A2(G179), .A3(new_n337), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT16), .ZN(new_n342));
  INV_X1    g0142(.A(G68), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT78), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n344), .B(new_n278), .C1(new_n319), .C2(new_n320), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT7), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n346), .A2(G20), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n319), .A2(new_n320), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n348), .A2(G33), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT78), .B1(new_n278), .B2(KEYINPUT3), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n345), .B(new_n347), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n346), .B1(new_n280), .B2(G20), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n343), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g0153(.A(G58), .B(G68), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n254), .A2(G159), .B1(new_n354), .B2(G20), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n342), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n333), .A2(new_n208), .A3(new_n318), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT7), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(G68), .B1(new_n358), .B2(KEYINPUT7), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n355), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n357), .B(new_n263), .C1(new_n362), .C2(new_n342), .ZN(new_n363));
  INV_X1    g0163(.A(new_n255), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n207), .B2(G20), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n365), .A2(new_n269), .B1(new_n364), .B2(new_n268), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n341), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT18), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n363), .A2(new_n366), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n336), .A2(G190), .A3(new_n337), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n338), .A2(G200), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n370), .A2(KEYINPUT17), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT18), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n341), .A2(new_n367), .A3(new_n374), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n372), .A2(new_n363), .A3(new_n366), .A4(new_n371), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT17), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n369), .A2(new_n373), .A3(new_n375), .A4(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n254), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n380), .A2(new_n250), .ZN(new_n381));
  INV_X1    g0181(.A(G77), .ZN(new_n382));
  OAI22_X1  g0182(.A1(new_n256), .A2(new_n382), .B1(new_n208), .B2(G68), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n263), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT11), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n385), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT12), .B1(new_n267), .B2(G68), .ZN(new_n388));
  OR3_X1    g0188(.A1(new_n267), .A2(KEYINPUT12), .A3(G68), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n343), .B1(new_n207), .B2(G20), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n388), .A2(new_n389), .B1(new_n269), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n386), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n285), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n232), .A2(G1698), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n280), .B(new_n394), .C1(G226), .C2(G1698), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G97), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n393), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n291), .A2(G238), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n397), .A2(new_n289), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT13), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n399), .A2(new_n400), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT14), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n405), .A3(G169), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n402), .A2(G179), .A3(new_n403), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n405), .B1(new_n404), .B2(G169), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n392), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(G190), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n404), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n296), .B1(new_n402), .B2(new_n403), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n412), .A2(new_n413), .A3(new_n392), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n380), .A2(new_n364), .ZN(new_n416));
  XNOR2_X1  g0216(.A(KEYINPUT15), .B(G87), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n220), .A2(new_n208), .B1(new_n417), .B2(new_n256), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n263), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n269), .ZN(new_n420));
  OAI21_X1  g0220(.A(G77), .B1(new_n208), .B2(G1), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n219), .A2(KEYINPUT73), .A3(new_n267), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT73), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(new_n220), .B2(new_n268), .ZN(new_n424));
  OAI221_X1 g0224(.A(new_n419), .B1(new_n420), .B2(new_n421), .C1(new_n422), .C2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(G232), .A2(G1698), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n282), .A2(G238), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n280), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n428), .B(new_n285), .C1(G107), .C2(new_n280), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n289), .B1(G244), .B2(new_n291), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n425), .B1(new_n432), .B2(G190), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n296), .B2(new_n432), .ZN(new_n434));
  INV_X1    g0234(.A(G169), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n425), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n432), .A2(new_n308), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n410), .A2(new_n415), .A3(new_n434), .A4(new_n439), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n311), .A2(new_n379), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G45), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(G1), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT5), .B(G41), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n285), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G257), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n445), .A2(new_n444), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n285), .A2(new_n287), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n282), .A2(G244), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n452), .B1(new_n333), .B2(new_n318), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT80), .B1(new_n453), .B2(KEYINPUT4), .ZN(new_n454));
  INV_X1    g0254(.A(new_n452), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n322), .B1(new_n348), .B2(G33), .ZN(new_n456));
  INV_X1    g0256(.A(new_n318), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT80), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT4), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G250), .ZN(new_n462));
  OAI22_X1  g0262(.A1(new_n452), .A2(new_n460), .B1(new_n462), .B2(new_n282), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n280), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n454), .A2(new_n461), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n451), .B1(new_n468), .B2(new_n285), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n308), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT4), .B1(new_n323), .B2(new_n455), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n466), .B1(new_n471), .B2(new_n459), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n393), .B1(new_n472), .B2(new_n454), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n435), .B1(new_n473), .B2(new_n451), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n267), .A2(G97), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n262), .A2(new_n216), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n476), .B(new_n267), .C1(G1), .C2(new_n278), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n475), .B1(new_n478), .B2(G97), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT6), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n480), .A2(new_n202), .A3(G107), .ZN(new_n481));
  XNOR2_X1  g0281(.A(G97), .B(G107), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n481), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  OAI22_X1  g0283(.A1(new_n380), .A2(new_n382), .B1(new_n483), .B2(new_n208), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n351), .A2(new_n352), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n484), .B1(new_n485), .B2(G107), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n479), .B1(new_n486), .B2(new_n476), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n470), .A2(new_n474), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(G200), .B1(new_n473), .B2(new_n451), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n468), .A2(new_n285), .ZN(new_n490));
  INV_X1    g0290(.A(new_n451), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n490), .A2(G190), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n487), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n489), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT81), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n489), .A2(new_n492), .A3(KEYINPUT81), .A4(new_n493), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n488), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n221), .A2(G1698), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(G238), .B2(G1698), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n500), .B1(new_n333), .B2(new_n318), .ZN(new_n501));
  INV_X1    g0301(.A(G116), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n278), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n285), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n285), .A2(new_n462), .A3(new_n444), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n505), .B1(new_n449), .B2(new_n444), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n435), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(G179), .B2(new_n507), .ZN(new_n509));
  INV_X1    g0309(.A(new_n417), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n478), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n510), .A2(new_n267), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n256), .A2(KEYINPUT19), .A3(new_n202), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n396), .A2(new_n208), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n204), .B2(G87), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n514), .B1(new_n516), .B2(KEYINPUT19), .ZN(new_n517));
  AOI21_X1  g0317(.A(G20), .B1(new_n333), .B2(new_n318), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(G68), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n263), .B1(new_n519), .B2(KEYINPUT82), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n323), .A2(new_n208), .A3(G68), .ZN(new_n521));
  INV_X1    g0321(.A(new_n517), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(KEYINPUT82), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n511), .B(new_n513), .C1(new_n520), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT83), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT82), .ZN(new_n527));
  AOI211_X1 g0327(.A(G20), .B(new_n343), .C1(new_n333), .C2(new_n318), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n527), .B1(new_n528), .B2(new_n517), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(new_n263), .A3(new_n523), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT83), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n530), .A2(new_n531), .A3(new_n511), .A4(new_n513), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n509), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n504), .A2(G190), .A3(new_n506), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT84), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n504), .A2(KEYINPUT84), .A3(G190), .A4(new_n506), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n521), .A2(new_n522), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n476), .B1(new_n539), .B2(new_n527), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n512), .B1(new_n540), .B2(new_n523), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n478), .A2(G87), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n507), .A2(G200), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n538), .A2(new_n541), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n533), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n498), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n462), .A2(new_n282), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(G257), .B2(new_n282), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n333), .B2(new_n318), .ZN(new_n550));
  INV_X1    g0350(.A(G294), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n278), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n285), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n446), .A2(G264), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n450), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT87), .B1(new_n555), .B2(G169), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n553), .A2(G179), .A3(new_n450), .A4(new_n554), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n555), .A2(KEYINPUT87), .A3(G169), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n503), .A2(new_n208), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT23), .B1(new_n203), .B2(G20), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n203), .A2(KEYINPUT23), .A3(G20), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n561), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n312), .A2(G20), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT22), .B1(new_n280), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(KEYINPUT22), .A2(G87), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  AOI211_X1 g0370(.A(KEYINPUT86), .B(new_n568), .C1(new_n518), .C2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT86), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n323), .A2(new_n208), .A3(new_n570), .ZN(new_n573));
  INV_X1    g0373(.A(new_n568), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n566), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT24), .ZN(new_n577));
  AOI211_X1 g0377(.A(G20), .B(new_n569), .C1(new_n333), .C2(new_n318), .ZN(new_n578));
  OAI21_X1  g0378(.A(KEYINPUT86), .B1(new_n578), .B2(new_n568), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n573), .A2(new_n572), .A3(new_n574), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT24), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n582), .A3(new_n566), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n476), .B1(new_n577), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT25), .B1(new_n268), .B2(new_n203), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n268), .A2(KEYINPUT25), .A3(new_n203), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n478), .A2(G107), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n560), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n582), .B1(new_n581), .B2(new_n566), .ZN(new_n591));
  AOI211_X1 g0391(.A(KEYINPUT24), .B(new_n565), .C1(new_n579), .C2(new_n580), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n263), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n555), .A2(new_n296), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(G190), .B2(new_n555), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n588), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n267), .A2(new_n502), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n478), .B2(new_n502), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n465), .B(new_n208), .C1(G33), .C2(new_n202), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n502), .A2(G20), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n599), .A2(new_n263), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT20), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n263), .A3(new_n600), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT20), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n602), .A2(KEYINPUT85), .A3(new_n605), .ZN(new_n606));
  OR3_X1    g0406(.A1(new_n601), .A2(KEYINPUT85), .A3(KEYINPUT20), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n598), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  OR2_X1    g0408(.A1(G257), .A2(G1698), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(G264), .B2(new_n282), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n333), .B2(new_n318), .ZN(new_n611));
  INV_X1    g0411(.A(G303), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n280), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n285), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n446), .A2(G270), .B1(new_n448), .B2(new_n449), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n608), .A2(new_n616), .A3(KEYINPUT21), .A4(G169), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n608), .A2(G179), .A3(new_n614), .A4(new_n615), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n608), .B1(G200), .B2(new_n616), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n411), .B2(new_n616), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n608), .A2(new_n616), .A3(G169), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT21), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n619), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n590), .A2(new_n596), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n442), .A2(new_n547), .A3(new_n627), .ZN(G372));
  OAI21_X1  g0428(.A(new_n410), .B1(new_n414), .B2(new_n439), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n629), .A2(new_n378), .A3(new_n373), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n369), .A2(new_n375), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n307), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n310), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n509), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n531), .B1(new_n541), .B2(new_n511), .ZN(new_n636));
  AND4_X1   g0436(.A1(new_n531), .A2(new_n530), .A3(new_n511), .A4(new_n513), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT89), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT89), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n533), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n638), .A2(new_n488), .A3(new_n544), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n638), .A2(new_n488), .A3(new_n544), .A4(KEYINPUT26), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n642), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n596), .A2(new_n638), .A3(new_n544), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT88), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n559), .A2(new_n558), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(new_n556), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n651), .B1(new_n593), .B2(new_n588), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n619), .A2(new_n624), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n649), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n653), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n590), .A2(KEYINPUT88), .A3(new_n655), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n648), .A2(new_n654), .A3(new_n498), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n647), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n634), .B1(new_n442), .B2(new_n659), .ZN(G369));
  NAND3_X1  g0460(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT90), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(G343), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(G343), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n608), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n653), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n625), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n673), .B1(new_n674), .B2(new_n672), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n671), .B1(new_n584), .B2(new_n589), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n590), .A2(new_n678), .A3(new_n596), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n652), .A2(new_n671), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n590), .A2(new_n596), .A3(new_n653), .A4(new_n670), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n652), .A2(new_n670), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n682), .A2(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n211), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n204), .A2(G87), .A3(G116), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT91), .Z(new_n692));
  NAND3_X1  g0492(.A1(new_n690), .A2(new_n692), .A3(G1), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n214), .B2(new_n690), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT93), .ZN(new_n695));
  XNOR2_X1  g0495(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n504), .A2(new_n553), .A3(new_n506), .A4(new_n554), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n614), .A2(G179), .A3(new_n615), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n700), .A2(new_n469), .A3(KEYINPUT30), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT94), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT94), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n700), .A2(new_n469), .A3(new_n703), .A4(KEYINPUT30), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT95), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n700), .A2(new_n469), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  INV_X1    g0508(.A(new_n469), .ZN(new_n709));
  AND4_X1   g0509(.A1(new_n308), .A2(new_n555), .A3(new_n616), .A4(new_n507), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n707), .A2(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n705), .A2(new_n706), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n706), .B1(new_n705), .B2(new_n711), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(KEYINPUT31), .B1(new_n714), .B2(new_n671), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n705), .A2(new_n711), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n671), .A2(KEYINPUT31), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n590), .A2(new_n596), .A3(new_n625), .A4(new_n670), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n718), .B1(new_n547), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(G330), .B1(new_n715), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT96), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n639), .A2(new_n723), .A3(new_n641), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n526), .A2(new_n532), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n640), .B1(new_n725), .B2(new_n635), .ZN(new_n726));
  AOI211_X1 g0526(.A(KEYINPUT89), .B(new_n509), .C1(new_n526), .C2(new_n532), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT96), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n645), .A2(new_n646), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n590), .A2(new_n655), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n498), .A2(new_n731), .A3(new_n546), .A4(new_n596), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT97), .ZN(new_n734));
  AND3_X1   g0534(.A1(new_n733), .A2(new_n734), .A3(new_n670), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n734), .B1(new_n733), .B2(new_n670), .ZN(new_n736));
  OAI21_X1  g0536(.A(KEYINPUT29), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n671), .B1(new_n647), .B2(new_n657), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(KEYINPUT29), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n722), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n697), .B1(new_n741), .B2(G1), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT98), .ZN(G364));
  NAND2_X1  g0543(.A1(new_n208), .A2(G13), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT99), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G45), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(KEYINPUT100), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n207), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n746), .A2(KEYINPUT100), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n689), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n677), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(G330), .B2(new_n675), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n216), .B1(G20), .B2(new_n435), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n208), .A2(G179), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(G190), .A3(G200), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n756), .A2(new_n411), .A3(G200), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n758), .A2(G87), .B1(new_n760), .B2(G107), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n208), .A2(new_n308), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G190), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n761), .B1(new_n343), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G58), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n762), .A2(G190), .A3(new_n296), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n763), .A2(new_n411), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n280), .B1(new_n767), .B2(new_n768), .C1(new_n770), .C2(new_n250), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n411), .A2(new_n296), .A3(G20), .A4(G179), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT102), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n772), .A2(new_n773), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n766), .B(new_n771), .C1(new_n219), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n308), .A2(new_n296), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT103), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n781), .A2(new_n208), .A3(G190), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G159), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(KEYINPUT104), .B(KEYINPUT32), .ZN(new_n786));
  OAI21_X1  g0586(.A(G20), .B1(new_n781), .B2(new_n411), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n785), .A2(new_n786), .B1(G97), .B2(new_n787), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n779), .B(new_n788), .C1(new_n785), .C2(new_n786), .ZN(new_n789));
  INV_X1    g0589(.A(new_n768), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n280), .B1(new_n790), .B2(G322), .ZN(new_n791));
  XNOR2_X1  g0591(.A(KEYINPUT105), .B(G326), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n791), .B1(new_n770), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(G311), .B2(new_n778), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n787), .A2(G294), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n782), .A2(G329), .ZN(new_n796));
  INV_X1    g0596(.A(G283), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n797), .A2(new_n759), .B1(new_n757), .B2(new_n612), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT33), .B(G317), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n798), .B1(new_n764), .B2(new_n799), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n794), .A2(new_n795), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n755), .B1(new_n789), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G13), .A2(G33), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G20), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n754), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n247), .A2(G45), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT101), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n323), .A2(new_n688), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n809), .B(new_n810), .C1(G45), .C2(new_n214), .ZN(new_n811));
  INV_X1    g0611(.A(new_n280), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n688), .A2(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n813), .A2(G355), .B1(new_n502), .B2(new_n688), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n807), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n751), .ZN(new_n816));
  NOR3_X1   g0616(.A1(new_n802), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n805), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n675), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n753), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G396));
  NAND2_X1  g0621(.A1(new_n425), .A2(new_n671), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n434), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n439), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n437), .A2(new_n438), .A3(new_n670), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n738), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n654), .A2(new_n656), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n498), .A2(new_n546), .A3(new_n596), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n726), .A2(new_n727), .ZN(new_n832));
  AOI21_X1  g0632(.A(KEYINPUT26), .B1(new_n546), .B2(new_n488), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n470), .A2(new_n474), .A3(new_n487), .ZN(new_n834));
  NOR4_X1   g0634(.A1(new_n533), .A2(new_n545), .A3(new_n834), .A4(new_n644), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n832), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n670), .B(new_n827), .C1(new_n831), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n828), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n751), .B1(new_n838), .B2(new_n721), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n721), .B2(new_n838), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n754), .A2(new_n803), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n816), .B1(new_n382), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n759), .A2(new_n343), .ZN(new_n843));
  INV_X1    g0643(.A(new_n323), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n843), .B(new_n844), .C1(G50), .C2(new_n758), .ZN(new_n845));
  INV_X1    g0645(.A(new_n787), .ZN(new_n846));
  INV_X1    g0646(.A(G132), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n845), .B1(new_n767), .B2(new_n846), .C1(new_n847), .C2(new_n783), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT34), .ZN(new_n849));
  AOI22_X1  g0649(.A1(G137), .A2(new_n769), .B1(new_n790), .B2(G143), .ZN(new_n850));
  INV_X1    g0650(.A(G150), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n850), .B1(new_n851), .B2(new_n765), .C1(new_n777), .C2(new_n784), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n848), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n852), .A2(new_n849), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n777), .A2(new_n502), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n812), .B1(new_n551), .B2(new_n768), .C1(new_n770), .C2(new_n612), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n855), .B(new_n856), .C1(G311), .C2(new_n782), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n764), .A2(G283), .B1(new_n760), .B2(G87), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n203), .B2(new_n757), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n787), .B2(G97), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n853), .A2(new_n854), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n842), .B1(new_n755), .B2(new_n861), .C1(new_n827), .C2(new_n804), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n840), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(G384));
  INV_X1    g0664(.A(new_n483), .ZN(new_n865));
  OR2_X1    g0665(.A1(new_n865), .A2(KEYINPUT35), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(KEYINPUT35), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n866), .A2(G116), .A3(new_n217), .A4(new_n867), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT36), .Z(new_n869));
  OAI211_X1 g0669(.A(new_n219), .B(new_n215), .C1(new_n767), .C2(new_n343), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n250), .A2(G68), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n207), .B(G13), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n409), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n874), .A2(new_n407), .A3(new_n406), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n392), .B(new_n671), .C1(new_n875), .C2(new_n414), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n392), .A2(new_n671), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n410), .A2(new_n415), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n826), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n626), .A2(new_n498), .A3(new_n546), .A4(new_n670), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n716), .A2(KEYINPUT95), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n705), .A2(new_n706), .A3(new_n711), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(new_n882), .A3(new_n717), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n879), .B1(new_n715), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT107), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n879), .B(KEYINPUT107), .C1(new_n715), .C2(new_n884), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT38), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n379), .A2(new_n367), .A3(new_n665), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n367), .A2(new_n665), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n368), .A2(new_n891), .A3(new_n376), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT37), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n892), .B(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n889), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n263), .B1(new_n362), .B2(new_n342), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n844), .A2(new_n346), .A3(new_n208), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(G68), .A3(new_n359), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT16), .B1(new_n898), .B2(new_n355), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n366), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n665), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n379), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n368), .A2(new_n891), .A3(new_n893), .A4(new_n376), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n341), .A2(new_n900), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n905), .A2(new_n901), .A3(new_n376), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n904), .B1(new_n906), .B2(new_n893), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n903), .A2(new_n907), .A3(KEYINPUT38), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n895), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n887), .A2(KEYINPUT40), .A3(new_n888), .A4(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n903), .A2(new_n907), .A3(KEYINPUT38), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT38), .B1(new_n903), .B2(new_n907), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n911), .B1(new_n885), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n712), .A2(new_n713), .A3(new_n670), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n880), .B(new_n883), .C1(new_n917), .C2(KEYINPUT31), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n441), .A2(new_n918), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n916), .A2(new_n919), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n920), .A2(G330), .A3(new_n921), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT108), .Z(new_n923));
  NAND3_X1  g0723(.A1(new_n737), .A2(new_n441), .A3(new_n740), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT106), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n737), .A2(KEYINPUT106), .A3(new_n441), .A4(new_n740), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n633), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n631), .A2(new_n664), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT39), .B1(new_n895), .B2(new_n908), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT39), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n912), .A2(new_n913), .A3(new_n931), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n875), .A2(new_n392), .A3(new_n670), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n825), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n738), .B2(new_n827), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n876), .A2(new_n878), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NOR3_X1   g0739(.A1(new_n937), .A2(new_n914), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n935), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n928), .B(new_n941), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n923), .A2(new_n942), .B1(new_n207), .B2(new_n745), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT109), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n923), .A2(new_n942), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n943), .A2(KEYINPUT109), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n873), .B1(new_n946), .B2(new_n947), .ZN(G367));
  AND2_X1   g0748(.A1(new_n239), .A2(new_n810), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n806), .B1(new_n211), .B2(new_n417), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n751), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(G317), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n844), .B1(new_n202), .B2(new_n759), .C1(new_n783), .C2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT115), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n765), .A2(new_n551), .B1(new_n612), .B2(new_n768), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(G311), .B2(new_n769), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT46), .B1(new_n758), .B2(G116), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n778), .B2(G283), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n758), .A2(KEYINPUT46), .A3(G116), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n787), .A2(G107), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n956), .A2(new_n958), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n280), .B1(new_n768), .B2(new_n851), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(G58), .B2(new_n758), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n782), .A2(G137), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n963), .B(new_n964), .C1(new_n250), .C2(new_n777), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n787), .A2(G68), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n769), .A2(G143), .B1(new_n760), .B2(new_n219), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n966), .B(new_n967), .C1(new_n784), .C2(new_n765), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n954), .A2(new_n961), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT47), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n951), .B1(new_n970), .B2(new_n754), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n670), .B1(new_n541), .B2(new_n542), .ZN(new_n972));
  MUX2_X1   g0772(.A(new_n546), .B(new_n642), .S(new_n972), .Z(new_n973));
  OAI21_X1  g0773(.A(new_n971), .B1(new_n973), .B2(new_n818), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n487), .A2(new_n671), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n498), .A2(new_n975), .B1(new_n488), .B2(new_n671), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n976), .A2(new_n685), .B1(KEYINPUT111), .B2(KEYINPUT44), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(KEYINPUT111), .B(KEYINPUT44), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n976), .A2(new_n685), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n978), .A2(KEYINPUT112), .A3(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT112), .ZN(new_n982));
  INV_X1    g0782(.A(new_n980), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n982), .B1(new_n983), .B2(new_n977), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n498), .A2(new_n975), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n488), .A2(new_n671), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n686), .A2(new_n988), .A3(KEYINPUT45), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT45), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n976), .B2(new_n685), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n985), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n682), .B(KEYINPUT113), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n993), .A2(KEYINPUT114), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT114), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n981), .A2(new_n984), .B1(new_n989), .B2(new_n991), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n997), .B1(new_n998), .B2(new_n994), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n682), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n996), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n679), .B(new_n680), .C1(new_n655), .C2(new_n671), .ZN(new_n1002));
  AND3_X1   g0802(.A1(new_n1002), .A2(new_n676), .A3(new_n683), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n676), .B1(new_n1002), .B2(new_n683), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n741), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n741), .B1(new_n1001), .B2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n689), .B(KEYINPUT41), .Z(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n750), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(KEYINPUT42), .B1(new_n976), .B2(new_n683), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n590), .B1(new_n496), .B2(new_n497), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n670), .B1(new_n1013), .B2(new_n488), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  NOR3_X1   g0815(.A1(new_n976), .A2(KEYINPUT42), .A3(new_n683), .ZN(new_n1016));
  OR3_X1    g0816(.A1(new_n1015), .A2(KEYINPUT110), .A3(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n973), .B(KEYINPUT43), .ZN(new_n1018));
  OAI21_X1  g0818(.A(KEYINPUT110), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1019));
  AND3_X1   g0819(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n682), .A2(new_n976), .ZN(new_n1023));
  OR3_X1    g0823(.A1(new_n1020), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1023), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n974), .B1(new_n1011), .B2(new_n1026), .ZN(G387));
  AOI21_X1  g0827(.A(new_n690), .B1(new_n741), .B2(new_n1006), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n733), .A2(new_n670), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(KEYINPUT97), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n733), .A2(new_n734), .A3(new_n670), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n739), .B1(new_n1032), .B2(KEYINPUT29), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1005), .B1(new_n1033), .B2(new_n722), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1028), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n810), .B1(new_n235), .B2(new_n443), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n813), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1036), .B1(new_n692), .B2(new_n1037), .ZN(new_n1038));
  OR3_X1    g0838(.A1(new_n364), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1039));
  OAI21_X1  g0839(.A(KEYINPUT50), .B1(new_n364), .B2(G50), .ZN(new_n1040));
  AOI21_X1  g0840(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n692), .A2(new_n1039), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1038), .A2(new_n1042), .B1(new_n203), .B2(new_n688), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n751), .B1(new_n1043), .B2(new_n807), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n323), .B1(G116), .B2(new_n760), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n846), .A2(new_n797), .B1(new_n551), .B2(new_n757), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G311), .A2(new_n764), .B1(new_n790), .B2(G317), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n769), .A2(G322), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(new_n612), .C2(new_n777), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT48), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1046), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n1050), .B2(new_n1049), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT49), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1045), .B1(new_n783), .B2(new_n792), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n787), .A2(new_n510), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n250), .B2(new_n768), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT116), .Z(new_n1058));
  OAI221_X1 g0858(.A(new_n323), .B1(new_n343), .B2(new_n777), .C1(new_n783), .C2(new_n851), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n770), .A2(new_n784), .B1(new_n759), .B2(new_n202), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n765), .A2(new_n364), .B1(new_n220), .B2(new_n757), .ZN(new_n1061));
  OR3_X1    g0861(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n1054), .A2(new_n1055), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1044), .B1(new_n1063), .B2(new_n754), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n681), .B2(new_n818), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n750), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1065), .B1(new_n1005), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1035), .A2(new_n1068), .ZN(G393));
  AND2_X1   g0869(.A1(new_n244), .A2(new_n810), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n806), .B1(new_n202), .B2(new_n211), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n751), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n765), .A2(new_n612), .B1(new_n757), .B2(new_n797), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n280), .B(new_n1073), .C1(G107), .C2(new_n760), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G294), .A2(new_n778), .B1(new_n782), .B2(G322), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1074), .B(new_n1075), .C1(new_n502), .C2(new_n846), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G317), .A2(new_n769), .B1(new_n790), .B2(G311), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT52), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G150), .A2(new_n769), .B1(new_n790), .B2(G159), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(KEYINPUT117), .B(KEYINPUT51), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1079), .B(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n787), .A2(G77), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n765), .A2(new_n250), .B1(new_n759), .B2(new_n312), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G68), .B2(new_n758), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1081), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n782), .A2(G143), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1086), .B(new_n323), .C1(new_n364), .C2(new_n777), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n1076), .A2(new_n1078), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1072), .B1(new_n1088), .B2(new_n754), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n988), .B2(new_n818), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n993), .A2(new_n677), .A3(new_n681), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n1000), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1090), .B1(new_n1092), .B2(new_n1066), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n690), .B1(new_n1092), .B2(new_n1007), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n1033), .A2(new_n722), .A3(new_n1005), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1095), .A2(new_n996), .A3(new_n1000), .A4(new_n999), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1093), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(G390));
  AND2_X1   g0898(.A1(new_n918), .A2(G330), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n441), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n633), .B(new_n1101), .C1(new_n926), .C2(new_n927), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1030), .A2(new_n1031), .A3(new_n825), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(new_n824), .A3(new_n938), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n934), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n895), .B2(new_n908), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT118), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n939), .B1(new_n837), .B2(new_n825), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1108), .B1(new_n1109), .B2(new_n1105), .ZN(new_n1110));
  OAI211_X1 g0910(.A(KEYINPUT118), .B(new_n934), .C1(new_n937), .C2(new_n939), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1110), .A2(new_n933), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n879), .B(G330), .C1(new_n715), .C2(new_n884), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(KEYINPUT119), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT119), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n918), .A2(new_n1116), .A3(G330), .A4(new_n879), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1113), .A2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(G330), .B(new_n827), .C1(new_n715), .C2(new_n720), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n1120), .A2(new_n939), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1107), .A2(new_n1112), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n918), .A2(G330), .A3(new_n827), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n939), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n735), .A2(new_n736), .A3(new_n936), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n824), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1121), .B(new_n1124), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1120), .A2(new_n939), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1115), .A2(new_n1128), .A3(new_n1117), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n937), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1102), .A2(new_n1119), .A3(new_n1122), .A4(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n930), .A2(new_n932), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n934), .B1(new_n937), .B2(new_n939), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1134), .B1(new_n1135), .B2(new_n1108), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1136), .A2(new_n1111), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1118), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1122), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n926), .A2(new_n927), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1140), .A2(new_n1132), .A3(new_n634), .A4(new_n1100), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1133), .A2(new_n1142), .A3(new_n689), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1119), .A2(new_n750), .A3(new_n1122), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n841), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n751), .B1(new_n255), .B2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n770), .A2(new_n797), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n843), .B(new_n1147), .C1(G107), .C2(new_n764), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n782), .A2(G294), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n812), .B1(new_n757), .B2(new_n312), .C1(new_n502), .C2(new_n768), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n778), .B2(G97), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1148), .A2(new_n1082), .A3(new_n1149), .A4(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(G125), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n280), .B1(new_n250), .B2(new_n759), .C1(new_n783), .C2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT120), .ZN(new_n1155));
  INV_X1    g0955(.A(G128), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n770), .A2(new_n1156), .B1(new_n847), .B2(new_n768), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G137), .B2(new_n764), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n758), .A2(G150), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1159), .A2(KEYINPUT53), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT54), .B(G143), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n778), .A2(new_n1162), .B1(new_n1159), .B2(KEYINPUT53), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n787), .A2(G159), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1158), .A2(new_n1160), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1152), .B1(new_n1155), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1146), .B1(new_n1166), .B2(new_n754), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1134), .B2(new_n804), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n1144), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1143), .A2(new_n1169), .ZN(G378));
  NAND3_X1  g0970(.A1(new_n888), .A2(KEYINPUT40), .A3(new_n909), .ZN(new_n1171));
  AOI21_X1  g0971(.A(KEYINPUT107), .B1(new_n918), .B2(new_n879), .ZN(new_n1172));
  OAI211_X1 g0972(.A(G330), .B(new_n915), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT121), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n910), .A2(KEYINPUT121), .A3(G330), .A4(new_n915), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n311), .A2(new_n271), .A3(new_n665), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n271), .A2(new_n665), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n307), .A2(new_n310), .A3(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n1177), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1180), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1175), .A2(new_n1176), .A3(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1173), .B(new_n1174), .C1(new_n1181), .C2(new_n1182), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n941), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1184), .A2(new_n941), .A3(new_n1185), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1188), .A2(new_n750), .A3(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n751), .B1(G50), .B2(new_n1145), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n759), .A2(new_n767), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n765), .A2(new_n202), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(G116), .C2(new_n769), .ZN(new_n1194));
  INV_X1    g0994(.A(G41), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n768), .B2(new_n203), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1196), .B(new_n323), .C1(new_n219), .C2(new_n758), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n510), .A2(new_n778), .B1(new_n782), .B2(G283), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1194), .A2(new_n966), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT58), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1195), .B1(new_n844), .B2(new_n278), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1199), .A2(new_n1200), .B1(new_n250), .B2(new_n1201), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n770), .A2(new_n1153), .B1(new_n1156), .B2(new_n768), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n765), .A2(new_n847), .B1(new_n757), .B2(new_n1161), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(G137), .C2(new_n778), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n851), .B2(new_n846), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n278), .B(new_n1195), .C1(new_n759), .C2(new_n784), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n782), .B2(G124), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1202), .B1(new_n1200), .B2(new_n1199), .C1(new_n1210), .C2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1191), .B1(new_n1212), .B2(new_n754), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1183), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1213), .B1(new_n1214), .B2(new_n804), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1190), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(KEYINPUT106), .B1(new_n1033), .B2(new_n441), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n927), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n634), .B(new_n1100), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT122), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n928), .A2(KEYINPUT122), .A3(new_n1100), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1188), .A2(KEYINPUT57), .A3(new_n1189), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n689), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1221), .B(new_n1222), .C1(new_n1139), .C2(new_n1141), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1184), .A2(new_n941), .A3(new_n1185), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n941), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT57), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1216), .B1(new_n1227), .B2(new_n1232), .ZN(G375));
  NAND2_X1  g1033(.A1(new_n939), .A2(new_n803), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n751), .B1(G68), .B2(new_n1145), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1192), .B(new_n844), .C1(G137), .C2(new_n790), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n1156), .B2(new_n783), .C1(new_n851), .C2(new_n777), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n769), .A2(G132), .B1(new_n758), .B2(G159), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1238), .B1(new_n765), .B2(new_n1161), .C1(new_n846), .C2(new_n250), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n812), .B1(new_n768), .B2(new_n797), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G294), .B2(new_n769), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1241), .B1(new_n777), .B2(new_n203), .C1(new_n612), .C2(new_n783), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n758), .A2(G97), .B1(new_n760), .B2(G77), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1056), .B(new_n1243), .C1(new_n502), .C2(new_n765), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n1237), .A2(new_n1239), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1235), .B1(new_n1245), .B2(new_n754), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1132), .A2(new_n750), .B1(new_n1234), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1141), .A2(new_n1010), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1132), .B1(new_n928), .B2(new_n1100), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1247), .B1(new_n1248), .B2(new_n1249), .ZN(G381));
  OR4_X1    g1050(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n974), .B(new_n1097), .C1(new_n1011), .C2(new_n1026), .ZN(new_n1252));
  NOR4_X1   g1052(.A1(G375), .A2(new_n1251), .A3(G378), .A4(new_n1252), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1253), .B(KEYINPUT123), .ZN(G407));
  NAND2_X1  g1054(.A1(new_n1190), .A2(new_n1215), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1228), .A2(new_n1231), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT57), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1229), .A2(new_n1230), .A3(new_n1257), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n690), .B1(new_n1259), .B2(new_n1228), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1255), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(G378), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n667), .A2(new_n668), .A3(G213), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1261), .A2(new_n1262), .A3(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(G407), .A2(G213), .A3(new_n1265), .ZN(G409));
  OAI211_X1 g1066(.A(G378), .B(new_n1216), .C1(new_n1227), .C2(new_n1232), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1228), .A2(new_n1231), .A3(new_n1010), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1216), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1262), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1267), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1263), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1264), .A2(G2897), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1249), .B1(KEYINPUT60), .B2(new_n1141), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1132), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1219), .A2(KEYINPUT60), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n689), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G384), .B(new_n1247), .C1(new_n1275), .C2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1141), .A2(KEYINPUT60), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1219), .A2(new_n1276), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1283), .A2(new_n689), .A3(new_n1277), .ZN(new_n1284));
  AOI21_X1  g1084(.A(G384), .B1(new_n1284), .B2(new_n1247), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1274), .B1(new_n1280), .B2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1247), .B1(new_n1275), .B2(new_n1278), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n863), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(new_n1279), .A3(new_n1273), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1286), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1272), .A2(new_n1290), .A3(KEYINPUT125), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT125), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1264), .B1(new_n1267), .B2(new_n1270), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1286), .A2(new_n1289), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1292), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1291), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1288), .A2(new_n1279), .ZN(new_n1297));
  AOI211_X1 g1097(.A(new_n1264), .B(new_n1297), .C1(new_n1267), .C2(new_n1270), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(G393), .A2(G396), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT126), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n820), .B1(new_n1035), .B2(new_n1068), .ZN(new_n1301));
  NOR3_X1   g1101(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1300), .B1(new_n1299), .B2(new_n1301), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1252), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1026), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1009), .B1(new_n1096), .B2(new_n741), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1305), .B1(new_n1306), .B2(new_n750), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1097), .B1(new_n1307), .B2(new_n974), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1302), .B1(new_n1304), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT61), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(G387), .A2(G390), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1302), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1311), .A2(new_n1312), .A3(new_n1252), .A4(new_n1303), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1309), .A2(new_n1310), .A3(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT127), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1309), .A2(new_n1313), .A3(KEYINPUT127), .A4(new_n1310), .ZN(new_n1317));
  AOI22_X1  g1117(.A1(new_n1298), .A2(KEYINPUT63), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT124), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1319), .B1(new_n1298), .B2(KEYINPUT63), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1297), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1271), .A2(new_n1263), .A3(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT63), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1322), .A2(KEYINPUT124), .A3(new_n1323), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1296), .A2(new_n1318), .A3(new_n1320), .A4(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1322), .A2(KEYINPUT62), .ZN(new_n1326));
  AOI21_X1  g1126(.A(G378), .B1(new_n1216), .B2(new_n1268), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1327), .B1(new_n1261), .B2(G378), .ZN(new_n1328));
  OAI211_X1 g1128(.A(new_n1289), .B(new_n1286), .C1(new_n1328), .C2(new_n1264), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT62), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1293), .A2(new_n1330), .A3(new_n1321), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1326), .A2(new_n1310), .A3(new_n1329), .A4(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1309), .A2(new_n1313), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1325), .A2(new_n1334), .ZN(G405));
  NAND2_X1  g1135(.A1(G375), .A2(new_n1262), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1267), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(new_n1321), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1336), .A2(new_n1267), .A3(new_n1297), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  XNOR2_X1  g1140(.A(new_n1340), .B(new_n1333), .ZN(G402));
endmodule


