//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n573, new_n575, new_n576, new_n577, new_n578, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n598, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n631, new_n632, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT64), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G137), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT66), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(new_n460), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  INV_X1    g044(.A(new_n462), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(KEYINPUT65), .A2(G113), .A3(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(G2105), .B1(new_n472), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n479));
  INV_X1    g054(.A(G2104), .ZN(new_n480));
  NOR3_X1   g055(.A1(new_n479), .A2(new_n480), .A3(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  AOI21_X1  g057(.A(KEYINPUT67), .B1(new_n482), .B2(G2104), .ZN(new_n483));
  OAI21_X1  g058(.A(G101), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n468), .A2(new_n478), .A3(new_n484), .ZN(G160));
  AND2_X1   g060(.A1(new_n465), .A2(KEYINPUT68), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n465), .A2(KEYINPUT68), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  OAI21_X1  g065(.A(G2105), .B1(new_n486), .B2(new_n487), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n482), .A2(G112), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n490), .B(new_n493), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G162));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n502), .B1(new_n461), .B2(new_n462), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n502), .B(new_n505), .C1(new_n462), .C2(new_n461), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n500), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(G126), .A2(G2105), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n508), .B1(new_n461), .B2(new_n462), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT69), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n465), .A2(KEYINPUT69), .A3(new_n508), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(G164));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  OR2_X1    g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G50), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT70), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n520), .B(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  AND2_X1   g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G62), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OR2_X1    g103(.A1(KEYINPUT5), .A2(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(KEYINPUT5), .A2(G543), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n517), .A2(new_n518), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n528), .A2(G651), .B1(new_n531), .B2(G88), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n522), .A2(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT72), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT72), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n537), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT7), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n536), .A2(new_n541), .A3(new_n538), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(G63), .A2(G651), .ZN(new_n544));
  AND2_X1   g119(.A1(KEYINPUT6), .A2(G651), .ZN(new_n545));
  NOR2_X1   g120(.A1(KEYINPUT6), .A2(G651), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(G89), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  XNOR2_X1  g124(.A(KEYINPUT5), .B(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g126(.A(KEYINPUT71), .B(G51), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n519), .A2(new_n552), .ZN(new_n553));
  AND3_X1   g128(.A1(new_n543), .A2(new_n551), .A3(new_n553), .ZN(G168));
  XNOR2_X1  g129(.A(KEYINPUT6), .B(G651), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n555), .A2(new_n550), .A3(G90), .ZN(new_n556));
  OAI211_X1 g131(.A(G52), .B(G543), .C1(new_n545), .C2(new_n546), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(G651), .ZN(new_n559));
  OAI21_X1  g134(.A(G64), .B1(new_n524), .B2(new_n525), .ZN(new_n560));
  NAND2_X1  g135(.A1(G77), .A2(G543), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n558), .A2(new_n562), .ZN(G171));
  NAND3_X1  g138(.A1(new_n555), .A2(G43), .A3(G543), .ZN(new_n564));
  INV_X1    g139(.A(G81), .ZN(new_n565));
  OAI22_X1  g140(.A1(new_n546), .A2(new_n545), .B1(new_n524), .B2(new_n525), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n550), .A2(G56), .ZN(new_n568));
  NAND2_X1  g143(.A1(G68), .A2(G543), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n559), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G860), .ZN(G153));
  AND3_X1   g147(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G36), .ZN(G176));
  NAND2_X1  g149(.A1(G1), .A2(G3), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT74), .ZN(new_n576));
  XOR2_X1   g151(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n577));
  XNOR2_X1  g152(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n573), .A2(new_n578), .ZN(G188));
  NAND2_X1  g154(.A1(G78), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G65), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n526), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(new_n531), .B2(G91), .ZN(new_n583));
  OAI211_X1 g158(.A(G53), .B(G543), .C1(new_n545), .C2(new_n546), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT9), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT9), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n555), .A2(new_n586), .A3(G53), .A4(G543), .ZN(new_n587));
  AND3_X1   g162(.A1(new_n585), .A2(new_n587), .A3(KEYINPUT75), .ZN(new_n588));
  AOI21_X1  g163(.A(KEYINPUT75), .B1(new_n585), .B2(new_n587), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n583), .B1(new_n588), .B2(new_n589), .ZN(G299));
  INV_X1    g165(.A(KEYINPUT76), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n591), .B1(new_n558), .B2(new_n562), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n560), .A2(new_n561), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G651), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n594), .A2(KEYINPUT76), .A3(new_n557), .A4(new_n556), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G301));
  AOI22_X1  g172(.A1(new_n549), .A2(new_n550), .B1(new_n519), .B2(new_n552), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(new_n543), .ZN(G286));
  NAND2_X1  g174(.A1(new_n531), .A2(G87), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n550), .B2(G74), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n519), .A2(G49), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(G288));
  NAND3_X1  g178(.A1(new_n555), .A2(new_n550), .A3(G86), .ZN(new_n604));
  OAI211_X1 g179(.A(G48), .B(G543), .C1(new_n545), .C2(new_n546), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(G61), .B1(new_n524), .B2(new_n525), .ZN(new_n607));
  NAND2_X1  g182(.A1(G73), .A2(G543), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n559), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(G305));
  NAND2_X1  g186(.A1(new_n519), .A2(G47), .ZN(new_n612));
  INV_X1    g187(.A(G85), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n550), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n614));
  OAI221_X1 g189(.A(new_n612), .B1(new_n613), .B2(new_n566), .C1(new_n614), .C2(new_n559), .ZN(G290));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  INV_X1    g191(.A(G92), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n566), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g193(.A1(new_n555), .A2(new_n550), .A3(KEYINPUT10), .A4(G92), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n519), .A2(G54), .ZN(new_n621));
  INV_X1    g196(.A(G66), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n526), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(G79), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n624), .A2(new_n516), .ZN(new_n625));
  OAI21_X1  g200(.A(G651), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n620), .A2(new_n621), .A3(new_n626), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(G868), .B2(new_n596), .ZN(G284));
  AOI21_X1  g204(.A(new_n628), .B1(G868), .B2(new_n596), .ZN(G321));
  INV_X1    g205(.A(G868), .ZN(new_n631));
  NAND2_X1  g206(.A1(G299), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n631), .B2(G168), .ZN(G297));
  OAI21_X1  g208(.A(new_n632), .B1(new_n631), .B2(G168), .ZN(G280));
  AOI21_X1  g209(.A(new_n625), .B1(new_n550), .B2(G66), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n621), .B1(new_n635), .B2(new_n559), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n636), .B1(new_n618), .B2(new_n619), .ZN(new_n637));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(G860), .ZN(G148));
  NAND2_X1  g214(.A1(new_n531), .A2(G81), .ZN(new_n640));
  AOI22_X1  g215(.A1(new_n550), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n640), .B(new_n564), .C1(new_n559), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(new_n631), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n627), .A2(G559), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n643), .B1(new_n644), .B2(new_n631), .ZN(G323));
  XNOR2_X1  g220(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g221(.A1(new_n481), .A2(new_n483), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(new_n465), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT12), .Z(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT13), .Z(new_n650));
  INV_X1    g225(.A(G2100), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT77), .ZN(new_n653));
  INV_X1    g228(.A(G2096), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n489), .A2(G135), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n492), .A2(G123), .ZN(new_n656));
  OR2_X1    g231(.A1(G99), .A2(G2105), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n657), .B(G2104), .C1(G111), .C2(new_n482), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  AOI22_X1  g235(.A1(new_n650), .A2(new_n651), .B1(new_n654), .B2(new_n660), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n653), .B(new_n661), .C1(new_n654), .C2(new_n660), .ZN(G156));
  XNOR2_X1  g237(.A(G2427), .B(G2438), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2430), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT15), .B(G2435), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(KEYINPUT14), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1341), .B(G1348), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2443), .B(G2446), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT79), .ZN(new_n674));
  XOR2_X1   g249(.A(G2451), .B(G2454), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n672), .A2(new_n676), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n677), .A2(G14), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT80), .Z(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G401));
  XOR2_X1   g256(.A(G2084), .B(G2090), .Z(new_n682));
  XNOR2_X1  g257(.A(G2067), .B(G2678), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2072), .B(G2078), .Z(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT82), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT81), .B(KEYINPUT18), .Z(new_n688));
  OR2_X1    g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  OAI21_X1  g265(.A(KEYINPUT17), .B1(new_n682), .B2(new_n683), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n691), .A2(new_n685), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n685), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n692), .A2(new_n684), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n689), .A2(new_n690), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G2096), .B(G2100), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G227));
  XOR2_X1   g272(.A(G1991), .B(G1996), .Z(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1956), .B(G2474), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT83), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1961), .B(G1966), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1971), .B(G1976), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT19), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT20), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n703), .A2(new_n704), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n711), .A2(new_n707), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT84), .Z(new_n713));
  NAND3_X1  g288(.A1(new_n705), .A2(new_n711), .A3(new_n707), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n710), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(KEYINPUT85), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n715), .A2(KEYINPUT85), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n701), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n718), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n720), .A2(new_n716), .A3(new_n700), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n699), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(G1981), .B(G1986), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n719), .A2(new_n721), .A3(new_n699), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n724), .ZN(new_n727));
  INV_X1    g302(.A(new_n725), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(new_n722), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n726), .A2(new_n729), .ZN(G229));
  INV_X1    g305(.A(G16), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G22), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G166), .B2(new_n731), .ZN(new_n733));
  INV_X1    g308(.A(G1971), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(G16), .A2(G23), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT88), .Z(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G288), .B2(new_n731), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT33), .B(G1976), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n735), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n731), .A2(G6), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n610), .B2(new_n731), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT87), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT32), .B(G1981), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  OR3_X1    g321(.A1(new_n741), .A2(KEYINPUT34), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G25), .A2(G29), .ZN(new_n748));
  OAI21_X1  g323(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n749));
  INV_X1    g324(.A(G107), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(G2105), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n489), .B2(G131), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT86), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n492), .B2(G119), .ZN(new_n754));
  INV_X1    g329(.A(G119), .ZN(new_n755));
  NOR3_X1   g330(.A1(new_n491), .A2(KEYINPUT86), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n752), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n748), .B1(new_n758), .B2(G29), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT35), .B(G1991), .Z(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n759), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n731), .A2(G24), .ZN(new_n763));
  INV_X1    g338(.A(G290), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n731), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1986), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(KEYINPUT34), .B1(new_n741), .B2(new_n746), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n747), .A2(new_n767), .A3(KEYINPUT90), .A4(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT89), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n747), .A2(new_n767), .A3(new_n768), .ZN(new_n773));
  OAI21_X1  g348(.A(KEYINPUT36), .B1(new_n773), .B2(new_n770), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n771), .A2(KEYINPUT36), .ZN(new_n776));
  NOR2_X1   g351(.A1(KEYINPUT96), .A2(G2090), .ZN(new_n777));
  INV_X1    g352(.A(G29), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G35), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G162), .B2(new_n778), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n780), .A2(KEYINPUT29), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(KEYINPUT29), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n777), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(KEYINPUT96), .A2(G2090), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n778), .A2(G32), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n489), .A2(G141), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n492), .A2(G129), .ZN(new_n788));
  NAND3_X1  g363(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT26), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n647), .A2(G105), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n787), .A2(new_n788), .A3(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n786), .B1(new_n795), .B2(new_n778), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT27), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1996), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n571), .A2(G16), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G16), .B2(G19), .ZN(new_n800));
  INV_X1    g375(.A(G1341), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(KEYINPUT31), .A2(G11), .ZN(new_n803));
  AND2_X1   g378(.A1(KEYINPUT31), .A2(G11), .ZN(new_n804));
  INV_X1    g379(.A(G28), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(KEYINPUT30), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT30), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n778), .B1(new_n807), .B2(G28), .ZN(new_n808));
  OAI221_X1 g383(.A(new_n802), .B1(new_n803), .B2(new_n804), .C1(new_n806), .C2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n637), .A2(G16), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G4), .B2(G16), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n809), .B1(G1348), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(G29), .A2(G33), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT92), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n489), .A2(G139), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT93), .B(KEYINPUT25), .Z(new_n817));
  NAND3_X1  g392(.A1(new_n482), .A2(G103), .A3(G2104), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n816), .B(new_n819), .C1(new_n482), .C2(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n815), .B1(new_n821), .B2(new_n778), .ZN(new_n822));
  INV_X1    g397(.A(G2072), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(G160), .A2(G29), .ZN(new_n825));
  INV_X1    g400(.A(G34), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n826), .A2(KEYINPUT24), .ZN(new_n827));
  AOI21_X1  g402(.A(G29), .B1(new_n826), .B2(KEYINPUT24), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n827), .B1(new_n828), .B2(KEYINPUT94), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(KEYINPUT94), .B2(new_n828), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n825), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n824), .B1(G2084), .B2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G2078), .ZN(new_n834));
  NAND2_X1  g409(.A1(G164), .A2(G29), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(G27), .B2(G29), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n822), .A2(new_n823), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n659), .A2(new_n778), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n731), .A2(G5), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(G171), .B2(new_n731), .ZN(new_n840));
  OAI22_X1  g415(.A1(new_n800), .A2(new_n801), .B1(G1961), .B2(new_n840), .ZN(new_n841));
  AOI211_X1 g416(.A(new_n838), .B(new_n841), .C1(G1961), .C2(new_n840), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n813), .A2(new_n833), .A3(new_n837), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n731), .A2(G20), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT23), .Z(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(G299), .B2(G16), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(G1956), .Z(new_n847));
  NOR2_X1   g422(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(G16), .A2(G21), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(G168), .B2(G16), .ZN(new_n850));
  INV_X1    g425(.A(G1966), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  OAI221_X1 g427(.A(new_n852), .B1(new_n834), .B2(new_n836), .C1(G1348), .C2(new_n812), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n778), .A2(G26), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT28), .Z(new_n855));
  OR2_X1    g430(.A1(G104), .A2(G2105), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n856), .B(G2104), .C1(G116), .C2(new_n482), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT91), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n858), .B1(new_n492), .B2(G128), .ZN(new_n859));
  INV_X1    g434(.A(G140), .ZN(new_n860));
  INV_X1    g435(.A(new_n489), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n855), .B1(new_n862), .B2(G29), .ZN(new_n863));
  INV_X1    g438(.A(G2067), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G2084), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n831), .A2(new_n866), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT95), .Z(new_n868));
  NOR3_X1   g443(.A1(new_n853), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  AND4_X1   g444(.A1(new_n785), .A2(new_n798), .A3(new_n848), .A4(new_n869), .ZN(new_n870));
  AND3_X1   g445(.A1(new_n775), .A2(new_n776), .A3(new_n870), .ZN(G311));
  NAND3_X1  g446(.A1(new_n775), .A2(new_n776), .A3(new_n870), .ZN(G150));
  INV_X1    g447(.A(KEYINPUT97), .ZN(new_n873));
  OAI211_X1 g448(.A(G55), .B(G543), .C1(new_n545), .C2(new_n546), .ZN(new_n874));
  INV_X1    g449(.A(G93), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n874), .B1(new_n566), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(G67), .B1(new_n524), .B2(new_n525), .ZN(new_n877));
  NAND2_X1  g452(.A1(G80), .A2(G543), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n559), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n873), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(G67), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n881), .B1(new_n529), .B2(new_n530), .ZN(new_n882));
  INV_X1    g457(.A(new_n878), .ZN(new_n883));
  OAI21_X1  g458(.A(G651), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n555), .A2(new_n550), .A3(G93), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n884), .A2(KEYINPUT97), .A3(new_n874), .A4(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n571), .A2(new_n880), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n874), .A3(new_n885), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n642), .A2(new_n873), .A3(new_n888), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT38), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n637), .A2(G559), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n893), .A2(KEYINPUT39), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(KEYINPUT39), .ZN(new_n895));
  XOR2_X1   g470(.A(KEYINPUT98), .B(G860), .Z(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n888), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n898), .A2(new_n896), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT37), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(G145));
  XNOR2_X1  g476(.A(new_n795), .B(new_n821), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT100), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n757), .B(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n649), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n757), .B(KEYINPUT100), .ZN(new_n907));
  INV_X1    g482(.A(new_n649), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n903), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n862), .B(new_n514), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n489), .A2(G142), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n492), .A2(G130), .ZN(new_n914));
  NOR3_X1   g489(.A1(new_n482), .A2(KEYINPUT99), .A3(G118), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT99), .B1(new_n482), .B2(G118), .ZN(new_n916));
  OR2_X1    g491(.A1(G106), .A2(G2105), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(G2104), .A3(new_n917), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n913), .B(new_n914), .C1(new_n915), .C2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n912), .B(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n906), .A2(new_n909), .A3(new_n903), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n911), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n920), .ZN(new_n923));
  INV_X1    g498(.A(new_n921), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n923), .B1(new_n924), .B2(new_n910), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n660), .B(new_n496), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(G160), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G37), .ZN(new_n930));
  INV_X1    g505(.A(new_n928), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n922), .A2(new_n925), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g509(.A(new_n890), .B(new_n644), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n585), .A2(new_n587), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT75), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n585), .A2(new_n587), .A3(KEYINPUT75), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(new_n627), .A3(new_n583), .ZN(new_n941));
  NAND2_X1  g516(.A1(G299), .A2(new_n637), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n935), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT101), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(G299), .B2(new_n637), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n940), .A2(new_n627), .A3(KEYINPUT101), .A4(new_n583), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(new_n942), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT41), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n949), .B1(G299), .B2(new_n637), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n948), .A2(new_n949), .B1(new_n941), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n944), .B1(new_n951), .B2(new_n935), .ZN(new_n952));
  NOR2_X1   g527(.A1(KEYINPUT102), .A2(KEYINPUT42), .ZN(new_n953));
  OR2_X1    g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n953), .ZN(new_n955));
  INV_X1    g530(.A(G288), .ZN(new_n956));
  NAND2_X1  g531(.A1(G305), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n610), .A2(G288), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n522), .A2(G290), .A3(new_n532), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(G290), .B1(new_n522), .B2(new_n532), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(G303), .A2(new_n764), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n964), .A2(new_n957), .A3(new_n958), .A4(new_n960), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(KEYINPUT102), .A2(KEYINPUT42), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n954), .A2(new_n955), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n970), .B1(new_n954), .B2(new_n955), .ZN(new_n972));
  OAI21_X1  g547(.A(G868), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n898), .A2(G868), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(new_n975), .ZN(G295));
  NAND2_X1  g551(.A1(G295), .A2(KEYINPUT103), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT103), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n973), .A2(new_n978), .A3(new_n975), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(G331));
  INV_X1    g555(.A(KEYINPUT107), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT104), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n531), .A2(G90), .B1(new_n519), .B2(G52), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n598), .A2(new_n543), .B1(new_n983), .B2(new_n594), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(new_n596), .B2(G168), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n982), .B1(new_n890), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n887), .A2(new_n889), .ZN(new_n987));
  AOI21_X1  g562(.A(G286), .B1(new_n592), .B2(new_n595), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n987), .B1(new_n988), .B2(new_n984), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n596), .A2(G168), .ZN(new_n990));
  INV_X1    g565(.A(new_n984), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n990), .A2(new_n991), .A3(new_n889), .A4(new_n887), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n986), .B1(new_n993), .B2(new_n982), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT105), .B1(new_n994), .B2(new_n951), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n948), .A2(new_n949), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n950), .A2(new_n941), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT105), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT104), .B1(new_n989), .B2(new_n992), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n998), .B(new_n999), .C1(new_n1000), .C2(new_n986), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n995), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n943), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n966), .B1(new_n993), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n981), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  AOI211_X1 g581(.A(KEYINPUT107), .B(new_n1004), .C1(new_n995), .C2(new_n1001), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n993), .A2(new_n1003), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1009), .B1(new_n995), .B2(new_n1001), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n963), .A2(new_n965), .A3(KEYINPUT106), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT106), .B1(new_n963), .B2(new_n965), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n930), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT43), .B1(new_n1008), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n994), .A2(new_n943), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1003), .A2(KEYINPUT41), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n946), .A2(new_n950), .A3(new_n947), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n993), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1013), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1020), .A2(KEYINPUT43), .A3(G37), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT108), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1021), .B(KEYINPUT108), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1015), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OR2_X1    g603(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1014), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT43), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1020), .A2(G37), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT43), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1008), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT44), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1028), .A2(new_n1035), .ZN(G397));
  INV_X1    g611(.A(G1384), .ZN(new_n1037));
  INV_X1    g612(.A(new_n500), .ZN(new_n1038));
  INV_X1    g613(.A(new_n506), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n505), .B1(new_n465), .B2(new_n502), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1038), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n511), .A2(new_n512), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1037), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n468), .A2(new_n478), .A3(G40), .A4(new_n484), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n862), .B(new_n864), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1048), .B1(new_n1049), .B2(new_n795), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT46), .B1(new_n1048), .B2(G1996), .ZN(new_n1051));
  OR3_X1    g626(.A1(new_n1048), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1050), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1053), .B(KEYINPUT47), .ZN(new_n1054));
  INV_X1    g629(.A(G1986), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1047), .A2(new_n1055), .A3(new_n764), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1056), .B(KEYINPUT126), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT48), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1060));
  XOR2_X1   g635(.A(new_n794), .B(G1996), .Z(new_n1061));
  AND2_X1   g636(.A1(new_n1061), .A2(new_n1049), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n758), .A2(new_n760), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n757), .A2(new_n761), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  AOI211_X1 g640(.A(new_n1059), .B(new_n1060), .C1(new_n1047), .C2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1063), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1062), .B1(KEYINPUT125), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT125), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1063), .A2(new_n1069), .ZN(new_n1070));
  OAI22_X1  g645(.A1(new_n1068), .A2(new_n1070), .B1(G2067), .B2(new_n862), .ZN(new_n1071));
  AOI211_X1 g646(.A(new_n1054), .B(new_n1066), .C1(new_n1047), .C2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n600), .A2(G1976), .A3(new_n601), .A4(new_n602), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1073), .B(KEYINPUT112), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT111), .ZN(new_n1075));
  AND4_X1   g650(.A1(G40), .A2(new_n468), .A3(new_n478), .A4(new_n484), .ZN(new_n1076));
  AOI21_X1  g651(.A(G1384), .B1(new_n507), .B2(new_n513), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1075), .B1(new_n1078), .B2(G8), .ZN(new_n1079));
  INV_X1    g654(.A(G8), .ZN(new_n1080));
  AOI211_X1 g655(.A(KEYINPUT111), .B(new_n1080), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1074), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT113), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(G8), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT111), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1078), .A2(new_n1075), .A3(G8), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1088), .A2(KEYINPUT113), .A3(new_n1074), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1084), .A2(KEYINPUT52), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(G303), .A2(G8), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT55), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1091), .B(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G2090), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1077), .A2(KEYINPUT50), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT50), .ZN(new_n1096));
  AOI211_X1 g671(.A(new_n1096), .B(G1384), .C1(new_n507), .C2(new_n513), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1094), .B(new_n1076), .C1(new_n1095), .C2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1046), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1077), .A2(KEYINPUT45), .ZN(new_n1100));
  AOI21_X1  g675(.A(G1971), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT110), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1098), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  AOI211_X1 g678(.A(KEYINPUT110), .B(G1971), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1104));
  OAI211_X1 g679(.A(G8), .B(new_n1093), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(G1981), .B1(new_n606), .B2(new_n609), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  OAI211_X1 g683(.A(KEYINPUT116), .B(G1981), .C1(new_n606), .C2(new_n609), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G61), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(new_n529), .B2(new_n530), .ZN(new_n1112));
  INV_X1    g687(.A(new_n608), .ZN(new_n1113));
  OAI21_X1  g688(.A(G651), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT114), .B(G1981), .Z(new_n1115));
  NAND4_X1  g690(.A1(new_n1114), .A2(new_n604), .A3(new_n605), .A4(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT115), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n604), .A2(new_n605), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT115), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1118), .A2(new_n1119), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1110), .A2(new_n1121), .A3(KEYINPUT49), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT117), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT117), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1110), .A2(new_n1121), .A3(new_n1124), .A4(KEYINPUT49), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1110), .A2(new_n1121), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT49), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1086), .A2(new_n1087), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1074), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1130), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1131));
  INV_X1    g706(.A(G1976), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT52), .B1(G288), .B2(new_n1132), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1126), .A2(new_n1129), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1091), .B(KEYINPUT55), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1043), .A2(new_n1096), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1077), .A2(KEYINPUT50), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1046), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1045), .A2(new_n1100), .A3(new_n1076), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1094), .A2(new_n1138), .B1(new_n1139), .B2(new_n734), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1135), .B1(new_n1140), .B2(new_n1080), .ZN(new_n1141));
  AND4_X1   g716(.A1(new_n1090), .A2(new_n1105), .A3(new_n1134), .A4(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT51), .ZN(new_n1143));
  NOR2_X1   g718(.A1(G168), .A2(new_n1080), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT121), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1044), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1037), .B(new_n1146), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1147), .B(new_n1076), .C1(KEYINPUT45), .C2(new_n1077), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1138), .A2(new_n866), .B1(new_n1148), .B2(new_n851), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1143), .B(new_n1145), .C1(new_n1149), .C2(new_n1080), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT51), .B1(new_n1149), .B2(new_n1145), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1144), .B(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1148), .A2(new_n851), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n866), .B(new_n1076), .C1(new_n1095), .C2(new_n1097), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1153), .B1(new_n1156), .B2(G8), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1150), .B1(new_n1151), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT53), .ZN(new_n1161));
  OR3_X1    g736(.A1(new_n1148), .A2(new_n1161), .A3(G2078), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1076), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1163));
  INV_X1    g738(.A(G1961), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1161), .B1(new_n1139), .B2(G2078), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1162), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n596), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1168), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1150), .B(KEYINPUT62), .C1(new_n1151), .C2(new_n1157), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1142), .A2(new_n1160), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(KEYINPUT124), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n956), .A2(new_n1132), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1173), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1121), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1088), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT52), .B1(new_n1131), .B2(KEYINPUT113), .ZN(new_n1179));
  AOI211_X1 g754(.A(new_n1083), .B(new_n1130), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1177), .B(new_n1178), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1176), .B1(new_n1181), .B2(new_n1105), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(KEYINPUT118), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT118), .ZN(new_n1184));
  OAI211_X1 g759(.A(new_n1176), .B(new_n1184), .C1(new_n1181), .C2(new_n1105), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1181), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1156), .A2(G8), .A3(G168), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT63), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(G8), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(new_n1135), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1187), .A2(new_n1105), .A3(new_n1190), .A4(new_n1192), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1090), .A2(new_n1105), .A3(new_n1134), .A4(new_n1141), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1189), .B1(new_n1194), .B2(new_n1188), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1172), .A2(new_n1186), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT124), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1160), .A2(new_n1198), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1199));
  OAI22_X1  g774(.A1(new_n1138), .A2(G1348), .B1(G2067), .B2(new_n1078), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT120), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  OAI221_X1 g777(.A(KEYINPUT120), .B1(G2067), .B2(new_n1078), .C1(new_n1138), .C2(G1348), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n627), .B1(new_n1204), .B2(KEYINPUT60), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT60), .ZN(new_n1206));
  AOI211_X1 g781(.A(new_n1206), .B(new_n637), .C1(new_n1202), .C2(new_n1203), .ZN(new_n1207));
  OAI22_X1  g782(.A1(new_n1205), .A2(new_n1207), .B1(KEYINPUT60), .B2(new_n1204), .ZN(new_n1208));
  XOR2_X1   g783(.A(KEYINPUT58), .B(G1341), .Z(new_n1209));
  NAND2_X1  g784(.A1(new_n1078), .A2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1210), .B1(new_n1139), .B2(G1996), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1211), .A2(new_n571), .ZN(new_n1212));
  XNOR2_X1  g787(.A(new_n1212), .B(KEYINPUT59), .ZN(new_n1213));
  XOR2_X1   g788(.A(KEYINPUT56), .B(G2072), .Z(new_n1214));
  OAI22_X1  g789(.A1(new_n1138), .A2(G1956), .B1(new_n1139), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT57), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n583), .B1(KEYINPUT119), .B2(new_n936), .ZN(new_n1217));
  AND2_X1   g792(.A1(new_n936), .A2(KEYINPUT119), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1216), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n940), .A2(KEYINPUT57), .A3(new_n583), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g796(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1215), .A2(new_n1222), .ZN(new_n1223));
  OAI221_X1 g798(.A(new_n1221), .B1(new_n1139), .B2(new_n1214), .C1(G1956), .C2(new_n1138), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g800(.A(KEYINPUT61), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1223), .A2(new_n1224), .A3(KEYINPUT61), .ZN(new_n1228));
  AND3_X1   g803(.A1(new_n1213), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  OAI21_X1  g804(.A(new_n1223), .B1(new_n1204), .B2(new_n627), .ZN(new_n1230));
  AOI22_X1  g805(.A1(new_n1208), .A2(new_n1229), .B1(new_n1230), .B2(new_n1224), .ZN(new_n1231));
  INV_X1    g806(.A(KEYINPUT54), .ZN(new_n1232));
  INV_X1    g807(.A(new_n1167), .ZN(new_n1233));
  AOI21_X1  g808(.A(new_n1232), .B1(new_n1233), .B2(G301), .ZN(new_n1234));
  NAND4_X1  g809(.A1(new_n1099), .A2(KEYINPUT53), .A3(new_n834), .A4(new_n1100), .ZN(new_n1235));
  AND3_X1   g810(.A1(new_n1163), .A2(KEYINPUT122), .A3(new_n1164), .ZN(new_n1236));
  AOI21_X1  g811(.A(KEYINPUT122), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1237));
  OAI211_X1 g812(.A(new_n1166), .B(new_n1235), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1238));
  INV_X1    g813(.A(KEYINPUT123), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g815(.A1(new_n1240), .A2(G171), .ZN(new_n1241));
  NOR2_X1   g816(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1242));
  OAI21_X1  g817(.A(new_n1234), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g818(.A(new_n1168), .B1(new_n1238), .B2(new_n596), .ZN(new_n1244));
  AOI21_X1  g819(.A(new_n1158), .B1(new_n1244), .B2(new_n1232), .ZN(new_n1245));
  NAND2_X1  g820(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g821(.A(new_n1199), .B1(new_n1231), .B2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g822(.A(new_n1197), .B1(new_n1247), .B2(new_n1142), .ZN(new_n1248));
  INV_X1    g823(.A(new_n1065), .ZN(new_n1249));
  XNOR2_X1  g824(.A(G290), .B(new_n1055), .ZN(new_n1250));
  AOI21_X1  g825(.A(new_n1048), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g826(.A(new_n1072), .B1(new_n1248), .B2(new_n1251), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g827(.A(G319), .ZN(new_n1254));
  NOR2_X1   g828(.A1(G227), .A2(new_n1254), .ZN(new_n1255));
  XNOR2_X1  g829(.A(new_n1255), .B(KEYINPUT127), .ZN(new_n1256));
  NAND2_X1  g830(.A1(new_n1256), .A2(new_n680), .ZN(new_n1257));
  AOI21_X1  g831(.A(new_n1257), .B1(new_n726), .B2(new_n729), .ZN(new_n1258));
  AND3_X1   g832(.A1(new_n1026), .A2(new_n933), .A3(new_n1258), .ZN(G308));
  NAND3_X1  g833(.A1(new_n1026), .A2(new_n1258), .A3(new_n933), .ZN(G225));
endmodule


