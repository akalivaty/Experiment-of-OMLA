//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974;
  INV_X1    g000(.A(G227gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT24), .ZN(new_n206));
  INV_X1    g005(.A(G183gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G190gat), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G183gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n206), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n206), .A2(G183gat), .A3(G190gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n205), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G183gat), .B(G190gat), .ZN(new_n215));
  OAI211_X1 g014(.A(KEYINPUT64), .B(new_n212), .C1(new_n215), .C2(new_n206), .ZN(new_n216));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n220));
  INV_X1    g019(.A(G169gat), .ZN(new_n221));
  INV_X1    g020(.A(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n219), .A2(new_n220), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(new_n223), .B2(new_n224), .ZN(new_n227));
  NOR2_X1   g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n228), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n214), .A2(new_n216), .A3(new_n225), .A4(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT25), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n232), .B1(new_n228), .B2(KEYINPUT23), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n225), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n212), .B1(new_n215), .B2(new_n206), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n233), .A2(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n241));
  OAI21_X1  g040(.A(G134gat), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(G127gat), .ZN(new_n243));
  INV_X1    g042(.A(G134gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G113gat), .B(G120gat), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n242), .B(new_n245), .C1(KEYINPUT1), .C2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G120gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(G113gat), .ZN(new_n249));
  INV_X1    g048(.A(G113gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G120gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n249), .A2(new_n251), .A3(KEYINPUT69), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT1), .ZN(new_n253));
  XNOR2_X1  g052(.A(G127gat), .B(G134gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(new_n248), .A3(G113gat), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n252), .A2(new_n253), .A3(new_n254), .A4(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n247), .A2(new_n257), .ZN(new_n258));
  OR2_X1    g057(.A1(new_n223), .A2(KEYINPUT26), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n219), .A2(new_n220), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n223), .A2(KEYINPUT26), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(KEYINPUT27), .B(G183gat), .Z(new_n263));
  OAI21_X1  g062(.A(KEYINPUT28), .B1(new_n263), .B2(G190gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265));
  OR3_X1    g064(.A1(new_n207), .A2(KEYINPUT67), .A3(KEYINPUT27), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT27), .B1(new_n207), .B2(KEYINPUT67), .ZN(new_n267));
  NOR2_X1   g066(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n262), .A2(new_n264), .A3(new_n265), .A4(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n239), .A2(new_n258), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n258), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n237), .B1(new_n231), .B2(new_n232), .ZN(new_n273));
  INV_X1    g072(.A(new_n270), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n204), .B1(new_n271), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT34), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI211_X1 g077(.A(KEYINPUT34), .B(new_n204), .C1(new_n271), .C2(new_n275), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XOR2_X1   g079(.A(G15gat), .B(G43gat), .Z(new_n281));
  XNOR2_X1  g080(.A(G71gat), .B(G99gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n271), .A2(new_n204), .A3(new_n275), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT33), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n280), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n285), .A2(KEYINPUT32), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n287), .B1(new_n278), .B2(new_n279), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n289), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n291), .B1(new_n289), .B2(new_n292), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT36), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n289), .A2(new_n292), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n290), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n289), .A2(new_n291), .A3(new_n292), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT36), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G225gat), .A2(G233gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT2), .ZN(new_n306));
  INV_X1    g105(.A(G141gat), .ZN(new_n307));
  INV_X1    g106(.A(G148gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G141gat), .A2(G148gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n306), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  OR3_X1    g110(.A1(KEYINPUT74), .A2(G155gat), .A3(G162gat), .ZN(new_n312));
  INV_X1    g111(.A(G155gat), .ZN(new_n313));
  INV_X1    g112(.A(G162gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT74), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n311), .A2(new_n305), .A3(new_n312), .A4(new_n316), .ZN(new_n317));
  AND2_X1   g116(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n305), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  XOR2_X1   g118(.A(G141gat), .B(G148gat), .Z(new_n320));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n258), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n317), .A2(new_n247), .A3(new_n323), .A4(new_n257), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n304), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT5), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT76), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n304), .ZN(new_n330));
  AND4_X1   g129(.A1(new_n257), .A2(new_n317), .A3(new_n247), .A4(new_n323), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n323), .A2(new_n317), .B1(new_n247), .B2(new_n257), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT76), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT5), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n324), .A2(KEYINPUT3), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT3), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n317), .A2(new_n323), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n258), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n324), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n340), .A2(new_n272), .A3(KEYINPUT4), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT4), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n339), .A2(new_n341), .A3(new_n304), .A4(new_n343), .ZN(new_n344));
  AND3_X1   g143(.A1(new_n329), .A2(new_n335), .A3(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT77), .B1(new_n344), .B2(KEYINPUT5), .ZN(new_n346));
  OR2_X1    g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G1gat), .B(G29gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT0), .ZN(new_n349));
  XNOR2_X1  g148(.A(G57gat), .B(G85gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n329), .A2(new_n335), .A3(new_n352), .A4(new_n344), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n347), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT6), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n353), .B1(new_n345), .B2(new_n346), .ZN(new_n356));
  INV_X1    g155(.A(new_n351), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n354), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n347), .A2(KEYINPUT6), .A3(new_n351), .A4(new_n353), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT71), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n239), .A2(new_n362), .A3(new_n270), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT71), .B1(new_n273), .B2(new_n274), .ZN(new_n364));
  INV_X1    g163(.A(G226gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n365), .A2(new_n203), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(KEYINPUT29), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n363), .A2(new_n364), .A3(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G197gat), .B(G204gat), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT22), .ZN(new_n370));
  INV_X1    g169(.A(G211gat), .ZN(new_n371));
  INV_X1    g170(.A(G218gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G211gat), .B(G218gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT70), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n375), .A2(new_n369), .A3(new_n373), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n374), .A2(KEYINPUT70), .A3(new_n376), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n239), .A2(new_n270), .A3(new_n366), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n368), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT72), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n368), .A2(KEYINPUT72), .A3(new_n382), .A4(new_n383), .ZN(new_n387));
  INV_X1    g186(.A(new_n382), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n362), .B1(new_n239), .B2(new_n270), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n273), .A2(KEYINPUT71), .A3(new_n274), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n366), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n239), .A2(new_n270), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n367), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n386), .A2(new_n387), .B1(new_n388), .B2(new_n394), .ZN(new_n395));
  XOR2_X1   g194(.A(G8gat), .B(G36gat), .Z(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(KEYINPUT73), .ZN(new_n397));
  XNOR2_X1  g196(.A(G64gat), .B(G92gat), .ZN(new_n398));
  XOR2_X1   g197(.A(new_n397), .B(new_n398), .Z(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n395), .A2(KEYINPUT30), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n395), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n399), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n387), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n394), .A2(new_n388), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n400), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT30), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n361), .A2(new_n401), .A3(new_n403), .A4(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT78), .ZN(new_n410));
  NAND2_X1  g209(.A1(G228gat), .A2(G233gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n377), .A2(new_n379), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT29), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n340), .B1(new_n414), .B2(new_n337), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n413), .A2(new_n338), .B1(new_n380), .B2(new_n381), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n411), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OR2_X1    g216(.A1(new_n416), .A2(new_n411), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n380), .A2(new_n413), .A3(new_n381), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n340), .B1(new_n419), .B2(new_n337), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n417), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n410), .B1(new_n421), .B2(G22gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(G78gat), .B(G106gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT31), .B(G50gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT79), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT79), .ZN(new_n428));
  INV_X1    g227(.A(G22gat), .ZN(new_n429));
  OR3_X1    g228(.A1(new_n420), .A2(new_n411), .A3(new_n416), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n429), .B1(new_n430), .B2(new_n417), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n428), .B(new_n425), .C1(new_n431), .C2(new_n410), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n421), .A2(G22gat), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(new_n431), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n427), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n434), .B1(new_n427), .B2(new_n432), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n409), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n303), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT84), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n351), .B(KEYINPUT80), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n353), .B(new_n442), .C1(new_n345), .C2(new_n346), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n358), .A2(new_n355), .A3(new_n443), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n444), .A2(new_n360), .A3(new_n406), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT82), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n368), .A2(new_n388), .A3(new_n383), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT37), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n388), .B1(new_n391), .B2(new_n393), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n393), .ZN(new_n451));
  INV_X1    g250(.A(new_n366), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n452), .B1(new_n363), .B2(new_n364), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n382), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n454), .A2(KEYINPUT82), .A3(KEYINPUT37), .A4(new_n447), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT37), .B1(new_n394), .B2(new_n388), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n400), .B1(new_n404), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT38), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n456), .A2(new_n458), .A3(KEYINPUT83), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n460), .ZN(new_n461));
  AOI211_X1 g260(.A(KEYINPUT38), .B(new_n400), .C1(new_n404), .C2(new_n457), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT83), .B1(new_n462), .B2(new_n456), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n440), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT83), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n458), .A2(new_n459), .ZN(new_n466));
  INV_X1    g265(.A(new_n456), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n468), .A2(KEYINPUT84), .A3(new_n460), .A4(new_n445), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n402), .A2(KEYINPUT37), .ZN(new_n470));
  INV_X1    g269(.A(new_n458), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT38), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n464), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n341), .A2(new_n343), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n304), .B1(new_n474), .B2(new_n339), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT39), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n331), .A2(new_n332), .A3(new_n330), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI211_X1 g277(.A(new_n442), .B(new_n478), .C1(new_n476), .C2(new_n475), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT40), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n443), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT81), .ZN(new_n482));
  OR3_X1    g281(.A1(new_n479), .A2(new_n482), .A3(KEYINPUT40), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n482), .B1(new_n479), .B2(KEYINPUT40), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n403), .A2(new_n408), .A3(new_n401), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n437), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n439), .B1(new_n473), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n436), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n427), .A2(new_n432), .A3(new_n434), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT35), .B1(new_n444), .B2(new_n360), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n295), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT85), .B1(new_n493), .B2(new_n486), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n491), .A2(new_n295), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT35), .B1(new_n495), .B2(new_n409), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n300), .A2(new_n437), .ZN(new_n497));
  INV_X1    g296(.A(new_n486), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT85), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n497), .A2(new_n498), .A3(new_n499), .A4(new_n492), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n494), .A2(new_n496), .A3(new_n500), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n488), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n503));
  NAND2_X1  g302(.A1(G229gat), .A2(G233gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT15), .ZN(new_n507));
  INV_X1    g306(.A(G50gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(G43gat), .ZN(new_n509));
  INV_X1    g308(.A(G43gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(G50gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OR3_X1    g311(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n507), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n509), .A2(new_n511), .A3(KEYINPUT15), .ZN(new_n516));
  NAND2_X1  g315(.A1(G29gat), .A2(G36gat), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n515), .A2(KEYINPUT88), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT88), .ZN(new_n519));
  XNOR2_X1  g318(.A(G43gat), .B(G50gat), .ZN(new_n520));
  INV_X1    g319(.A(new_n514), .ZN(new_n521));
  NOR3_X1   g320(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n522));
  OAI22_X1  g321(.A1(new_n520), .A2(KEYINPUT15), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n516), .A2(new_n517), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n519), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n518), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n514), .A2(KEYINPUT87), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT87), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n528), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n527), .A2(new_n513), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n516), .B1(new_n530), .B2(new_n517), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G15gat), .B(G22gat), .ZN(new_n534));
  INV_X1    g333(.A(G1gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT16), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT89), .B1(new_n534), .B2(G1gat), .ZN(new_n539));
  OAI21_X1  g338(.A(G8gat), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n534), .A2(G1gat), .ZN(new_n541));
  INV_X1    g340(.A(G8gat), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n541), .A2(new_n537), .A3(KEYINPUT89), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n533), .A2(new_n544), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n526), .A2(new_n532), .B1(new_n540), .B2(new_n543), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n506), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT93), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT93), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n549), .B(new_n506), .C1(new_n545), .C2(new_n546), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(KEYINPUT91), .A2(KEYINPUT18), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n533), .A2(KEYINPUT17), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n526), .A2(new_n554), .A3(new_n532), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT90), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n540), .A2(new_n543), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(new_n540), .B2(new_n543), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n546), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n552), .B1(new_n561), .B2(new_n504), .ZN(new_n562));
  INV_X1    g361(.A(new_n546), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n554), .B1(new_n526), .B2(new_n532), .ZN(new_n564));
  AOI211_X1 g363(.A(KEYINPUT17), .B(new_n531), .C1(new_n518), .C2(new_n525), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n560), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AND4_X1   g365(.A1(new_n563), .A2(new_n566), .A3(new_n504), .A4(new_n552), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n551), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G113gat), .B(G141gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G169gat), .B(G197gat), .Z(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT12), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n568), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n551), .B(new_n574), .C1(new_n562), .C2(new_n567), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n579), .A2(KEYINPUT94), .ZN(new_n580));
  XOR2_X1   g379(.A(G71gat), .B(G78gat), .Z(new_n581));
  AOI21_X1  g380(.A(new_n580), .B1(new_n581), .B2(KEYINPUT95), .ZN(new_n582));
  XNOR2_X1  g381(.A(G71gat), .B(G78gat), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT95), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n579), .A2(KEYINPUT94), .ZN(new_n586));
  NAND2_X1  g385(.A1(G57gat), .A2(G64gat), .ZN(new_n587));
  OR2_X1    g386(.A1(G57gat), .A2(G64gat), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n582), .A2(new_n585), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n584), .B(new_n583), .C1(new_n591), .C2(new_n580), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n593), .A2(KEYINPUT21), .ZN(new_n594));
  NAND2_X1  g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(new_n243), .ZN(new_n597));
  XNOR2_X1  g396(.A(G183gat), .B(G211gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n544), .B1(new_n593), .B2(KEYINPUT21), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n600), .B(KEYINPUT96), .Z(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(new_n313), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n601), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n599), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G190gat), .B(G218gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT100), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT41), .ZN(new_n608));
  NAND2_X1  g407(.A1(G232gat), .A2(G233gat), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G85gat), .A2(G92gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT97), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT97), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n613), .A2(G85gat), .A3(G92gat), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n612), .A2(new_n614), .A3(KEYINPUT7), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT7), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n611), .A2(KEYINPUT97), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(G85gat), .ZN(new_n618));
  INV_X1    g417(.A(G92gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G99gat), .A2(G106gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT8), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n617), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n615), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(G99gat), .ZN(new_n625));
  INV_X1    g424(.A(G106gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n621), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT98), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT98), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n627), .A2(new_n630), .A3(new_n621), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n624), .A2(new_n632), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n629), .B(new_n631), .C1(new_n615), .C2(new_n623), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n633), .A2(new_n634), .A3(KEYINPUT99), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT99), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n624), .A2(new_n636), .A3(new_n632), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n610), .B1(new_n638), .B2(new_n533), .ZN(new_n639));
  INV_X1    g438(.A(new_n556), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n639), .B1(new_n640), .B2(new_n638), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n606), .A2(KEYINPUT100), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(G134gat), .B(G162gat), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n609), .A2(new_n608), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n641), .A2(new_n642), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n643), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n646), .B1(new_n643), .B2(new_n647), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(G230gat), .A2(G233gat), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n652), .B(KEYINPUT101), .Z(new_n653));
  NAND4_X1  g452(.A1(new_n635), .A2(new_n592), .A3(new_n590), .A4(new_n637), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT10), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n593), .A2(new_n633), .A3(new_n634), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n638), .A2(KEYINPUT10), .A3(new_n593), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n654), .A2(new_n656), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n659), .B1(new_n653), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G120gat), .B(G148gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(G176gat), .B(G204gat), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n662), .B(new_n663), .Z(new_n664));
  OR2_X1    g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n661), .A2(new_n664), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n605), .A2(new_n651), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n502), .A2(new_n578), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT102), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n502), .A2(new_n673), .A3(new_n578), .A4(new_n670), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n361), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g477(.A(KEYINPUT16), .B(G8gat), .Z(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  AOI211_X1 g479(.A(new_n498), .B(new_n680), .C1(new_n672), .C2(new_n674), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n681), .A2(KEYINPUT42), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n542), .B1(new_n675), .B2(new_n486), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT42), .B1(new_n683), .B2(new_n681), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(G1325gat));
  INV_X1    g484(.A(G15gat), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n675), .A2(new_n686), .A3(new_n295), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n303), .B1(new_n672), .B2(new_n674), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(new_n688), .B2(new_n686), .ZN(G1326gat));
  NAND2_X1  g488(.A1(new_n675), .A2(new_n437), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT103), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT103), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n675), .A2(new_n692), .A3(new_n437), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT43), .B(G22gat), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n694), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n692), .B1(new_n675), .B2(new_n437), .ZN(new_n697));
  AOI211_X1 g496(.A(KEYINPUT103), .B(new_n491), .C1(new_n672), .C2(new_n674), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n695), .A2(new_n699), .ZN(G1327gat));
  OAI21_X1  g499(.A(new_n650), .B1(new_n488), .B2(new_n501), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n578), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n605), .A2(new_n704), .A3(new_n667), .ZN(new_n705));
  OAI211_X1 g504(.A(KEYINPUT44), .B(new_n650), .C1(new_n488), .C2(new_n501), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n703), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G29gat), .B1(new_n707), .B2(new_n361), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n502), .A2(new_n650), .A3(new_n705), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n361), .A2(G29gat), .ZN(new_n711));
  OR3_X1    g510(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n709), .B2(new_n711), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n708), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT104), .ZN(G1328gat));
  OR2_X1    g514(.A1(new_n651), .A2(G36gat), .ZN(new_n716));
  NOR4_X1   g515(.A1(new_n716), .A2(new_n498), .A3(new_n605), .A4(new_n667), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n502), .A2(new_n578), .A3(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(G36gat), .B1(new_n707), .B2(new_n498), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1329gat));
  INV_X1    g523(.A(new_n709), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n725), .A2(new_n510), .A3(new_n295), .ZN(new_n726));
  INV_X1    g525(.A(new_n303), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n703), .A2(new_n727), .A3(new_n705), .A4(new_n706), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G43gat), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n728), .A2(new_n729), .ZN(new_n732));
  OAI211_X1 g531(.A(KEYINPUT47), .B(new_n726), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n728), .A2(G43gat), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n726), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(KEYINPUT47), .B2(new_n735), .ZN(G1330gat));
  NAND3_X1  g535(.A1(new_n725), .A2(new_n508), .A3(new_n437), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT48), .B1(new_n737), .B2(KEYINPUT107), .ZN(new_n738));
  OAI21_X1  g537(.A(G50gat), .B1(new_n707), .B2(new_n491), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n737), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n738), .B(new_n740), .ZN(G1331gat));
  INV_X1    g540(.A(new_n605), .ZN(new_n742));
  NOR4_X1   g541(.A1(new_n742), .A2(new_n578), .A3(new_n650), .A4(new_n668), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n502), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n676), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT108), .B(G57gat), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1332gat));
  INV_X1    g546(.A(KEYINPUT49), .ZN(new_n748));
  INV_X1    g547(.A(G64gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n486), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT109), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n744), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n748), .A2(new_n749), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1333gat));
  NAND4_X1  g553(.A1(new_n502), .A2(G71gat), .A3(new_n727), .A4(new_n743), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n744), .A2(new_n295), .ZN(new_n758));
  INV_X1    g557(.A(G71gat), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT50), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n757), .A2(new_n763), .A3(new_n760), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(G1334gat));
  NAND2_X1  g564(.A1(new_n744), .A2(new_n437), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g566(.A1(new_n605), .A2(new_n578), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n668), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n703), .A2(new_n706), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT111), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n703), .A2(new_n773), .A3(new_n706), .A4(new_n770), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n772), .A2(new_n676), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n772), .A2(KEYINPUT112), .A3(new_n676), .A4(new_n774), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(G85gat), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n502), .A2(new_n780), .A3(new_n650), .A4(new_n768), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT51), .B1(new_n701), .B2(new_n769), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(new_n667), .A3(new_n782), .ZN(new_n783));
  OR3_X1    g582(.A1(new_n783), .A2(G85gat), .A3(new_n361), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n779), .A2(new_n784), .ZN(G1336gat));
  OAI21_X1  g584(.A(G92gat), .B1(new_n771), .B2(new_n498), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n486), .A2(new_n619), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n786), .B(new_n787), .C1(new_n783), .C2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n783), .A2(new_n788), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n772), .A2(new_n486), .A3(new_n774), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n791), .B2(G92gat), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n789), .B1(new_n792), .B2(new_n787), .ZN(G1337gat));
  NAND4_X1  g592(.A1(new_n772), .A2(G99gat), .A3(new_n727), .A4(new_n774), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n625), .B1(new_n783), .B2(new_n300), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT113), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n794), .A2(new_n798), .A3(new_n795), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1338gat));
  XOR2_X1   g599(.A(KEYINPUT114), .B(G106gat), .Z(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(new_n771), .B2(new_n491), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n437), .A2(new_n626), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n802), .B(new_n803), .C1(new_n783), .C2(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n783), .A2(new_n804), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n772), .A2(new_n437), .A3(new_n774), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n806), .B1(new_n807), .B2(new_n801), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n805), .B1(new_n808), .B2(new_n803), .ZN(G1339gat));
  NAND3_X1  g608(.A1(new_n657), .A2(new_n653), .A3(new_n658), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n657), .A2(new_n658), .ZN(new_n812));
  INV_X1    g611(.A(new_n653), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n657), .A2(new_n658), .A3(new_n815), .A4(new_n653), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n811), .A2(new_n814), .A3(KEYINPUT54), .A4(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n664), .B1(new_n659), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT55), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n817), .A2(KEYINPUT55), .A3(new_n819), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n666), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n820), .B1(new_n822), .B2(KEYINPUT116), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n821), .A2(new_n824), .A3(new_n666), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n823), .A2(new_n578), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n827), .B1(new_n561), .B2(new_n504), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n504), .B1(new_n566), .B2(new_n563), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT117), .ZN(new_n830));
  OR3_X1    g629(.A1(new_n545), .A2(new_n546), .A3(new_n506), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n573), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT118), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n831), .B1(new_n829), .B2(KEYINPUT117), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n561), .A2(new_n827), .A3(new_n504), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n835), .B(new_n573), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n834), .A2(new_n667), .A3(new_n577), .A4(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n650), .B1(new_n826), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n577), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n835), .B1(new_n832), .B2(new_n573), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AND4_X1   g642(.A1(new_n650), .A2(new_n823), .A3(new_n843), .A4(new_n825), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n742), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n670), .A2(new_n704), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n437), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AND4_X1   g646(.A1(new_n676), .A2(new_n847), .A3(new_n498), .A4(new_n295), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n578), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n667), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g651(.A1(new_n848), .A2(new_n605), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT119), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n240), .A2(new_n241), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n854), .B(new_n855), .ZN(G1342gat));
  INV_X1    g655(.A(KEYINPUT56), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n650), .B1(new_n857), .B2(new_n244), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n858), .A2(new_n361), .A3(new_n300), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n847), .A2(new_n498), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n857), .A2(new_n244), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n860), .B(new_n861), .ZN(G1343gat));
  NOR3_X1   g661(.A1(new_n727), .A2(new_n361), .A3(new_n486), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n845), .A2(new_n846), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT57), .B1(new_n864), .B2(new_n437), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n491), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n823), .A2(new_n843), .A3(new_n650), .A4(new_n825), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n820), .B1(new_n576), .B2(new_n577), .ZN(new_n871));
  INV_X1    g670(.A(new_n822), .ZN(new_n872));
  AOI22_X1  g671(.A1(new_n843), .A2(new_n667), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n870), .B1(new_n873), .B2(new_n650), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n874), .A2(new_n742), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n669), .A2(new_n578), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n869), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n865), .B2(new_n866), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n578), .B(new_n863), .C1(new_n867), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(G141gat), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n864), .A2(new_n437), .A3(new_n863), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n578), .A2(new_n307), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT121), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(KEYINPUT58), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT58), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n880), .A2(new_n888), .A3(new_n885), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(G1344gat));
  OAI21_X1  g689(.A(new_n863), .B1(new_n867), .B2(new_n878), .ZN(new_n891));
  OAI21_X1  g690(.A(G148gat), .B1(new_n891), .B2(new_n668), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n882), .A2(new_n308), .A3(new_n667), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n871), .A2(new_n872), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n650), .B1(new_n897), .B2(new_n839), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n896), .B1(new_n844), .B2(new_n898), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n870), .B(KEYINPUT122), .C1(new_n873), .C2(new_n650), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(new_n742), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n491), .B1(new_n901), .B2(new_n846), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT123), .B1(new_n902), .B2(KEYINPUT57), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n605), .B1(new_n874), .B2(new_n896), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n876), .B1(new_n905), .B2(new_n900), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n904), .B(new_n868), .C1(new_n906), .C2(new_n491), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n864), .A2(new_n869), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n903), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n909), .A2(new_n667), .A3(new_n863), .ZN(new_n910));
  NAND2_X1  g709(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n894), .B(new_n895), .C1(new_n910), .C2(new_n911), .ZN(G1345gat));
  OAI21_X1  g711(.A(G155gat), .B1(new_n891), .B2(new_n742), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n882), .A2(new_n313), .A3(new_n605), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1346gat));
  OAI21_X1  g714(.A(G162gat), .B1(new_n891), .B2(new_n651), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n882), .A2(new_n314), .A3(new_n650), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1347gat));
  AOI21_X1  g717(.A(new_n676), .B1(new_n845), .B2(new_n846), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n495), .A2(new_n498), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n578), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n486), .A2(new_n361), .ZN(new_n924));
  XOR2_X1   g723(.A(new_n924), .B(KEYINPUT124), .Z(new_n925));
  NOR2_X1   g724(.A1(new_n925), .A2(new_n300), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n847), .A2(new_n926), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n927), .A2(KEYINPUT125), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(KEYINPUT125), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n704), .A2(new_n221), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n923), .B1(new_n930), .B2(new_n931), .ZN(G1348gat));
  NAND2_X1  g731(.A1(new_n928), .A2(new_n929), .ZN(new_n933));
  OAI21_X1  g732(.A(G176gat), .B1(new_n933), .B2(new_n668), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n922), .A2(new_n222), .A3(new_n667), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1349gat));
  OAI21_X1  g735(.A(G183gat), .B1(new_n933), .B2(new_n742), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n921), .A2(new_n263), .A3(new_n742), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT60), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT60), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n937), .A2(new_n942), .A3(new_n939), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1350gat));
  NAND3_X1  g743(.A1(new_n922), .A2(new_n209), .A3(new_n650), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n650), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n946), .B1(new_n947), .B2(G190gat), .ZN(new_n948));
  AOI211_X1 g747(.A(KEYINPUT61), .B(new_n209), .C1(new_n930), .C2(new_n650), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(G1351gat));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n925), .A2(new_n727), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n909), .A2(new_n578), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G197gat), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n919), .A2(new_n437), .A3(new_n486), .A4(new_n303), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n955), .A2(G197gat), .A3(new_n704), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n951), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  AOI211_X1 g757(.A(KEYINPUT126), .B(new_n956), .C1(new_n953), .C2(G197gat), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n958), .A2(new_n959), .ZN(G1352gat));
  NAND2_X1  g759(.A1(new_n909), .A2(new_n952), .ZN(new_n961));
  OAI21_X1  g760(.A(G204gat), .B1(new_n961), .B2(new_n668), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n955), .A2(G204gat), .A3(new_n668), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT62), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n964), .ZN(G1353gat));
  OAI21_X1  g764(.A(G211gat), .B1(new_n961), .B2(new_n742), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(KEYINPUT63), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT63), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n968), .B(G211gat), .C1(new_n961), .C2(new_n742), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n955), .A2(G211gat), .A3(new_n742), .ZN(new_n970));
  XOR2_X1   g769(.A(new_n970), .B(KEYINPUT127), .Z(new_n971));
  NAND3_X1  g770(.A1(new_n967), .A2(new_n969), .A3(new_n971), .ZN(G1354gat));
  OAI21_X1  g771(.A(G218gat), .B1(new_n961), .B2(new_n651), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n650), .A2(new_n372), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n973), .B1(new_n955), .B2(new_n974), .ZN(G1355gat));
endmodule


