//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  XNOR2_X1  g012(.A(KEYINPUT67), .B(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XNOR2_X1  g015(.A(KEYINPUT68), .B(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  AND2_X1   g017(.A1(G2072), .A2(G2078), .ZN(new_n443));
  NAND3_X1  g018(.A1(new_n443), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n463), .A2(G2105), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n466), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n469), .B1(new_n464), .B2(new_n465), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT69), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(G113), .A3(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g050(.A(G2105), .B1(new_n470), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n468), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n466), .A2(G136), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT70), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G112), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n465), .ZN(new_n484));
  NOR2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(G2105), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n483), .B1(new_n488), .B2(G124), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n480), .A2(new_n489), .ZN(G162));
  NAND2_X1  g065(.A1(KEYINPUT4), .A2(G138), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(new_n464), .B2(new_n465), .ZN(new_n492));
  AND2_X1   g067(.A1(G102), .A2(G2104), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n487), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n464), .B2(new_n465), .ZN(new_n496));
  AND2_X1   g071(.A1(G114), .A2(G2104), .ZN(new_n497));
  OAI21_X1  g072(.A(G2105), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(G138), .B(new_n487), .C1(new_n484), .C2(new_n485), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n494), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  NAND2_X1  g078(.A1(G75), .A2(G543), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G62), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n504), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G651), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n513), .A2(new_n507), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G88), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(G50), .A3(G543), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n517), .A2(KEYINPUT71), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(KEYINPUT71), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n510), .B(new_n515), .C1(new_n518), .C2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  XOR2_X1   g098(.A(KEYINPUT72), .B(G51), .Z(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n523), .A2(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n516), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n507), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT73), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n528), .B(new_n532), .C1(new_n507), .C2(new_n529), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(G168));
  XNOR2_X1  g109(.A(KEYINPUT5), .B(G543), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n535), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G651), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n516), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n512), .A2(new_n511), .B1(new_n505), .B2(new_n506), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n539), .A2(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(KEYINPUT74), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT74), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n546), .B1(new_n538), .B2(new_n543), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n545), .A2(new_n547), .ZN(G171));
  AOI22_X1  g123(.A1(new_n535), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n537), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n539), .A2(new_n551), .B1(new_n541), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND2_X1  g134(.A1(new_n523), .A2(G53), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n507), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(G651), .A2(new_n564), .B1(new_n514), .B2(G91), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  INV_X1    g142(.A(G168), .ZN(G286));
  OR2_X1    g143(.A1(new_n535), .A2(G74), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n569), .A2(G651), .B1(new_n523), .B2(G49), .ZN(new_n570));
  AND3_X1   g145(.A1(new_n514), .A2(KEYINPUT75), .A3(G87), .ZN(new_n571));
  AOI21_X1  g146(.A(KEYINPUT75), .B1(new_n514), .B2(G87), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(G288));
  OAI211_X1 g148(.A(G48), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n574));
  INV_X1    g149(.A(G86), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n541), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n535), .B2(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n577), .B1(new_n580), .B2(new_n537), .ZN(new_n581));
  OAI21_X1  g156(.A(G61), .B1(new_n505), .B2(new_n506), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(new_n578), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n583), .A2(KEYINPUT76), .A3(G651), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n576), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n535), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n537), .ZN(new_n588));
  INV_X1    g163(.A(G47), .ZN(new_n589));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n539), .A2(new_n589), .B1(new_n541), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G290));
  INV_X1    g168(.A(G54), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n594), .B1(new_n539), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n523), .A2(KEYINPUT78), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n507), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n596), .A2(new_n597), .B1(G651), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT77), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n514), .A2(new_n602), .A3(G92), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT77), .B1(new_n541), .B2(new_n605), .ZN(new_n606));
  AND3_X1   g181(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n604), .B1(new_n603), .B2(new_n606), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n601), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g186(.A(new_n610), .B1(G868), .B2(G171), .ZN(G321));
  NOR2_X1   g187(.A1(G299), .A2(G868), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g189(.A(new_n613), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g190(.A(new_n601), .ZN(new_n616));
  INV_X1    g191(.A(new_n608), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G860), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT79), .ZN(G148));
  NAND2_X1  g197(.A1(new_n619), .A2(new_n620), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g201(.A(new_n486), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(new_n467), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2100), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n488), .A2(G123), .B1(G135), .B2(new_n466), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(G111), .ZN(new_n635));
  AOI22_X1  g210(.A1(new_n634), .A2(KEYINPUT81), .B1(new_n635), .B2(G2105), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(KEYINPUT81), .B2(new_n634), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(KEYINPUT82), .B(G2096), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n632), .A2(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT83), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2427), .B(G2430), .Z(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(KEYINPUT14), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n648), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(new_n656), .A3(G14), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT84), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G401));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT85), .ZN(new_n661));
  NOR2_X1   g236(.A1(G2072), .A2(G2078), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n443), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2084), .B(G2090), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n661), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT18), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n661), .A2(new_n663), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n663), .B(KEYINPUT17), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n667), .B(new_n664), .C1(new_n661), .C2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n664), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n668), .A2(new_n661), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n666), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2096), .B(G2100), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT20), .ZN(new_n682));
  INV_X1    g257(.A(new_n677), .ZN(new_n683));
  INV_X1    g258(.A(new_n680), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n678), .A2(new_n679), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n682), .B(new_n686), .C1(new_n683), .C2(new_n685), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT87), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT88), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n689), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  MUX2_X1   g271(.A(G23), .B(G288), .S(G16), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT33), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1976), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G6), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n585), .B2(new_n700), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT32), .B(G1981), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  INV_X1    g280(.A(G22), .ZN(new_n706));
  OR3_X1    g281(.A1(new_n706), .A2(KEYINPUT91), .A3(G16), .ZN(new_n707));
  OAI21_X1  g282(.A(KEYINPUT91), .B1(new_n706), .B2(G16), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n707), .B(new_n708), .C1(G166), .C2(new_n700), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n709), .A2(G1971), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(G1971), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n699), .A2(new_n704), .A3(new_n705), .A4(new_n712), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n713), .A2(KEYINPUT34), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(KEYINPUT34), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G25), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT89), .Z(new_n718));
  OR2_X1    g293(.A1(G95), .A2(G2105), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n719), .B(G2104), .C1(G107), .C2(new_n487), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT90), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n488), .A2(G119), .B1(G131), .B2(new_n466), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n718), .B1(new_n723), .B2(G29), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT35), .B(G1991), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n724), .B(new_n725), .Z(new_n726));
  NOR2_X1   g301(.A1(new_n592), .A2(new_n700), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n700), .B2(G24), .ZN(new_n728));
  INV_X1    g303(.A(G1986), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  NOR3_X1   g306(.A1(new_n726), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n714), .A2(new_n715), .A3(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT92), .B(KEYINPUT36), .Z(new_n734));
  AND2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n716), .A2(G26), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT28), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n488), .A2(G128), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n466), .A2(G140), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n487), .A2(G116), .ZN(new_n740));
  OAI21_X1  g315(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n738), .B(new_n739), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT94), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n737), .B1(new_n743), .B2(G29), .ZN(new_n744));
  INV_X1    g319(.A(G2067), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n716), .A2(G27), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G164), .B2(new_n716), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G2078), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT95), .B(KEYINPUT24), .ZN(new_n750));
  INV_X1    g325(.A(G34), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n716), .B1(new_n750), .B2(new_n751), .ZN(new_n753));
  OAI22_X1  g328(.A1(G160), .A2(new_n716), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G2084), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n716), .A2(G33), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n627), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n757), .A2(new_n487), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n487), .A2(G103), .A3(G2104), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT25), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n466), .A2(G139), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n756), .B1(new_n763), .B2(new_n716), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G2072), .ZN(new_n765));
  NOR4_X1   g340(.A1(new_n746), .A2(new_n749), .A3(new_n755), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n716), .A2(G35), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G162), .B2(new_n716), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT29), .B(G2090), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G4), .A2(G16), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n619), .B2(G16), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n772), .A2(G1348), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT30), .B(G28), .ZN(new_n774));
  OR2_X1    g349(.A1(KEYINPUT31), .A2(G11), .ZN(new_n775));
  NAND2_X1  g350(.A1(KEYINPUT31), .A2(G11), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n774), .A2(new_n716), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n638), .B2(new_n716), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT100), .Z(new_n779));
  NOR3_X1   g354(.A1(new_n770), .A2(new_n773), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G5), .A2(G16), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G171), .B2(G16), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1961), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G1348), .B2(new_n772), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n700), .A2(G20), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT23), .Z(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G299), .B2(G16), .ZN(new_n787));
  INV_X1    g362(.A(G1956), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G16), .A2(G19), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n554), .B2(G16), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT93), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n792), .A2(G1341), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n792), .A2(G1341), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n789), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n766), .A2(new_n780), .A3(new_n784), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n716), .A2(G32), .ZN(new_n797));
  NAND3_X1  g372(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT26), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n467), .A2(G105), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT97), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n627), .A2(G2105), .ZN(new_n803));
  INV_X1    g378(.A(G129), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n488), .A2(KEYINPUT97), .A3(G129), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n801), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n466), .A2(G141), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT96), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT98), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n807), .A2(new_n809), .A3(KEYINPUT98), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n797), .B1(new_n815), .B2(new_n716), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT27), .B(G1996), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  AND3_X1   g393(.A1(G168), .A2(KEYINPUT99), .A3(G16), .ZN(new_n819));
  AOI21_X1  g394(.A(KEYINPUT99), .B1(G168), .B2(G16), .ZN(new_n820));
  OAI22_X1  g395(.A1(new_n819), .A2(new_n820), .B1(G16), .B2(G21), .ZN(new_n821));
  INV_X1    g396(.A(G1966), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n796), .A2(new_n818), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n733), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n735), .A2(new_n826), .ZN(G311));
  OR2_X1    g402(.A1(new_n735), .A2(new_n826), .ZN(G150));
  NOR2_X1   g403(.A1(new_n609), .A2(new_n620), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT38), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n535), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(new_n537), .ZN(new_n832));
  INV_X1    g407(.A(G55), .ZN(new_n833));
  INV_X1    g408(.A(G93), .ZN(new_n834));
  OAI22_X1  g409(.A1(new_n539), .A2(new_n833), .B1(new_n541), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n554), .B(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n830), .B(new_n837), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n839));
  INV_X1    g414(.A(G860), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n836), .A2(new_n840), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT37), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(G145));
  NAND3_X1  g420(.A1(new_n812), .A2(G164), .A3(new_n813), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n743), .ZN(new_n848));
  AOI21_X1  g423(.A(G164), .B1(new_n812), .B2(new_n813), .ZN(new_n849));
  NOR3_X1   g424(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n814), .A2(new_n502), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n743), .B1(new_n851), .B2(new_n846), .ZN(new_n852));
  OAI22_X1  g427(.A1(new_n850), .A2(new_n852), .B1(new_n758), .B2(new_n762), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n488), .A2(G130), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n466), .A2(G142), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n487), .A2(G118), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n854), .B(new_n855), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n723), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n630), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n848), .B1(new_n847), .B2(new_n849), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n851), .A2(new_n743), .A3(new_n846), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n861), .A2(new_n763), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n853), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(KEYINPUT101), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n853), .A2(new_n863), .ZN(new_n866));
  INV_X1    g441(.A(new_n860), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n866), .A2(KEYINPUT101), .A3(new_n867), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n638), .B(G160), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(G162), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(G37), .ZN(new_n875));
  INV_X1    g450(.A(new_n873), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n864), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n860), .B1(new_n853), .B2(new_n863), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(KEYINPUT40), .B1(new_n874), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n876), .B1(new_n869), .B2(new_n870), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT40), .ZN(new_n883));
  NOR3_X1   g458(.A1(new_n882), .A2(new_n883), .A3(new_n879), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n881), .A2(new_n884), .ZN(G395));
  NAND2_X1  g460(.A1(new_n619), .A2(G299), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT9), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n560), .B(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n565), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n609), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n887), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n891), .A2(new_n609), .A3(KEYINPUT103), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n886), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n894), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n895), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(KEYINPUT104), .A3(new_n894), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(new_n554), .B(new_n836), .Z(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT102), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(new_n623), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT105), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n886), .A2(new_n892), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n904), .A2(KEYINPUT105), .A3(new_n907), .ZN(new_n913));
  XNOR2_X1  g488(.A(G288), .B(new_n592), .ZN(new_n914));
  XNOR2_X1  g489(.A(G303), .B(new_n585), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n915), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT107), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n919), .A2(new_n924), .A3(new_n921), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n923), .A2(new_n925), .A3(new_n927), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n912), .A2(new_n913), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n931), .B1(new_n912), .B2(new_n913), .ZN(new_n933));
  OAI21_X1  g508(.A(G868), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(G868), .B2(new_n836), .ZN(G295));
  OAI21_X1  g510(.A(new_n934), .B1(G868), .B2(new_n836), .ZN(G331));
  INV_X1    g511(.A(KEYINPUT109), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n531), .A2(new_n545), .A3(new_n533), .A4(new_n547), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n533), .A2(new_n531), .B1(new_n545), .B2(new_n547), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n837), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n942));
  NAND2_X1  g517(.A1(G168), .A2(G171), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n905), .A2(new_n943), .A3(new_n938), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n905), .A2(new_n943), .A3(KEYINPUT108), .A4(new_n938), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(new_n902), .B2(new_n903), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n941), .A2(new_n909), .A3(new_n944), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n937), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n903), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT104), .B1(new_n899), .B2(new_n894), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n952), .A2(new_n953), .A3(new_n895), .ZN(new_n954));
  OAI211_X1 g529(.A(KEYINPUT109), .B(new_n949), .C1(new_n954), .C2(new_n947), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n917), .A2(KEYINPUT110), .A3(new_n918), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n957));
  INV_X1    g532(.A(new_n918), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n957), .B1(new_n958), .B2(new_n916), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n951), .A2(new_n955), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n948), .A2(new_n950), .ZN(new_n962));
  AOI21_X1  g537(.A(G37), .B1(new_n962), .B2(new_n919), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT43), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n910), .B1(new_n945), .B2(new_n946), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n897), .A2(KEYINPUT41), .A3(new_n886), .A4(new_n898), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n909), .A2(new_n894), .ZN(new_n967));
  AOI22_X1  g542(.A1(new_n966), .A2(new_n967), .B1(new_n944), .B2(new_n941), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n960), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT111), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n971), .B(new_n960), .C1(new_n965), .C2(new_n968), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n919), .B(new_n949), .C1(new_n954), .C2(new_n947), .ZN(new_n974));
  AND4_X1   g549(.A1(KEYINPUT43), .A2(new_n973), .A3(new_n875), .A4(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT44), .B1(new_n964), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n961), .B2(new_n963), .ZN(new_n979));
  AND4_X1   g554(.A1(new_n978), .A2(new_n973), .A3(new_n875), .A4(new_n974), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n976), .A2(new_n981), .ZN(G397));
  XNOR2_X1  g557(.A(new_n743), .B(new_n745), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n468), .A2(new_n476), .A3(G40), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n468), .A2(new_n476), .A3(KEYINPUT112), .A4(G40), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G1384), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n502), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  OR3_X1    g569(.A1(new_n983), .A2(KEYINPUT114), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G1996), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n994), .B1(new_n814), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(new_n996), .B2(new_n814), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT114), .B1(new_n983), .B2(new_n994), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n995), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  XOR2_X1   g575(.A(new_n723), .B(new_n725), .Z(new_n1001));
  OAI21_X1  g576(.A(new_n1000), .B1(new_n994), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n993), .A2(G1986), .A3(G290), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n993), .A2(new_n729), .A3(new_n592), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g580(.A(new_n1005), .B(KEYINPUT113), .Z(new_n1006));
  NOR2_X1   g581(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT126), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n502), .A2(new_n1009), .A3(new_n989), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1009), .B1(new_n502), .B2(new_n989), .ZN(new_n1011));
  NOR4_X1   g586(.A1(new_n988), .A2(new_n1010), .A3(new_n1011), .A4(G2084), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT119), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT45), .B1(new_n502), .B2(new_n989), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1013), .B1(new_n988), .B2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n992), .A2(KEYINPUT119), .A3(new_n986), .A4(new_n987), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n989), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1012), .B1(new_n1018), .B2(new_n822), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT51), .B1(new_n1019), .B2(G168), .ZN(new_n1020));
  INV_X1    g595(.A(G8), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(new_n1019), .B2(G168), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT62), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1027));
  AOI211_X1 g602(.A(G286), .B(new_n1012), .C1(new_n1018), .C2(new_n822), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT51), .B1(new_n1028), .B2(new_n1021), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT62), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  AND3_X1   g606(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n992), .A2(new_n986), .A3(new_n987), .A4(new_n1017), .ZN(new_n1035));
  INV_X1    g610(.A(G1971), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n986), .A2(new_n987), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n502), .A2(new_n1009), .A3(new_n989), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1011), .ZN(new_n1040));
  XNOR2_X1  g615(.A(KEYINPUT115), .B(G2090), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  AOI211_X1 g617(.A(new_n1021), .B(new_n1034), .C1(new_n1037), .C2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1034), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n989), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n988), .A2(new_n1045), .A3(new_n1014), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1042), .B1(new_n1046), .B2(G1971), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1044), .B1(new_n1047), .B2(G8), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1043), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G2078), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT53), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .A4(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1054), .B1(new_n1035), .B2(G2078), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1056));
  INV_X1    g631(.A(G1961), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1053), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G171), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n986), .A2(new_n989), .A3(new_n502), .A4(new_n987), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n570), .B(G1976), .C1(new_n571), .C2(new_n572), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(G8), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT52), .ZN(new_n1065));
  INV_X1    g640(.A(G1976), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT52), .B1(G288), .B2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1067), .A2(G8), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1062), .A2(G8), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n537), .B1(new_n582), .B2(new_n578), .ZN(new_n1071));
  OAI21_X1  g646(.A(G1981), .B1(new_n576), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g649(.A(KEYINPUT116), .B(G1981), .C1(new_n576), .C2(new_n1071), .ZN(new_n1075));
  INV_X1    g650(.A(G1981), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1074), .A2(new_n1075), .B1(new_n585), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT117), .B1(new_n1077), .B2(KEYINPUT49), .ZN(new_n1078));
  INV_X1    g653(.A(new_n576), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1071), .A2(KEYINPUT76), .ZN(new_n1080));
  AOI211_X1 g655(.A(new_n577), .B(new_n537), .C1(new_n582), .C2(new_n578), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1079), .B(new_n1076), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1075), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n516), .A2(new_n535), .A3(G86), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1084), .B(new_n574), .C1(new_n580), .C2(new_n537), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT116), .B1(new_n1085), .B2(G1981), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1082), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT49), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1070), .B1(new_n1078), .B2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(KEYINPUT49), .B(new_n1082), .C1(new_n1083), .C2(new_n1086), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1095), .A2(KEYINPUT118), .A3(KEYINPUT49), .A4(new_n1082), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1069), .B1(new_n1091), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1049), .A2(new_n1061), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  AND4_X1   g675(.A1(new_n1008), .A2(new_n1026), .A3(new_n1031), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1099), .B1(new_n1102), .B2(KEYINPUT62), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1008), .B1(new_n1103), .B2(new_n1031), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1106), .B(KEYINPUT57), .C1(new_n889), .C2(new_n890), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(KEYINPUT57), .ZN(new_n1108));
  OR2_X1    g683(.A1(new_n1106), .A2(KEYINPUT57), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n561), .A2(new_n565), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT56), .B(G2072), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1046), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1056), .A2(new_n788), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1062), .A2(G2067), .ZN(new_n1117));
  INV_X1    g692(.A(G1348), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1117), .B1(new_n1056), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1119), .A2(new_n609), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1112), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1116), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT61), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n988), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1124), .A2(G1956), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1113), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1035), .A2(new_n1126), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1125), .A2(new_n1127), .A3(new_n1111), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1123), .B1(new_n1128), .B2(new_n1116), .ZN(new_n1129));
  XOR2_X1   g704(.A(KEYINPUT58), .B(G1341), .Z(new_n1130));
  NAND2_X1  g705(.A1(new_n1062), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1062), .A2(KEYINPUT123), .A3(new_n1130), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT122), .B(G1996), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1133), .B(new_n1134), .C1(new_n1035), .C2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n554), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT59), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1111), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1140), .A2(KEYINPUT61), .A3(new_n1121), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1124), .A2(G1348), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1142), .B1(new_n1143), .B2(new_n1117), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1119), .A2(KEYINPUT60), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1144), .A2(new_n1145), .A3(new_n619), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1129), .A2(new_n1139), .A3(new_n1141), .A4(new_n1146), .ZN(new_n1147));
  OAI22_X1  g722(.A1(new_n1137), .A2(new_n1138), .B1(new_n619), .B2(new_n1145), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1122), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  OR4_X1    g724(.A1(new_n1014), .A2(new_n1045), .A3(new_n984), .A4(new_n1051), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1055), .A2(new_n1150), .A3(new_n1058), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1151), .A2(G171), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1053), .A2(new_n1055), .A3(new_n1058), .A4(G301), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT54), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT125), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1151), .A2(G171), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT125), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1156), .A2(new_n1157), .A3(KEYINPUT54), .A4(new_n1153), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n1151), .A2(G171), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT54), .B1(new_n1160), .B2(new_n1060), .ZN(new_n1161));
  AOI22_X1  g736(.A1(new_n1124), .A2(new_n1041), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1034), .B1(new_n1162), .B2(new_n1021), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1078), .A2(new_n1090), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1070), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1164), .A2(new_n1097), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1069), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n988), .A2(new_n1014), .ZN(new_n1168));
  AOI21_X1  g743(.A(G1971), .B1(new_n1168), .B2(new_n1017), .ZN(new_n1169));
  AND4_X1   g744(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1170));
  OAI211_X1 g745(.A(G8), .B(new_n1044), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1163), .A2(new_n1166), .A3(new_n1167), .A4(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1161), .A2(new_n1172), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1149), .A2(new_n1102), .A3(new_n1159), .A4(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1043), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1082), .ZN(new_n1176));
  NOR2_X1   g751(.A1(G288), .A2(G1976), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1176), .B1(new_n1166), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1175), .B1(new_n1178), .B2(new_n1070), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT63), .ZN(new_n1180));
  NAND2_X1  g755(.A1(G168), .A2(G8), .ZN(new_n1181));
  OR2_X1    g756(.A1(new_n1019), .A2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1180), .B1(new_n1172), .B2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1019), .A2(new_n1181), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1049), .A2(KEYINPUT63), .A3(new_n1098), .A4(new_n1184), .ZN(new_n1185));
  AOI211_X1 g760(.A(KEYINPUT120), .B(new_n1179), .C1(new_n1183), .C2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT120), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1179), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1174), .B1(new_n1186), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1007), .B1(new_n1105), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n994), .B1(new_n983), .B2(new_n815), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT46), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n993), .A2(new_n996), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1193), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1196), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1197));
  XOR2_X1   g772(.A(new_n1197), .B(KEYINPUT47), .Z(new_n1198));
  NOR2_X1   g773(.A1(new_n723), .A2(new_n725), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1000), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n848), .A2(new_n745), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n994), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  XOR2_X1   g777(.A(new_n1004), .B(KEYINPUT48), .Z(new_n1203));
  NOR2_X1   g778(.A1(new_n1002), .A2(new_n1203), .ZN(new_n1204));
  NOR3_X1   g779(.A1(new_n1198), .A2(new_n1202), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1192), .A2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g781(.A1(new_n979), .A2(new_n980), .ZN(new_n1208));
  NOR2_X1   g782(.A1(G227), .A2(new_n460), .ZN(new_n1209));
  XNOR2_X1  g783(.A(new_n1209), .B(KEYINPUT127), .ZN(new_n1210));
  NOR3_X1   g784(.A1(G401), .A2(new_n1210), .A3(G229), .ZN(new_n1211));
  OAI21_X1  g785(.A(new_n1211), .B1(new_n882), .B2(new_n879), .ZN(new_n1212));
  NOR2_X1   g786(.A1(new_n1208), .A2(new_n1212), .ZN(G308));
  OAI221_X1 g787(.A(new_n1211), .B1(new_n882), .B2(new_n879), .C1(new_n979), .C2(new_n980), .ZN(G225));
endmodule


