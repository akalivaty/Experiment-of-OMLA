//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1283, new_n1284,
    new_n1285, new_n1287, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1347,
    new_n1348, new_n1349, new_n1350;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n202), .A2(G77), .A3(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT65), .Z(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n204), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(new_n210), .A2(new_n211), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(G50), .ZN(new_n225));
  INV_X1    g0025(.A(G226), .ZN(new_n226));
  INV_X1    g0026(.A(G77), .ZN(new_n227));
  INV_X1    g0027(.A(G244), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n208), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n217), .B1(new_n211), .B2(new_n210), .C1(new_n230), .C2(KEYINPUT1), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT67), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n238), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n236), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT9), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  AND3_X1   g0051(.A1(new_n251), .A2(KEYINPUT69), .A3(new_n214), .ZN(new_n252));
  AOI21_X1  g0052(.A(KEYINPUT69), .B1(new_n251), .B2(new_n214), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT70), .A2(G58), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(KEYINPUT8), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G20), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n256), .A2(new_n258), .B1(G150), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n215), .B1(new_n201), .B2(new_n203), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT71), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n261), .A2(new_n262), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n254), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G13), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(new_n215), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n251), .A2(new_n214), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT69), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n251), .A2(KEYINPUT69), .A3(new_n214), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n225), .B1(new_n267), .B2(G20), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n274), .A2(new_n275), .B1(new_n225), .B2(new_n269), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n266), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  OAI211_X1 g0078(.A(G1), .B(G13), .C1(new_n257), .C2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT3), .B(G33), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G223), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  OR2_X1    g0085(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT3), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n286), .A2(new_n287), .A3(new_n289), .A4(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G222), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n291), .A2(new_n292), .B1(new_n227), .B2(new_n281), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n280), .B1(new_n285), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G45), .ZN(new_n295));
  AOI21_X1  g0095(.A(G1), .B1(new_n278), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G274), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n280), .A2(new_n296), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n298), .B1(new_n299), .B2(G226), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G200), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT79), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n250), .A2(new_n277), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(new_n250), .B2(new_n277), .ZN(new_n305));
  INV_X1    g0105(.A(new_n301), .ZN(new_n306));
  AOI21_X1  g0106(.A(KEYINPUT78), .B1(new_n306), .B2(G190), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n307), .B1(new_n303), .B2(new_n302), .ZN(new_n308));
  OR3_X1    g0108(.A1(new_n305), .A2(KEYINPUT10), .A3(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT10), .B1(new_n305), .B2(new_n308), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT72), .B(G179), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT73), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n314), .B(new_n277), .C1(G169), .C2(new_n306), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n298), .B1(new_n299), .B2(G238), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n287), .A2(new_n289), .A3(G232), .A4(G1698), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G97), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n318), .B(new_n319), .C1(new_n291), .C2(new_n226), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT80), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AND2_X1   g0122(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n323));
  NOR2_X1   g0123(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(new_n281), .A3(G226), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n326), .A2(KEYINPUT80), .A3(new_n318), .A4(new_n319), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n280), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n317), .B1(new_n322), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT13), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n320), .A2(new_n321), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(new_n327), .A3(new_n280), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(new_n333), .A3(new_n317), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n330), .A2(G190), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT81), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT81), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n330), .A2(new_n337), .A3(G190), .A4(new_n334), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT76), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n274), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G13), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n342), .A2(G1), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G20), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n344), .B1(new_n252), .B2(new_n253), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT76), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n267), .A2(G20), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n341), .A2(new_n346), .A3(G68), .A4(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G68), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n343), .A2(G20), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT12), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n258), .A2(G77), .ZN(new_n352));
  INV_X1    g0152(.A(new_n259), .ZN(new_n353));
  OAI221_X1 g0153(.A(new_n352), .B1(new_n215), .B2(G68), .C1(new_n225), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n254), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT11), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n351), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(new_n356), .B2(new_n355), .ZN(new_n358));
  AND3_X1   g0158(.A1(new_n332), .A2(new_n333), .A3(new_n317), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n333), .B1(new_n332), .B2(new_n317), .ZN(new_n360));
  OAI21_X1  g0160(.A(G200), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n339), .A2(new_n348), .A3(new_n358), .A4(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n358), .A2(new_n348), .ZN(new_n363));
  INV_X1    g0163(.A(G169), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n330), .B2(new_n334), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT14), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n330), .A2(new_n334), .ZN(new_n367));
  INV_X1    g0167(.A(G179), .ZN(new_n368));
  OAI22_X1  g0168(.A1(new_n365), .A2(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(G169), .B1(new_n359), .B2(new_n360), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n370), .A2(KEYINPUT14), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n363), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n362), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n298), .B1(new_n299), .B2(G232), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n286), .A2(new_n290), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n375), .A2(new_n283), .B1(new_n226), .B2(new_n284), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n288), .A2(G33), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT82), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n257), .B2(KEYINPUT3), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n288), .A2(KEYINPUT82), .A3(G33), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n377), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n376), .A2(new_n381), .B1(G33), .B2(G87), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n374), .B(new_n312), .C1(new_n382), .C2(new_n279), .ZN(new_n383));
  INV_X1    g0183(.A(new_n296), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n279), .ZN(new_n385));
  INV_X1    g0185(.A(G232), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n297), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n325), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n288), .A2(KEYINPUT82), .A3(G33), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT82), .B1(new_n288), .B2(G33), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n287), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI22_X1  g0191(.A1(new_n388), .A2(new_n391), .B1(new_n257), .B2(new_n219), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n387), .B1(new_n392), .B2(new_n280), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n383), .B1(new_n393), .B2(G169), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n391), .A2(new_n395), .A3(new_n215), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT7), .B1(new_n381), .B2(G20), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(new_n397), .A3(G68), .ZN(new_n398));
  INV_X1    g0198(.A(G58), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n399), .A2(new_n349), .ZN(new_n400));
  OR2_X1    g0200(.A1(new_n400), .A2(new_n203), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n401), .A2(G20), .B1(G159), .B2(new_n259), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n398), .A2(KEYINPUT16), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n402), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT84), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n287), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n289), .A2(KEYINPUT84), .ZN(new_n408));
  OAI211_X1 g0208(.A(KEYINPUT7), .B(new_n215), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n215), .B1(new_n377), .B2(new_n405), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT83), .B1(new_n410), .B2(new_n395), .ZN(new_n411));
  AOI21_X1  g0211(.A(G20), .B1(new_n287), .B2(new_n289), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT83), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n412), .A2(new_n413), .A3(KEYINPUT7), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n409), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n404), .B1(new_n415), .B2(G68), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n254), .B(new_n403), .C1(new_n416), .C2(KEYINPUT16), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n256), .A2(new_n347), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n345), .A2(new_n418), .B1(new_n344), .B2(new_n256), .ZN(new_n419));
  XNOR2_X1  g0219(.A(new_n419), .B(KEYINPUT85), .ZN(new_n420));
  AOI211_X1 g0220(.A(KEYINPUT18), .B(new_n394), .C1(new_n417), .C2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT18), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n415), .A2(G68), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT16), .B1(new_n423), .B2(new_n402), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n403), .A2(new_n254), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n420), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n394), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n422), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n421), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(G190), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n374), .B(new_n430), .C1(new_n382), .C2(new_n279), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n393), .B2(G200), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n420), .B(new_n432), .C1(new_n424), .C2(new_n425), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n433), .B(KEYINPUT17), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g0235(.A(KEYINPUT8), .B(G58), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n436), .A2(new_n353), .B1(new_n215), .B2(new_n227), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT74), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n219), .A2(KEYINPUT15), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT15), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(G87), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT75), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n439), .A2(new_n441), .A3(KEYINPUT75), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(new_n258), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT74), .ZN(new_n447));
  OAI221_X1 g0247(.A(new_n447), .B1(new_n215), .B2(new_n227), .C1(new_n436), .C2(new_n353), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n438), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n449), .A2(new_n254), .B1(new_n227), .B2(new_n269), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n341), .A2(new_n346), .A3(G77), .A4(new_n347), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n297), .B1(new_n385), .B2(new_n228), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n281), .A2(G238), .A3(G1698), .ZN(new_n454));
  INV_X1    g0254(.A(G107), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n281), .A2(G232), .ZN(new_n456));
  OAI221_X1 g0256(.A(new_n454), .B1(new_n455), .B2(new_n281), .C1(new_n456), .C2(new_n375), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n453), .B1(new_n457), .B2(new_n280), .ZN(new_n458));
  INV_X1    g0258(.A(new_n312), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OR2_X1    g0260(.A1(new_n458), .A2(new_n364), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n452), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT77), .B1(new_n450), .B2(new_n451), .ZN(new_n464));
  OAI22_X1  g0264(.A1(new_n456), .A2(new_n375), .B1(new_n455), .B2(new_n281), .ZN(new_n465));
  INV_X1    g0265(.A(new_n454), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n280), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n453), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n467), .A2(G190), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G200), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n469), .B1(new_n458), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n464), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n452), .A2(KEYINPUT77), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n463), .A2(new_n474), .ZN(new_n475));
  NOR4_X1   g0275(.A1(new_n316), .A2(new_n373), .A3(new_n435), .A4(new_n475), .ZN(new_n476));
  XOR2_X1   g0276(.A(KEYINPUT90), .B(KEYINPUT25), .Z(new_n477));
  NAND3_X1  g0277(.A1(new_n343), .A2(G20), .A3(new_n455), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT91), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n477), .A2(new_n478), .ZN(new_n480));
  OR2_X1    g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n480), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n267), .A2(G33), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n344), .B(new_n483), .C1(new_n252), .C2(new_n253), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n481), .B(new_n482), .C1(new_n455), .C2(new_n484), .ZN(new_n485));
  XOR2_X1   g0285(.A(KEYINPUT88), .B(KEYINPUT24), .Z(new_n486));
  OAI21_X1  g0286(.A(KEYINPUT23), .B1(new_n215), .B2(G107), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT23), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(new_n455), .A3(G20), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n215), .A2(G33), .A3(G116), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n487), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT22), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n287), .A2(new_n289), .A3(new_n215), .A4(G87), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n379), .A2(new_n380), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n492), .A2(new_n219), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n495), .A2(new_n215), .A3(new_n287), .A4(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n486), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n493), .A2(new_n492), .ZN(new_n499));
  INV_X1    g0299(.A(new_n491), .ZN(new_n500));
  AND4_X1   g0300(.A1(new_n497), .A2(new_n499), .A3(new_n500), .A4(new_n486), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n254), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT89), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(KEYINPUT89), .B(new_n254), .C1(new_n498), .C2(new_n501), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n485), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n267), .A2(G45), .ZN(new_n507));
  OR2_X1    g0307(.A1(KEYINPUT5), .A2(G41), .ZN(new_n508));
  NAND2_X1  g0308(.A1(KEYINPUT5), .A2(G41), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n280), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G264), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(G274), .ZN(new_n513));
  OAI22_X1  g0313(.A1(new_n375), .A2(new_n220), .B1(new_n222), .B2(new_n284), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n514), .A2(new_n381), .B1(G33), .B2(G294), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n512), .B(new_n513), .C1(new_n515), .C2(new_n279), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n516), .A2(G169), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n516), .A2(new_n368), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OR2_X1    g0319(.A1(new_n506), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n516), .A2(new_n470), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(G190), .B2(new_n516), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n506), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G283), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n287), .A2(new_n289), .A3(G250), .A4(G1698), .ZN(new_n527));
  NAND2_X1  g0327(.A1(KEYINPUT4), .A2(G244), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n526), .B(new_n527), .C1(new_n291), .C2(new_n528), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n323), .A2(new_n324), .A3(new_n228), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT4), .B1(new_n381), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n280), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n511), .A2(G257), .B1(G274), .B2(new_n510), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n532), .A2(new_n430), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(G200), .B1(new_n532), .B2(new_n533), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n413), .B1(new_n412), .B2(KEYINPUT7), .ZN(new_n537));
  OAI211_X1 g0337(.A(KEYINPUT83), .B(new_n395), .C1(new_n281), .C2(G20), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n455), .B1(new_n539), .B2(new_n409), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT6), .ZN(new_n541));
  NOR3_X1   g0341(.A1(new_n541), .A2(new_n221), .A3(G107), .ZN(new_n542));
  XNOR2_X1  g0342(.A(G97), .B(G107), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  OAI22_X1  g0344(.A1(new_n544), .A2(new_n215), .B1(new_n227), .B2(new_n353), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n254), .B1(new_n540), .B2(new_n545), .ZN(new_n546));
  MUX2_X1   g0346(.A(new_n344), .B(new_n484), .S(G97), .Z(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OR2_X1    g0348(.A1(new_n536), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n507), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G274), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n507), .A2(G250), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n279), .ZN(new_n554));
  INV_X1    g0354(.A(G116), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n257), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n286), .A2(G238), .A3(new_n290), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n228), .A2(new_n284), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n556), .B1(new_n560), .B2(new_n381), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n430), .B(new_n554), .C1(new_n561), .C2(new_n279), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n280), .B1(new_n552), .B2(new_n551), .ZN(new_n563));
  INV_X1    g0363(.A(new_n556), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n558), .B1(new_n325), .B2(G238), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n564), .B1(new_n565), .B2(new_n391), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n563), .B1(new_n566), .B2(new_n280), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n562), .B1(new_n567), .B2(G200), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n495), .A2(new_n215), .A3(G68), .A4(new_n287), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT19), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n215), .B1(new_n319), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(G87), .A2(G97), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n455), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n215), .A2(G33), .A3(G97), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n571), .A2(new_n573), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n254), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n444), .A2(new_n445), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n269), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n274), .A2(G87), .A3(new_n483), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n568), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT86), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n484), .B2(new_n578), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n439), .A2(new_n441), .A3(KEYINPUT75), .ZN(new_n585));
  AOI21_X1  g0385(.A(KEYINPUT75), .B1(new_n439), .B2(new_n441), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n274), .A2(new_n587), .A3(KEYINPUT86), .A4(new_n483), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n577), .A2(new_n584), .A3(new_n588), .A4(new_n579), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n554), .B1(new_n561), .B2(new_n279), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n364), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n312), .B(new_n554), .C1(new_n561), .C2(new_n279), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n589), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n582), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n532), .A2(new_n533), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G169), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n532), .A2(new_n459), .A3(new_n533), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n548), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n549), .A2(new_n595), .A3(new_n600), .ZN(new_n601));
  NOR3_X1   g0401(.A1(new_n323), .A2(new_n324), .A3(new_n222), .ZN(new_n602));
  AND2_X1   g0402(.A1(G264), .A2(G1698), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n381), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n282), .A2(G303), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n280), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n511), .A2(G270), .B1(G274), .B2(new_n510), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n269), .A2(new_n555), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n526), .B(new_n215), .C1(G33), .C2(new_n221), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT87), .ZN(new_n612));
  AOI21_X1  g0412(.A(G20), .B1(new_n257), .B2(G97), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT87), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n614), .A3(new_n526), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n251), .A2(new_n214), .B1(G20), .B2(new_n555), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n616), .A2(KEYINPUT20), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT20), .B1(new_n616), .B2(new_n617), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n610), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n555), .B1(new_n267), .B2(G33), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n341), .A2(new_n346), .A3(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(G169), .B(new_n609), .C1(new_n620), .C2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT21), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n279), .B1(new_n604), .B2(new_n605), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n508), .A2(new_n509), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n550), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n279), .ZN(new_n628));
  INV_X1    g0428(.A(G270), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n513), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(KEYINPUT21), .B(G169), .C1(new_n625), .C2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n607), .A2(G179), .A3(new_n608), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n341), .A2(new_n346), .A3(new_n621), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n634), .B(new_n610), .C1(new_n619), .C2(new_n618), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n623), .A2(new_n624), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n635), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n609), .A2(G190), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n625), .A2(new_n630), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(G200), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n637), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n636), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n601), .A2(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n476), .A2(new_n525), .A3(new_n643), .ZN(G372));
  NAND3_X1  g0444(.A1(new_n361), .A2(new_n348), .A3(new_n358), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n645), .B1(new_n336), .B2(new_n338), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n372), .B1(new_n646), .B2(new_n463), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n647), .A2(new_n434), .ZN(new_n648));
  INV_X1    g0448(.A(new_n429), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n311), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n650), .A2(new_n315), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n592), .B1(new_n567), .B2(G169), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT92), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n591), .A2(KEYINPUT92), .A3(new_n592), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(new_n589), .A3(new_n655), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n597), .A2(new_n598), .B1(new_n546), .B2(new_n547), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT93), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n576), .A2(new_n254), .B1(new_n269), .B2(new_n578), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT93), .B1(new_n662), .B2(new_n580), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n568), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n656), .A2(new_n657), .A3(new_n658), .A4(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(KEYINPUT26), .B1(new_n600), .B2(new_n594), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n665), .A2(new_n666), .A3(new_n656), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n636), .B1(new_n506), .B2(new_n519), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n536), .A2(new_n548), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(new_n657), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n584), .A2(new_n588), .ZN(new_n671));
  AOI22_X1  g0471(.A1(new_n652), .A2(new_n653), .B1(new_n662), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n659), .A2(new_n660), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n662), .A2(KEYINPUT93), .A3(new_n580), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n672), .A2(new_n655), .B1(new_n675), .B2(new_n568), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n668), .A2(new_n670), .A3(new_n523), .A4(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n667), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n476), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n651), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g0480(.A(new_n680), .B(KEYINPUT94), .Z(G369));
  OR3_X1    g0481(.A1(new_n268), .A2(KEYINPUT27), .A3(G20), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT27), .B1(new_n268), .B2(G20), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n637), .A2(new_n687), .ZN(new_n688));
  MUX2_X1   g0488(.A(new_n642), .B(new_n636), .S(new_n688), .Z(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT95), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n506), .A2(new_n687), .ZN(new_n693));
  OAI22_X1  g0493(.A1(new_n524), .A2(new_n693), .B1(new_n520), .B2(new_n687), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n524), .A2(new_n693), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n636), .A2(new_n686), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n520), .A2(new_n686), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT96), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n698), .A2(KEYINPUT96), .A3(new_n699), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n695), .A2(new_n704), .ZN(G399));
  INV_X1    g0505(.A(new_n209), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n572), .A2(new_n455), .A3(new_n555), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n708), .A2(G1), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n212), .B2(new_n708), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT31), .ZN(new_n714));
  INV_X1    g0514(.A(new_n632), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n514), .A2(new_n381), .ZN(new_n716));
  NAND2_X1  g0516(.A1(G33), .A2(G294), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n280), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n719), .A2(new_n512), .ZN(new_n720));
  INV_X1    g0520(.A(new_n596), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n715), .A2(new_n720), .A3(new_n721), .A4(new_n567), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n639), .A2(new_n567), .A3(new_n459), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(new_n516), .A3(new_n596), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n722), .B2(new_n723), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n714), .B(new_n686), .C1(new_n724), .C2(new_n727), .ZN(new_n728));
  NOR4_X1   g0528(.A1(new_n524), .A2(new_n601), .A3(new_n642), .A4(new_n686), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n686), .B1(new_n724), .B2(new_n727), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT31), .ZN(new_n731));
  OAI211_X1 g0531(.A(G330), .B(new_n728), .C1(new_n729), .C2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n657), .A2(new_n658), .A3(new_n593), .A4(new_n582), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT97), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n656), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n672), .A2(KEYINPUT97), .A3(new_n655), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n734), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n676), .A2(new_n657), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(KEYINPUT26), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n677), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n687), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT98), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n741), .A2(KEYINPUT98), .A3(new_n687), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(KEYINPUT29), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n686), .B1(new_n667), .B2(new_n677), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n748), .A2(KEYINPUT29), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n733), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n713), .B1(new_n750), .B2(G1), .ZN(G364));
  OR2_X1    g0551(.A1(new_n690), .A2(G330), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n342), .A2(G20), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G45), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n708), .A2(G1), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n752), .A2(new_n691), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(KEYINPUT99), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT99), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n752), .A2(new_n758), .A3(new_n691), .A4(new_n755), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n214), .B1(G20), .B2(new_n364), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n215), .A2(G190), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n459), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n470), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR4_X1   g0566(.A1(new_n312), .A2(new_n215), .A3(new_n430), .A4(G200), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n766), .A2(new_n349), .B1(new_n399), .B2(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n430), .A2(G179), .A3(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n215), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n221), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n470), .A2(G179), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(G20), .A3(G190), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n219), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n763), .A2(new_n773), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n281), .B1(new_n776), .B2(new_n455), .ZN(new_n777));
  NOR4_X1   g0577(.A1(new_n769), .A2(new_n772), .A3(new_n775), .A4(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT32), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G179), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n763), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G159), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n779), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n781), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n784), .A2(KEYINPUT32), .A3(G159), .ZN(new_n785));
  NOR4_X1   g0585(.A1(new_n312), .A2(new_n215), .A3(new_n430), .A4(new_n470), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n783), .A2(new_n785), .B1(new_n786), .B2(G50), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n764), .A2(G200), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n778), .B(new_n787), .C1(new_n227), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n767), .A2(G322), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT100), .ZN(new_n792));
  INV_X1    g0592(.A(G303), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n282), .B1(new_n774), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n791), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(G311), .B2(new_n788), .ZN(new_n796));
  INV_X1    g0596(.A(new_n776), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G283), .A2(new_n797), .B1(new_n784), .B2(G329), .ZN(new_n798));
  INV_X1    g0598(.A(G294), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n799), .B2(new_n771), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(G326), .B2(new_n786), .ZN(new_n801));
  XNOR2_X1  g0601(.A(KEYINPUT33), .B(G317), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n765), .A2(new_n802), .B1(new_n792), .B2(new_n794), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n796), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n762), .B1(new_n790), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G13), .A2(G33), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(G20), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n761), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n282), .A2(new_n706), .ZN(new_n810));
  AOI22_X1  g0610(.A1(G355), .A2(new_n810), .B1(new_n555), .B2(new_n706), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n213), .A2(G45), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(new_n245), .B2(G45), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n391), .A2(new_n209), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n811), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n755), .B(new_n805), .C1(new_n809), .C2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n808), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n690), .B2(new_n817), .ZN(new_n818));
  AND3_X1   g0618(.A1(new_n760), .A2(KEYINPUT101), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(KEYINPUT101), .B1(new_n760), .B2(new_n818), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G396));
  INV_X1    g0622(.A(new_n755), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n462), .A2(new_n687), .ZN(new_n824));
  INV_X1    g0624(.A(new_n452), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n472), .A2(new_n473), .B1(new_n825), .B2(new_n686), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n824), .B1(new_n826), .B2(new_n462), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n748), .A2(new_n828), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n686), .B(new_n827), .C1(new_n677), .C2(new_n667), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n823), .B1(new_n831), .B2(new_n733), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n732), .B1(new_n829), .B2(new_n830), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n762), .A2(new_n807), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n823), .B1(G77), .B2(new_n835), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n765), .A2(G150), .B1(G143), .B2(new_n767), .ZN(new_n837));
  INV_X1    g0637(.A(G137), .ZN(new_n838));
  INV_X1    g0638(.A(new_n786), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n837), .B1(new_n838), .B2(new_n839), .C1(new_n782), .C2(new_n789), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n840), .B(KEYINPUT34), .Z(new_n841));
  INV_X1    g0641(.A(new_n771), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n391), .B1(new_n842), .B2(G58), .ZN(new_n843));
  INV_X1    g0643(.A(new_n774), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n844), .A2(G50), .B1(new_n784), .B2(G132), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n797), .A2(G68), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n843), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n844), .A2(G107), .B1(new_n784), .B2(G311), .ZN(new_n848));
  INV_X1    g0648(.A(new_n772), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n797), .A2(G87), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n848), .A2(new_n849), .A3(new_n282), .A4(new_n850), .ZN(new_n851));
  AOI22_X1  g0651(.A1(G294), .A2(new_n767), .B1(new_n786), .B2(G303), .ZN(new_n852));
  INV_X1    g0652(.A(G283), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n852), .B1(new_n789), .B2(new_n555), .C1(new_n853), .C2(new_n766), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n841), .A2(new_n847), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n836), .B1(new_n855), .B2(new_n761), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n828), .B2(new_n807), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT102), .Z(new_n858));
  NOR2_X1   g0658(.A1(new_n834), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(G384));
  NOR2_X1   g0660(.A1(new_n753), .A2(new_n267), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT16), .B1(new_n398), .B2(new_n402), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n420), .B1(new_n425), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n684), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n429), .B2(new_n434), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n426), .A2(new_n427), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n426), .A2(new_n864), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n868), .A2(new_n869), .A3(new_n870), .A4(new_n433), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT105), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n871), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n863), .A2(new_n427), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n865), .A2(new_n874), .A3(new_n433), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT37), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT104), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n875), .A2(KEYINPUT104), .A3(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(KEYINPUT38), .B(new_n867), .C1(new_n873), .C2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  INV_X1    g0682(.A(new_n433), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n394), .B1(new_n417), .B2(new_n420), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n885), .A2(new_n872), .A3(new_n870), .A4(new_n869), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n871), .A2(KEYINPUT105), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n869), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n886), .A2(new_n887), .B1(KEYINPUT37), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n869), .B1(new_n429), .B2(new_n434), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n882), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n881), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n728), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n525), .A2(new_n643), .A3(new_n687), .ZN(new_n895));
  INV_X1    g0695(.A(new_n731), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n365), .A2(new_n366), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n370), .A2(KEYINPUT14), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n898), .B(new_n899), .C1(new_n368), .C2(new_n367), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n363), .B(new_n686), .C1(new_n646), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n363), .A2(new_n686), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n362), .A2(new_n372), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n897), .A2(new_n828), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT40), .B1(new_n893), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(KEYINPUT40), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n867), .B1(new_n873), .B2(new_n880), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n882), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n881), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n476), .A2(new_n897), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n912), .B(new_n913), .Z(new_n914));
  INV_X1    g0714(.A(G330), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n900), .A2(new_n363), .A3(new_n687), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT39), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n909), .B2(new_n881), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n881), .A2(new_n891), .A3(new_n920), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n429), .A2(new_n864), .ZN(new_n924));
  INV_X1    g0724(.A(new_n824), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n748), .B2(new_n828), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n901), .A2(new_n903), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT103), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT103), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n929), .B(new_n904), .C1(new_n830), .C2(new_n925), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n924), .B1(new_n931), .B2(new_n910), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n923), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n747), .A2(new_n476), .A3(new_n749), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n651), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n933), .B(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n861), .B1(new_n917), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n936), .B2(new_n917), .ZN(new_n938));
  INV_X1    g0738(.A(new_n544), .ZN(new_n939));
  OAI211_X1 g0739(.A(G116), .B(new_n216), .C1(new_n939), .C2(KEYINPUT35), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(KEYINPUT35), .B2(new_n939), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT36), .Z(new_n942));
  NOR2_X1   g0742(.A1(new_n202), .A2(new_n349), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n212), .A2(new_n227), .A3(new_n400), .ZN(new_n944));
  OAI211_X1 g0744(.A(G1), .B(new_n342), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n938), .A2(new_n942), .A3(new_n945), .ZN(G367));
  INV_X1    g0746(.A(KEYINPUT106), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n548), .A2(new_n686), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n670), .A2(new_n948), .ZN(new_n949));
  OR3_X1    g0749(.A1(new_n698), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n947), .B1(new_n698), .B2(new_n949), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n600), .B1(new_n949), .B2(new_n520), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n952), .A2(KEYINPUT42), .B1(new_n687), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT107), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n952), .B2(KEYINPUT42), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT42), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n950), .A2(KEYINPUT107), .A3(new_n957), .A4(new_n951), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n954), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n675), .A2(new_n687), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n656), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n676), .B2(new_n960), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT108), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n959), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n959), .B(new_n965), .C1(KEYINPUT43), .C2(new_n963), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n657), .A2(new_n686), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n949), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n970), .B1(new_n695), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n695), .A2(new_n973), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n968), .A2(new_n975), .A3(new_n969), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n707), .B(KEYINPUT41), .Z(new_n977));
  INV_X1    g0777(.A(new_n695), .ZN(new_n978));
  AND3_X1   g0778(.A1(new_n698), .A2(KEYINPUT96), .A3(new_n699), .ZN(new_n979));
  AOI21_X1  g0779(.A(KEYINPUT96), .B1(new_n698), .B2(new_n699), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n972), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n704), .A2(KEYINPUT45), .A3(new_n972), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n702), .A2(new_n703), .A3(new_n973), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT44), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT44), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n702), .A2(new_n988), .A3(new_n703), .A4(new_n973), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n978), .B1(new_n985), .B2(new_n990), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n987), .A2(new_n989), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n983), .A2(new_n984), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n992), .A2(new_n695), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n692), .A2(KEYINPUT109), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT109), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n691), .A2(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n694), .A2(new_n697), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n998), .A2(new_n698), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n995), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  OR3_X1    g0800(.A1(new_n999), .A2(new_n691), .A3(new_n996), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n991), .A2(new_n750), .A3(new_n994), .A4(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n977), .B1(new_n1003), .B2(new_n750), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n754), .A2(G1), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n974), .B(new_n976), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n241), .A2(new_n814), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n809), .B1(new_n578), .B2(new_n209), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n823), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n765), .A2(G159), .B1(G143), .B2(new_n786), .ZN(new_n1010));
  INV_X1    g0810(.A(G150), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1010), .B1(new_n1011), .B2(new_n768), .C1(new_n201), .C2(new_n789), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n771), .A2(new_n349), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n281), .B1(new_n774), .B2(new_n399), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n776), .A2(new_n227), .B1(new_n781), .B2(new_n838), .ZN(new_n1015));
  NOR4_X1   g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n788), .A2(G283), .B1(G311), .B2(new_n786), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n793), .B2(new_n768), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G97), .A2(new_n797), .B1(new_n784), .B2(G317), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n391), .B(new_n1019), .C1(new_n766), .C2(new_n799), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n844), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT46), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n774), .B2(new_n555), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1021), .B(new_n1023), .C1(new_n455), .C2(new_n771), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1018), .A2(new_n1020), .A3(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1016), .A2(new_n1025), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1026), .A2(KEYINPUT47), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n762), .B1(new_n1026), .B2(KEYINPUT47), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1009), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n817), .B2(new_n963), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1006), .A2(new_n1030), .ZN(G387));
  NAND2_X1  g0831(.A1(new_n844), .A2(G77), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n221), .B2(new_n776), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n391), .B(new_n1033), .C1(G150), .C2(new_n784), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n587), .A2(new_n842), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n765), .A2(new_n256), .B1(G50), .B2(new_n767), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n788), .A2(G68), .B1(G159), .B2(new_n786), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(KEYINPUT111), .B(G322), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n839), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n765), .A2(G311), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n788), .A2(G303), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n767), .A2(G317), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1045), .A2(KEYINPUT48), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n771), .A2(new_n853), .B1(new_n774), .B2(new_n799), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n1045), .B2(KEYINPUT48), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1046), .A2(KEYINPUT49), .A3(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G116), .A2(new_n797), .B1(new_n784), .B2(G326), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(new_n391), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(KEYINPUT49), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1038), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1053), .A2(KEYINPUT112), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(KEYINPUT112), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1054), .A2(new_n761), .A3(new_n1055), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n694), .A2(new_n817), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n710), .B(new_n295), .C1(new_n349), .C2(new_n227), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n436), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n225), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1058), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n814), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n236), .B2(new_n295), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n810), .A2(new_n709), .B1(new_n455), .B2(new_n706), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n755), .B1(new_n1067), .B2(new_n809), .ZN(new_n1068));
  AND3_X1   g0868(.A1(new_n1056), .A2(new_n1057), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1002), .A2(new_n750), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n707), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1002), .A2(new_n750), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1070), .B1(new_n1072), .B2(new_n1073), .ZN(G393));
  AND2_X1   g0874(.A1(new_n1003), .A2(new_n707), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n994), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n695), .B1(new_n992), .B2(new_n993), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1071), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(KEYINPUT115), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1078), .A2(new_n1003), .A3(KEYINPUT115), .A4(new_n707), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n973), .A2(new_n808), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n809), .B1(new_n221), .B2(new_n209), .C1(new_n248), .C2(new_n814), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n823), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G150), .A2(new_n786), .B1(new_n767), .B2(G159), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT51), .Z(new_n1086));
  OAI21_X1  g0886(.A(new_n850), .B1(new_n349), .B2(new_n774), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n842), .A2(G77), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n381), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1087), .B(new_n1089), .C1(G143), .C2(new_n784), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n202), .A2(new_n765), .B1(new_n788), .B2(new_n1059), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1086), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n765), .A2(G303), .B1(G116), .B2(new_n842), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(KEYINPUT114), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n774), .A2(new_n853), .B1(new_n781), .B2(new_n1039), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n281), .B(new_n1095), .C1(G107), .C2(new_n797), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1094), .B(new_n1096), .C1(new_n799), .C2(new_n789), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G311), .A2(new_n767), .B1(new_n786), .B2(G317), .ZN(new_n1098));
  XOR2_X1   g0898(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n1099));
  XNOR2_X1  g0899(.A(new_n1098), .B(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(KEYINPUT114), .B2(new_n1093), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1092), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1084), .B1(new_n1102), .B2(new_n761), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1081), .A2(new_n1005), .B1(new_n1082), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1080), .A2(new_n1104), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1079), .A2(new_n1105), .ZN(G390));
  NAND4_X1  g0906(.A1(new_n897), .A2(G330), .A3(new_n828), .A4(new_n904), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n748), .A2(new_n828), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n824), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n919), .B1(new_n1110), .B2(new_n904), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n921), .A2(new_n922), .A3(new_n1111), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n875), .A2(KEYINPUT104), .A3(KEYINPUT37), .ZN(new_n1113));
  AOI21_X1  g0913(.A(KEYINPUT104), .B1(new_n875), .B2(KEYINPUT37), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n886), .A2(new_n887), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n882), .B(new_n866), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n888), .A2(KEYINPUT37), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n871), .A2(KEYINPUT105), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n871), .A2(KEYINPUT105), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n890), .ZN(new_n1122));
  AOI21_X1  g0922(.A(KEYINPUT38), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n918), .B1(new_n1117), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n826), .A2(new_n462), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n734), .A2(new_n736), .A3(new_n737), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n658), .B1(new_n676), .B2(new_n657), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n743), .B(new_n686), .C1(new_n1129), .C2(new_n677), .ZN(new_n1130));
  AOI21_X1  g0930(.A(KEYINPUT98), .B1(new_n741), .B2(new_n687), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1126), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n824), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1124), .B1(new_n904), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1108), .B1(new_n1112), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n925), .B1(new_n746), .B2(new_n1126), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n918), .B(new_n892), .C1(new_n1136), .C2(new_n927), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1111), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1139));
  AOI21_X1  g0939(.A(KEYINPUT38), .B1(new_n1139), .B2(new_n867), .ZN(new_n1140));
  OAI21_X1  g0940(.A(KEYINPUT39), .B1(new_n1140), .B2(new_n1117), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n881), .A2(new_n891), .A3(new_n920), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1138), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1137), .A2(new_n1143), .A3(new_n1107), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1135), .A2(new_n1144), .A3(new_n1005), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT117), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1145), .B(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1135), .A2(new_n1144), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT116), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n927), .B1(new_n732), .B2(new_n827), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n1107), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n926), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1133), .A2(new_n1107), .A3(new_n1150), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n476), .A2(G330), .A3(new_n897), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n934), .A2(new_n651), .A3(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1148), .A2(new_n1149), .A3(new_n1158), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1135), .B(new_n1144), .C1(new_n1157), .C2(KEYINPUT116), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(new_n1160), .A3(new_n707), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n823), .B1(new_n256), .B2(new_n835), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n282), .B1(new_n784), .B2(G125), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n201), .B2(new_n776), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G159), .B2(new_n842), .ZN(new_n1165));
  INV_X1    g0965(.A(G132), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n768), .C1(new_n838), .C2(new_n766), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n774), .A2(new_n1011), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT53), .ZN(new_n1169));
  INV_X1    g0969(.A(G128), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT54), .B(G143), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1169), .B1(new_n1170), .B2(new_n839), .C1(new_n789), .C2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n775), .A2(new_n281), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n784), .A2(G294), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1173), .A2(new_n1088), .A3(new_n846), .A4(new_n1174), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(G116), .A2(new_n767), .B1(new_n786), .B2(G283), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1176), .B1(new_n789), .B2(new_n221), .C1(new_n455), .C2(new_n766), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n1167), .A2(new_n1172), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1162), .B1(new_n1178), .B2(new_n761), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n921), .A2(new_n922), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1179), .B1(new_n1181), .B2(new_n807), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1147), .A2(new_n1161), .A3(new_n1182), .ZN(G378));
  INV_X1    g0983(.A(new_n277), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1184), .A2(new_n684), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n316), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n316), .A2(new_n1185), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1188), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n923), .A2(new_n932), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1191), .B1(new_n923), .B2(new_n932), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n915), .B1(new_n906), .B2(new_n911), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n912), .A2(G330), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1191), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n931), .A2(new_n910), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n924), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n918), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1197), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n923), .A2(new_n932), .A3(new_n1191), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1196), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(KEYINPUT118), .B1(new_n1195), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1194), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1202), .A2(new_n1196), .A3(new_n1203), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT118), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1205), .A2(new_n1005), .A3(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1191), .A2(new_n806), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n823), .B1(new_n202), .B2(new_n835), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n771), .A2(new_n1011), .B1(new_n774), .B2(new_n1171), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n788), .A2(G137), .B1(G128), .B2(new_n767), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n1166), .B2(new_n766), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1213), .B(new_n1215), .C1(G125), .C2(new_n786), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT59), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n257), .B(new_n278), .C1(new_n776), .C2(new_n782), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G124), .B2(new_n784), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1218), .A2(new_n1219), .A3(new_n1221), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n765), .A2(G97), .B1(G107), .B2(new_n767), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n578), .B2(new_n789), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n797), .A2(G58), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n784), .A2(G283), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1032), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n278), .B(new_n391), .C1(new_n839), .C2(new_n555), .ZN(new_n1228));
  NOR4_X1   g1028(.A1(new_n1224), .A2(new_n1013), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(KEYINPUT58), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n1229), .A2(KEYINPUT58), .ZN(new_n1231));
  AOI21_X1  g1031(.A(G50), .B1(new_n257), .B2(new_n278), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n381), .B2(G41), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1222), .A2(new_n1230), .A3(new_n1231), .A4(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1212), .B1(new_n1234), .B2(new_n761), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1211), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1210), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1154), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1135), .A2(new_n1144), .A3(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1156), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1205), .A2(new_n1241), .A3(new_n1209), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT57), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1243), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n707), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1237), .B1(new_n1244), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(G375));
  OAI21_X1  g1051(.A(new_n823), .B1(G68), .B2(new_n835), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n767), .A2(G137), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1253), .B1(new_n1166), .B2(new_n839), .C1(new_n766), .C2(new_n1171), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT122), .ZN(new_n1255));
  OR2_X1    g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n381), .B1(new_n771), .B2(new_n225), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n1225), .B1(new_n1170), .B2(new_n781), .C1(new_n782), .C2(new_n774), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n1258), .B(new_n1259), .C1(G150), .C2(new_n788), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1256), .A2(new_n1257), .A3(new_n1260), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n455), .A2(new_n789), .B1(new_n766), .B2(new_n555), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n1262), .A2(KEYINPUT119), .B1(new_n799), .B2(new_n839), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(KEYINPUT119), .B2(new_n1262), .ZN(new_n1264));
  XOR2_X1   g1064(.A(new_n1264), .B(KEYINPUT120), .Z(new_n1265));
  OAI22_X1  g1065(.A1(new_n774), .A2(new_n221), .B1(new_n781), .B2(new_n793), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT121), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n767), .A2(G283), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n281), .B1(new_n797), .B2(G77), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1267), .A2(new_n1035), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1261), .B1(new_n1265), .B2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1252), .B1(new_n1271), .B2(new_n761), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n904), .B2(new_n807), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1005), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1273), .B1(new_n1154), .B2(new_n1274), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1275), .B(KEYINPUT123), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n977), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1158), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1277), .A2(new_n1280), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(KEYINPUT124), .ZN(G381));
  OR4_X1    g1082(.A1(G396), .A2(G387), .A3(G384), .A4(G393), .ZN(new_n1283));
  INV_X1    g1083(.A(G378), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1250), .A2(new_n1284), .ZN(new_n1285));
  OR4_X1    g1085(.A1(G390), .A2(new_n1283), .A3(new_n1285), .A4(G381), .ZN(G407));
  INV_X1    g1086(.A(G213), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1287), .A2(G343), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1285), .A2(new_n1289), .ZN(new_n1290));
  XOR2_X1   g1090(.A(new_n1290), .B(KEYINPUT125), .Z(new_n1291));
  NAND3_X1  g1091(.A1(new_n1291), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1092(.A(KEYINPUT60), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(new_n1279), .B(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1158), .A2(new_n707), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1277), .B(G384), .C1(new_n1294), .C2(new_n1295), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n859), .B1(new_n1297), .B2(new_n1276), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1248), .B1(new_n1243), .B2(new_n1242), .ZN(new_n1301));
  NOR3_X1   g1101(.A1(new_n1301), .A2(new_n1284), .A3(new_n1237), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1205), .A2(new_n1278), .A3(new_n1241), .A4(new_n1209), .ZN(new_n1303));
  AOI22_X1  g1103(.A1(new_n1246), .A2(new_n1005), .B1(new_n1211), .B2(new_n1235), .ZN(new_n1304));
  AOI21_X1  g1104(.A(G378), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n1289), .B(new_n1300), .C1(new_n1302), .C2(new_n1305), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT61), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1244), .A2(new_n1249), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1237), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1310), .A2(new_n1311), .A3(G378), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1305), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT62), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1314), .A2(new_n1315), .A3(new_n1289), .A4(new_n1300), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1288), .A2(G2897), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1296), .A2(new_n1298), .A3(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1317), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1305), .B1(new_n1250), .B2(G378), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1321), .B1(new_n1322), .B2(new_n1288), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1308), .A2(new_n1309), .A3(new_n1316), .A4(new_n1323), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1079), .A2(new_n1105), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(G387), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1006), .B(new_n1030), .C1(new_n1079), .C2(new_n1105), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(G393), .B(new_n821), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT126), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1326), .A2(new_n1327), .A3(new_n1330), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1325), .B(G387), .C1(new_n1329), .C2(new_n1328), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(G390), .A2(new_n1006), .A3(new_n1030), .A4(new_n1328), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1331), .A2(new_n1332), .A3(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1324), .A2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1334), .A2(new_n1309), .ZN(new_n1337));
  NOR3_X1   g1137(.A1(new_n1322), .A2(new_n1288), .A3(new_n1299), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1337), .B1(new_n1338), .B2(KEYINPUT63), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1320), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(new_n1318), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1341), .B1(new_n1314), .B2(new_n1289), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT63), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1306), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1339), .A2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1336), .A2(new_n1345), .ZN(G405));
  NAND2_X1  g1146(.A1(new_n1334), .A2(new_n1299), .ZN(new_n1347));
  NAND4_X1  g1147(.A1(new_n1331), .A2(new_n1333), .A3(new_n1332), .A4(new_n1300), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  XNOR2_X1  g1149(.A(new_n1250), .B(G378), .ZN(new_n1350));
  XNOR2_X1  g1150(.A(new_n1349), .B(new_n1350), .ZN(G402));
endmodule


