//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 1 0 0 0 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n633, new_n634, new_n635, new_n638, new_n640,
    new_n641, new_n642, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1202, new_n1203,
    new_n1204;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n460), .A2(G101), .A3(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n461), .B(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n464), .B1(new_n465), .B2(KEYINPUT68), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n460), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n463), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n460), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n472), .A2(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(new_n470), .A2(KEYINPUT70), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n466), .B2(new_n468), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G112), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n487));
  OR2_X1    g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n487), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n460), .B1(new_n466), .B2(new_n468), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n488), .A2(new_n489), .B1(G124), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n483), .A2(new_n491), .ZN(new_n492));
  XOR2_X1   g067(.A(new_n492), .B(KEYINPUT72), .Z(G162));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n494), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n473), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT76), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n473), .A2(KEYINPUT76), .A3(new_n495), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n501), .B1(new_n479), .B2(G138), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n490), .A2(G126), .ZN(new_n504));
  OAI21_X1  g079(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(G114), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n460), .B1(KEYINPUT73), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT73), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G114), .ZN(new_n509));
  AOI211_X1 g084(.A(KEYINPUT74), .B(new_n505), .C1(new_n507), .C2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT74), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n506), .A2(KEYINPUT73), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n509), .A2(new_n512), .A3(G2105), .ZN(new_n513));
  INV_X1    g088(.A(new_n505), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n504), .B1(new_n510), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT75), .ZN(new_n517));
  OAI21_X1  g092(.A(G2105), .B1(new_n508), .B2(G114), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n506), .A2(KEYINPUT73), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n514), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT74), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n513), .A2(new_n511), .A3(new_n514), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT75), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(new_n524), .A3(new_n504), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n503), .B1(new_n517), .B2(new_n525), .ZN(G164));
  INV_X1    g101(.A(G543), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT6), .ZN(new_n528));
  INV_X1    g103(.A(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(KEYINPUT6), .A2(G651), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G50), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT77), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n533), .B(new_n534), .ZN(new_n535));
  OR2_X1    g110(.A1(KEYINPUT5), .A2(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(KEYINPUT5), .A2(G543), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n538), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n530), .A2(new_n531), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(G88), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n539), .A2(new_n529), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n535), .A2(new_n543), .ZN(G166));
  INV_X1    g119(.A(new_n538), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n529), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n546), .A2(G63), .B1(G51), .B2(new_n532), .ZN(new_n547));
  NAND3_X1  g122(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT7), .ZN(new_n549));
  INV_X1    g124(.A(G89), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n541), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n547), .B1(KEYINPUT78), .B2(new_n551), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n551), .A2(KEYINPUT78), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n552), .A2(new_n553), .ZN(G168));
  AOI22_X1  g129(.A1(new_n538), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n529), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n532), .A2(G52), .ZN(new_n557));
  XOR2_X1   g132(.A(KEYINPUT79), .B(G90), .Z(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n541), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n556), .A2(new_n559), .ZN(G171));
  AOI22_X1  g135(.A1(new_n538), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(new_n529), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n532), .A2(G43), .ZN(new_n563));
  INV_X1    g138(.A(G81), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n541), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT80), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n565), .A2(new_n566), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n562), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G860), .ZN(G153));
  NAND4_X1  g146(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND4_X1  g149(.A1(G319), .A2(G483), .A3(G661), .A4(new_n574), .ZN(G188));
  NAND2_X1  g150(.A1(new_n532), .A2(G53), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT9), .ZN(new_n577));
  NAND2_X1  g152(.A1(G78), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G65), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n545), .B2(new_n579), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n538), .A2(new_n540), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n580), .A2(G651), .B1(new_n581), .B2(G91), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n577), .A2(new_n582), .ZN(G299));
  INV_X1    g158(.A(G171), .ZN(G301));
  INV_X1    g159(.A(G168), .ZN(G286));
  INV_X1    g160(.A(G166), .ZN(G303));
  OAI21_X1  g161(.A(G651), .B1(new_n538), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT81), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT81), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n589), .B(G651), .C1(new_n538), .C2(G74), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n532), .A2(G49), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n538), .A2(new_n540), .A3(G87), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n588), .A2(new_n590), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(KEYINPUT82), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n591), .A2(new_n592), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT82), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n595), .A2(new_n596), .A3(new_n588), .A4(new_n590), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G288));
  INV_X1    g174(.A(KEYINPUT83), .ZN(new_n600));
  INV_X1    g175(.A(G61), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(new_n536), .B2(new_n537), .ZN(new_n602));
  AND2_X1   g177(.A1(G73), .A2(G543), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n600), .B(G651), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n532), .A2(G48), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT84), .ZN(new_n607));
  INV_X1    g182(.A(G86), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n541), .B2(new_n608), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n538), .A2(new_n540), .A3(KEYINPUT84), .A4(G86), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(G651), .B1(new_n602), .B2(new_n603), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(KEYINPUT83), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n606), .A2(new_n611), .A3(new_n613), .ZN(G305));
  AOI22_X1  g189(.A1(new_n538), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n615), .A2(new_n529), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n532), .A2(G47), .ZN(new_n617));
  INV_X1    g192(.A(G85), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n541), .B2(new_n618), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n616), .A2(new_n619), .ZN(G290));
  INV_X1    g195(.A(G868), .ZN(new_n621));
  NOR2_X1   g196(.A1(G301), .A2(new_n621), .ZN(new_n622));
  AND3_X1   g197(.A1(new_n538), .A2(new_n540), .A3(G92), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT10), .ZN(new_n624));
  NAND2_X1  g199(.A1(G79), .A2(G543), .ZN(new_n625));
  INV_X1    g200(.A(G66), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n545), .B2(new_n626), .ZN(new_n627));
  AOI22_X1  g202(.A1(new_n627), .A2(G651), .B1(G54), .B2(new_n532), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT85), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n622), .B1(new_n630), .B2(new_n621), .ZN(G284));
  AOI21_X1  g206(.A(new_n622), .B1(new_n630), .B2(new_n621), .ZN(G321));
  INV_X1    g207(.A(G299), .ZN(new_n633));
  OAI21_X1  g208(.A(KEYINPUT86), .B1(new_n633), .B2(G868), .ZN(new_n634));
  NOR2_X1   g209(.A1(G168), .A2(new_n621), .ZN(new_n635));
  MUX2_X1   g210(.A(new_n634), .B(KEYINPUT86), .S(new_n635), .Z(G297));
  MUX2_X1   g211(.A(new_n634), .B(KEYINPUT86), .S(new_n635), .Z(G280));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n630), .B1(new_n638), .B2(G860), .ZN(G148));
  NAND2_X1  g214(.A1(new_n569), .A2(new_n621), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n630), .A2(new_n638), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n640), .B1(new_n642), .B2(new_n621), .ZN(G323));
  XNOR2_X1  g218(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g219(.A1(new_n482), .A2(G135), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n490), .A2(G123), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n460), .A2(G111), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n645), .B(new_n646), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT87), .B(G2096), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n460), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT12), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT13), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2100), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n651), .A2(new_n655), .ZN(G156));
  XOR2_X1   g231(.A(KEYINPUT15), .B(G2435), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2438), .ZN(new_n658));
  XOR2_X1   g233(.A(G2427), .B(G2430), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT88), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(KEYINPUT14), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2451), .B(G2454), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT16), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1341), .B(G1348), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n663), .B(new_n667), .Z(new_n668));
  XNOR2_X1  g243(.A(G2443), .B(G2446), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(new_n671), .A3(G14), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G401));
  XNOR2_X1  g248(.A(G2084), .B(G2090), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT89), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2072), .B(G2078), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2067), .B(G2678), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT18), .Z(new_n679));
  NOR2_X1   g254(.A1(new_n675), .A2(new_n677), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n675), .A2(new_n677), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n676), .B(KEYINPUT17), .Z(new_n683));
  NAND3_X1  g258(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n676), .B(KEYINPUT90), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n679), .B(new_n684), .C1(new_n681), .C2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G2096), .B(G2100), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n688), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(G227));
  XNOR2_X1  g266(.A(G1956), .B(G2474), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT91), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1961), .B(G1966), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1971), .B(G1976), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT19), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT20), .Z(new_n700));
  OR2_X1    g275(.A1(new_n693), .A2(new_n695), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n701), .A2(new_n698), .A3(new_n696), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n700), .B(new_n702), .C1(new_n698), .C2(new_n701), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1991), .B(G1996), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1981), .B(G1986), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n707), .A2(new_n709), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(G229));
  OAI21_X1  g287(.A(KEYINPUT100), .B1(G16), .B2(G21), .ZN(new_n713));
  NAND2_X1  g288(.A1(G168), .A2(G16), .ZN(new_n714));
  MUX2_X1   g289(.A(KEYINPUT100), .B(new_n713), .S(new_n714), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1966), .ZN(new_n716));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  NOR2_X1   g292(.A1(G171), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G5), .B2(new_n717), .ZN(new_n719));
  INV_X1    g294(.A(G1961), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  OAI22_X1  g296(.A1(new_n719), .A2(new_n720), .B1(new_n721), .B2(new_n649), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n719), .A2(new_n720), .ZN(new_n723));
  INV_X1    g298(.A(G28), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(KEYINPUT30), .ZN(new_n725));
  AOI21_X1  g300(.A(G29), .B1(new_n724), .B2(KEYINPUT30), .ZN(new_n726));
  OR2_X1    g301(.A1(KEYINPUT31), .A2(G11), .ZN(new_n727));
  NAND2_X1  g302(.A1(KEYINPUT31), .A2(G11), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n725), .A2(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n723), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G2084), .ZN(new_n731));
  NAND2_X1  g306(.A1(G160), .A2(G29), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT24), .B(G34), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(new_n721), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT97), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  AOI211_X1 g311(.A(new_n722), .B(new_n730), .C1(new_n731), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n482), .A2(G141), .ZN(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT26), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n460), .A2(G105), .A3(G2104), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT98), .ZN(new_n742));
  AOI211_X1 g317(.A(new_n740), .B(new_n742), .C1(G129), .C2(new_n490), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(new_n721), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n721), .B2(G32), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT27), .B(G1996), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n717), .A2(G20), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT23), .Z(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G299), .B2(G16), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1956), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n716), .A2(new_n737), .A3(new_n749), .A4(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT95), .ZN(new_n755));
  NOR2_X1   g330(.A1(G16), .A2(G19), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n570), .B2(G16), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT94), .B(G1341), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n721), .A2(G26), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT28), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n482), .A2(G140), .ZN(new_n762));
  OAI21_X1  g337(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n763));
  INV_X1    g338(.A(G116), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(G2105), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n490), .B2(G128), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n761), .B1(new_n767), .B2(G29), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G2067), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n630), .A2(G16), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G4), .B2(G16), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n771), .A2(G1348), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(G1348), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n759), .B(new_n769), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n754), .B1(new_n755), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n721), .A2(G27), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G164), .B2(new_n721), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT101), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G2078), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n482), .A2(G139), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT25), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n473), .A2(G127), .ZN(new_n784));
  AND2_X1   g359(.A1(G115), .A2(G2104), .ZN(new_n785));
  OAI21_X1  g360(.A(G2105), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT96), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n781), .B(new_n788), .C1(new_n787), .C2(new_n786), .ZN(new_n789));
  MUX2_X1   g364(.A(G33), .B(new_n789), .S(G29), .Z(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(G2072), .Z(new_n791));
  NOR2_X1   g366(.A1(new_n736), .A2(new_n731), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n747), .B2(new_n748), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT99), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n721), .A2(G35), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G162), .B2(new_n721), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT29), .Z(new_n798));
  INV_X1    g373(.A(G2090), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n795), .B(new_n800), .C1(new_n755), .C2(new_n774), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n780), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n798), .A2(new_n799), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT102), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n717), .A2(G22), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G166), .B2(new_n717), .ZN(new_n806));
  INV_X1    g381(.A(G1971), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(G6), .A2(G16), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G305), .B2(new_n717), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT32), .B(G1981), .Z(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  MUX2_X1   g388(.A(G23), .B(new_n593), .S(G16), .Z(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT33), .B(G1976), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n808), .A2(new_n812), .A3(new_n813), .A4(new_n816), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n482), .A2(G131), .ZN(new_n820));
  OAI21_X1  g395(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n821));
  INV_X1    g396(.A(G107), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n821), .B1(new_n822), .B2(G2105), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n490), .B2(G119), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G29), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G25), .B2(G29), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT35), .B(G1991), .Z(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n717), .A2(G24), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT92), .ZN(new_n832));
  INV_X1    g407(.A(G290), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(new_n717), .ZN(new_n834));
  AOI21_X1  g409(.A(KEYINPUT93), .B1(new_n834), .B2(G1986), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n830), .B(new_n835), .C1(G1986), .C2(new_n834), .ZN(new_n836));
  NOR4_X1   g411(.A1(new_n818), .A2(new_n819), .A3(new_n829), .A4(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT36), .Z(new_n838));
  AND3_X1   g413(.A1(new_n802), .A2(new_n804), .A3(new_n838), .ZN(G311));
  NAND3_X1  g414(.A1(new_n802), .A2(new_n804), .A3(new_n838), .ZN(G150));
  NAND2_X1  g415(.A1(new_n630), .A2(G559), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT103), .Z(new_n842));
  INV_X1    g417(.A(KEYINPUT38), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n841), .B(KEYINPUT103), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(KEYINPUT38), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n538), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n848), .A2(new_n529), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n532), .A2(G55), .ZN(new_n850));
  INV_X1    g425(.A(G93), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n850), .B1(new_n541), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n569), .A2(new_n854), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n562), .B(new_n853), .C1(new_n567), .C2(new_n568), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n847), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n857), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n844), .A2(new_n859), .A3(new_n846), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(KEYINPUT39), .A3(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT104), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n858), .A2(KEYINPUT104), .A3(KEYINPUT39), .A4(new_n860), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(KEYINPUT39), .B1(new_n858), .B2(new_n860), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n866), .A2(G860), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n854), .A2(G860), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(KEYINPUT37), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(G145));
  NAND2_X1  g446(.A1(new_n789), .A2(KEYINPUT105), .ZN(new_n872));
  AOI211_X1 g447(.A(new_n494), .B(G2105), .C1(new_n466), .C2(new_n468), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n498), .B(new_n499), .C1(new_n873), .C2(new_n501), .ZN(new_n874));
  INV_X1    g449(.A(G126), .ZN(new_n875));
  AOI211_X1 g450(.A(new_n875), .B(new_n460), .C1(new_n466), .C2(new_n468), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n876), .B1(new_n521), .B2(new_n522), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n872), .B(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n490), .A2(G130), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n460), .A2(G118), .ZN(new_n881));
  OAI21_X1  g456(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n883), .B1(new_n482), .B2(G142), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n653), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n879), .B(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n767), .B(new_n744), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n825), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n886), .A2(new_n888), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(G162), .B(new_n649), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(G160), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(G37), .ZN(new_n896));
  INV_X1    g471(.A(new_n891), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n897), .A2(new_n894), .A3(new_n889), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n895), .A2(KEYINPUT40), .A3(new_n896), .A4(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n896), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n892), .A2(new_n894), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n899), .A2(new_n903), .ZN(G395));
  NOR2_X1   g479(.A1(new_n854), .A2(G868), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n642), .A2(new_n857), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n641), .A2(new_n859), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n633), .B(new_n629), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT41), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n908), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n908), .B2(new_n911), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n906), .A2(new_n909), .A3(new_n907), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT106), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT109), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n916), .B(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n920), .B(new_n921), .C1(new_n914), .C2(new_n913), .ZN(new_n922));
  XNOR2_X1  g497(.A(G290), .B(new_n593), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g500(.A(G166), .B(G305), .Z(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n924), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g505(.A(new_n930), .B(KEYINPUT42), .Z(new_n931));
  NAND3_X1  g506(.A1(new_n918), .A2(new_n922), .A3(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n915), .A2(new_n917), .ZN(new_n933));
  INV_X1    g508(.A(new_n931), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n921), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n905), .B1(new_n936), .B2(G868), .ZN(G295));
  AOI21_X1  g512(.A(new_n905), .B1(new_n936), .B2(G868), .ZN(G331));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n939));
  INV_X1    g514(.A(new_n930), .ZN(new_n940));
  NOR2_X1   g515(.A1(G171), .A2(KEYINPUT110), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n859), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(G286), .B1(KEYINPUT110), .B2(G171), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n942), .B1(new_n855), .B2(new_n856), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n944), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n857), .A2(new_n941), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n948), .B1(new_n949), .B2(new_n945), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n911), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n947), .A2(new_n950), .A3(new_n909), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n940), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT111), .B1(new_n954), .B2(G37), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n952), .A2(new_n940), .A3(new_n953), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n947), .A2(new_n950), .A3(new_n909), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n910), .B1(new_n947), .B2(new_n950), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n930), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT111), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(new_n962), .A3(new_n896), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n955), .A2(new_n958), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n961), .A2(new_n956), .A3(new_n896), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n939), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n955), .A2(new_n963), .A3(new_n956), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n954), .A2(G37), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n968), .A2(KEYINPUT43), .B1(new_n969), .B2(new_n958), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n967), .B1(new_n970), .B2(new_n939), .ZN(G397));
  AOI211_X1 g546(.A(KEYINPUT75), .B(new_n876), .C1(new_n521), .C2(new_n522), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n524), .B1(new_n523), .B2(new_n504), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n874), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n975));
  INV_X1    g550(.A(G1384), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G40), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n472), .A2(new_n476), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n878), .A2(new_n976), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n980), .B1(new_n981), .B2(KEYINPUT50), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n977), .A2(new_n799), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(G164), .B2(G1384), .ZN(new_n985));
  AOI21_X1  g560(.A(G1384), .B1(new_n874), .B2(new_n877), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n980), .B1(new_n986), .B2(KEYINPUT45), .ZN(new_n987));
  AOI21_X1  g562(.A(G1971), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT119), .B1(new_n983), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT119), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n977), .A2(new_n982), .A3(new_n799), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n878), .A2(KEYINPUT45), .A3(new_n976), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n979), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n974), .A2(new_n976), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n993), .B1(new_n994), .B2(new_n984), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n990), .B(new_n991), .C1(new_n995), .C2(G1971), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n989), .A2(G8), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G8), .ZN(new_n998));
  NOR2_X1   g573(.A1(G166), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n997), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n998), .B1(new_n986), .B2(new_n979), .ZN(new_n1003));
  INV_X1    g578(.A(G1976), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n593), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n594), .A2(new_n597), .A3(new_n1004), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1008), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n581), .A2(G86), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n613), .A2(new_n1013), .A3(new_n604), .A4(new_n605), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(G1981), .ZN(new_n1015));
  INV_X1    g590(.A(G1981), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n606), .A2(new_n611), .A3(new_n1016), .A4(new_n613), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1015), .A2(new_n1017), .A3(KEYINPUT49), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT116), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1015), .A2(new_n1017), .A3(new_n1020), .A4(KEYINPUT49), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1003), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT49), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1012), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n985), .A2(new_n987), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n807), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n986), .A2(new_n1030), .A3(new_n975), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1031), .A2(new_n979), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n878), .A2(new_n975), .A3(new_n976), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT114), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1032), .A2(new_n799), .A3(new_n1033), .A4(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n998), .B1(new_n1029), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1001), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1027), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1032), .A2(new_n731), .A3(new_n1033), .A4(new_n1035), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n974), .A2(KEYINPUT45), .A3(new_n976), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n980), .B1(new_n981), .B2(new_n984), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1966), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1040), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(G8), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1047), .A2(G286), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1002), .A2(new_n1039), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT63), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI211_X1 g626(.A(new_n998), .B(new_n1001), .C1(new_n1029), .C2(new_n1036), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(new_n1050), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1006), .A2(KEYINPUT52), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1054), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1012), .A2(new_n1026), .A3(KEYINPUT117), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1053), .A2(new_n1060), .A3(new_n1048), .A4(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1035), .A2(new_n979), .A3(new_n1031), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n975), .B1(new_n974), .B2(new_n976), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1064), .A2(new_n1065), .A3(G2090), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1038), .B(G8), .C1(new_n1066), .C2(new_n988), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1067), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1026), .A2(new_n1004), .A3(new_n598), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1023), .B1(new_n1069), .B2(new_n1017), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1063), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1012), .A2(new_n1026), .A3(KEYINPUT117), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT117), .B1(new_n1012), .B2(new_n1026), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1052), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1070), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(new_n1075), .A3(KEYINPUT118), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1051), .A2(new_n1062), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(G168), .A2(new_n998), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1047), .B(new_n1079), .C1(KEYINPUT122), .C2(KEYINPUT51), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT51), .B1(new_n1079), .B2(KEYINPUT122), .ZN(new_n1081));
  OAI211_X1 g656(.A(G8), .B(new_n1081), .C1(new_n1046), .C2(G286), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1046), .A2(new_n1078), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1080), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT62), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1086));
  INV_X1    g661(.A(G2078), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n985), .A2(new_n1087), .A3(new_n987), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1086), .A2(new_n720), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1089), .A2(G2078), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1041), .A2(new_n1042), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(G301), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1002), .A2(new_n1039), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT62), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1080), .A2(new_n1082), .A3(new_n1095), .A4(new_n1083), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1085), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G1956), .ZN(new_n1098));
  NOR3_X1   g673(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n979), .B1(new_n986), .B2(new_n975), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT56), .B(G2072), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n985), .A2(new_n987), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  OR2_X1    g679(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n1105));
  NAND2_X1  g680(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n633), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(G299), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1104), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1064), .ZN(new_n1111));
  AOI21_X1  g686(.A(G1348), .B1(new_n1111), .B2(new_n1033), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n986), .A2(new_n979), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1113), .A2(G2067), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n630), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1109), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1101), .A2(new_n1116), .A3(new_n1103), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1110), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G1996), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n985), .A2(new_n1119), .A3(new_n987), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT58), .B(G1341), .Z(new_n1121));
  NAND2_X1  g696(.A1(new_n1113), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n569), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1123), .B(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1101), .A2(new_n1116), .A3(new_n1103), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1110), .A2(KEYINPUT61), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1116), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1128), .B1(new_n1117), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1125), .A2(new_n1127), .A3(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n1132));
  INV_X1    g707(.A(new_n630), .ZN(new_n1133));
  INV_X1    g708(.A(G1348), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1114), .B1(new_n1086), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT60), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1133), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1132), .B1(new_n1137), .B2(new_n1115), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1131), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1137), .A2(new_n1115), .A3(new_n1132), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1118), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1090), .A2(G301), .A3(new_n1092), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n981), .A2(new_n984), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n979), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n992), .A2(new_n1091), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT124), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1042), .A2(new_n1147), .A3(new_n992), .A4(new_n1091), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  AOI211_X1 g724(.A(KEYINPUT125), .B(G301), .C1(new_n1090), .C2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT125), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1086), .A2(new_n720), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1152), .A2(new_n1149), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1151), .B1(new_n1154), .B2(G171), .ZN(new_n1155));
  OAI211_X1 g730(.A(KEYINPUT54), .B(new_n1142), .C1(new_n1150), .C2(new_n1155), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1002), .A2(new_n1039), .ZN(new_n1157));
  XNOR2_X1  g732(.A(KEYINPUT123), .B(KEYINPUT54), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1154), .A2(G171), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1158), .B1(new_n1159), .B2(new_n1093), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1156), .A2(new_n1157), .A3(new_n1084), .A4(new_n1160), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1077), .B(new_n1097), .C1(new_n1141), .C2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1143), .A2(new_n980), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n1119), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1164), .A2(new_n744), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n1165), .B(KEYINPUT112), .Z(new_n1166));
  XNOR2_X1  g741(.A(new_n767), .B(G2067), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n1163), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT113), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1163), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1170), .A2(new_n1119), .A3(new_n745), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1166), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n825), .A2(new_n828), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n825), .A2(new_n828), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1163), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(G290), .B(G1986), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1176), .B1(new_n1163), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1162), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT46), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1164), .A2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(KEYINPUT126), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n745), .B1(new_n1180), .B2(G1996), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1163), .B1(new_n1167), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(KEYINPUT47), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1170), .A2(G1986), .A3(G290), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1187), .B(KEYINPUT48), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1186), .B1(new_n1176), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1190));
  OR2_X1    g765(.A1(new_n767), .A2(G2067), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1170), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1179), .A2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g769(.A1(new_n689), .A2(G319), .A3(new_n690), .ZN(new_n1196));
  XOR2_X1   g770(.A(new_n1196), .B(KEYINPUT127), .Z(new_n1197));
  NAND2_X1  g771(.A1(new_n1197), .A2(new_n672), .ZN(new_n1198));
  AOI21_X1  g772(.A(new_n1198), .B1(new_n710), .B2(new_n711), .ZN(new_n1199));
  OAI21_X1  g773(.A(new_n1199), .B1(new_n901), .B2(new_n902), .ZN(new_n1200));
  NOR2_X1   g774(.A1(new_n1200), .A2(new_n970), .ZN(G308));
  NAND3_X1  g775(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n1202));
  AND2_X1   g776(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n1203));
  AND2_X1   g777(.A1(new_n958), .A2(new_n969), .ZN(new_n1204));
  OAI211_X1 g778(.A(new_n1202), .B(new_n1199), .C1(new_n1203), .C2(new_n1204), .ZN(G225));
endmodule


