//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056;
  INV_X1    g000(.A(KEYINPUT78), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT71), .B(G217), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n189), .B1(G234), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT76), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT25), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G125), .ZN(new_n196));
  INV_X1    g010(.A(G125), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G140), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n198), .A3(KEYINPUT74), .ZN(new_n199));
  OR3_X1    g013(.A1(new_n197), .A2(KEYINPUT74), .A3(G140), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(KEYINPUT16), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT16), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n196), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n201), .A2(new_n206), .A3(new_n203), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(KEYINPUT75), .A3(new_n207), .ZN(new_n208));
  AOI211_X1 g022(.A(KEYINPUT75), .B(new_n206), .C1(new_n201), .C2(new_n203), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G119), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G128), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(KEYINPUT73), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(G128), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT23), .ZN(new_n215));
  OR2_X1    g029(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n216));
  AOI22_X1  g030(.A1(new_n213), .A2(new_n215), .B1(new_n212), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G110), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OR3_X1    g033(.A1(new_n211), .A2(KEYINPUT72), .A3(G128), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT72), .B1(new_n211), .B2(G128), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(new_n214), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT24), .B(G110), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n208), .A2(new_n210), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n217), .A2(new_n218), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n222), .A2(new_n223), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n196), .A2(new_n198), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n206), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n205), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT22), .B(G137), .ZN(new_n233));
  INV_X1    g047(.A(G221), .ZN(new_n234));
  INV_X1    g048(.A(G234), .ZN(new_n235));
  NOR3_X1   g049(.A1(new_n234), .A2(new_n235), .A3(G953), .ZN(new_n236));
  XOR2_X1   g050(.A(new_n233), .B(new_n236), .Z(new_n237));
  AND3_X1   g051(.A1(new_n226), .A2(new_n232), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n237), .B1(new_n226), .B2(new_n232), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(G902), .B1(new_n192), .B2(new_n193), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n194), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n226), .A2(new_n232), .ZN(new_n243));
  INV_X1    g057(.A(new_n237), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n226), .A2(new_n232), .A3(new_n237), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n245), .A2(new_n246), .A3(new_n241), .A4(new_n194), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n191), .B1(new_n242), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n191), .A2(G902), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT77), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n252), .B1(new_n238), .B2(new_n239), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n245), .A2(KEYINPUT77), .A3(new_n246), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n251), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n187), .B1(new_n249), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n191), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n245), .A2(new_n246), .A3(new_n241), .ZN(new_n259));
  INV_X1    g073(.A(new_n194), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n258), .B1(new_n261), .B2(new_n247), .ZN(new_n262));
  NOR3_X1   g076(.A1(new_n262), .A2(KEYINPUT78), .A3(new_n255), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G113), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT2), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT2), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G113), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(G116), .B(G119), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n269), .B1(new_n270), .B2(KEYINPUT67), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n211), .A2(G116), .ZN(new_n272));
  INV_X1    g086(.A(G116), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G119), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT2), .B(G113), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT67), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n271), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(KEYINPUT66), .A2(KEYINPUT30), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT66), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT30), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G128), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(KEYINPUT1), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n206), .A2(G143), .ZN(new_n287));
  INV_X1    g101(.A(G143), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G146), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n286), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT65), .ZN(new_n291));
  XNOR2_X1  g105(.A(G143), .B(G146), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT65), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n293), .A3(new_n286), .ZN(new_n294));
  INV_X1    g108(.A(new_n292), .ZN(new_n295));
  OAI21_X1  g109(.A(KEYINPUT1), .B1(new_n288), .B2(G146), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G128), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n291), .A2(new_n294), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G134), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT11), .B1(new_n299), .B2(G137), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT11), .ZN(new_n301));
  INV_X1    g115(.A(G137), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n302), .A3(G134), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G131), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n302), .A2(G134), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT64), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n309), .B1(new_n302), .B2(G134), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n302), .A2(G134), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n299), .A2(KEYINPUT64), .A3(G137), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G131), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n298), .A2(new_n315), .ZN(new_n316));
  AND2_X1   g130(.A1(KEYINPUT0), .A2(G128), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n287), .A2(new_n289), .A3(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT0), .B(G128), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n318), .B1(new_n292), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n304), .A2(new_n307), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G131), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n320), .B1(new_n322), .B2(new_n308), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n281), .B(new_n284), .C1(new_n316), .C2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n295), .A2(new_n297), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n293), .B1(new_n292), .B2(new_n286), .ZN(new_n326));
  AND4_X1   g140(.A1(new_n293), .A2(new_n286), .A3(new_n287), .A4(new_n289), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(new_n308), .A3(new_n314), .ZN(new_n329));
  INV_X1    g143(.A(new_n320), .ZN(new_n330));
  INV_X1    g144(.A(new_n308), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n305), .B1(new_n304), .B2(new_n307), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n329), .A2(new_n282), .A3(new_n333), .A4(new_n283), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n280), .B1(new_n324), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT31), .ZN(new_n336));
  NOR2_X1   g150(.A1(G237), .A2(G953), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G210), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(KEYINPUT27), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT26), .B(G101), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n339), .B(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n316), .A2(new_n323), .A3(new_n279), .ZN(new_n343));
  NOR4_X1   g157(.A1(new_n335), .A2(new_n336), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(G472), .A2(G902), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n346), .A2(KEYINPUT32), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n324), .A2(new_n334), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n279), .ZN(new_n349));
  INV_X1    g163(.A(new_n343), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n341), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n336), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT68), .B1(new_n316), .B2(new_n323), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT68), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n329), .A2(new_n354), .A3(new_n333), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(new_n355), .A3(new_n280), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT28), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n280), .B1(new_n329), .B2(new_n333), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT28), .B1(new_n343), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n341), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n345), .B(new_n347), .C1(new_n352), .C2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT70), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n345), .B(new_n346), .C1(new_n352), .C2(new_n361), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT69), .B(KEYINPUT32), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n329), .A2(new_n333), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n279), .B1(new_n368), .B2(KEYINPUT68), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT28), .B1(new_n369), .B2(new_n355), .ZN(new_n370));
  INV_X1    g184(.A(new_n359), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n357), .B1(new_n350), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n342), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n343), .B1(new_n348), .B2(new_n279), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT31), .B1(new_n374), .B2(new_n341), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n344), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(KEYINPUT70), .A3(new_n347), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n358), .A2(new_n341), .A3(new_n360), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT29), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n342), .B1(new_n335), .B2(new_n343), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n190), .B1(new_n378), .B2(new_n379), .ZN(new_n382));
  OAI21_X1  g196(.A(G472), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n364), .A2(new_n367), .A3(new_n377), .A4(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT9), .B(G234), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n234), .B1(new_n386), .B2(new_n190), .ZN(new_n387));
  INV_X1    g201(.A(G469), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(new_n190), .ZN(new_n389));
  INV_X1    g203(.A(G104), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT3), .B1(new_n390), .B2(G107), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT3), .ZN(new_n392));
  INV_X1    g206(.A(G107), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(G104), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n390), .A2(G107), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n391), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(G101), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT80), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT80), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n396), .A2(new_n400), .A3(new_n397), .A4(G101), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n397), .B1(new_n396), .B2(G101), .ZN(new_n403));
  INV_X1    g217(.A(G101), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n391), .A2(new_n394), .A3(new_n404), .A4(new_n395), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n320), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT10), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n296), .A2(KEYINPUT81), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT81), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n410), .B(KEYINPUT1), .C1(new_n288), .C2(G146), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(G128), .A3(new_n411), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n412), .A2(new_n295), .B1(new_n291), .B2(new_n294), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n390), .A2(G107), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n393), .A2(G104), .ZN(new_n415));
  OAI21_X1  g229(.A(G101), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n405), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n408), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n405), .A2(new_n416), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n328), .A2(KEYINPUT10), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n407), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n322), .A2(new_n308), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n422), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n407), .A2(new_n418), .A3(new_n424), .A4(new_n420), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G953), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G227), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(KEYINPUT79), .ZN(new_n429));
  XNOR2_X1  g243(.A(G110), .B(G140), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n429), .B(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n426), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n291), .A2(new_n294), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n434), .A2(new_n325), .A3(new_n417), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n411), .A2(G128), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n410), .B1(new_n287), .B2(KEYINPUT1), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n295), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n417), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(KEYINPUT12), .B(new_n422), .C1(new_n435), .C2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n434), .A2(new_n325), .A3(new_n417), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(new_n413), .B2(new_n417), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT12), .B1(new_n443), .B2(new_n422), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n425), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT82), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT82), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n447), .B(new_n425), .C1(new_n441), .C2(new_n444), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n433), .B1(new_n449), .B2(new_n432), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n389), .B1(new_n450), .B2(G469), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n431), .B(new_n425), .C1(new_n441), .C2(new_n444), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT83), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n426), .A2(new_n432), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n422), .B1(new_n435), .B2(new_n439), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT12), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n440), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n459), .A2(KEYINPUT83), .A3(new_n431), .A4(new_n425), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n454), .A2(new_n455), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n388), .A3(new_n190), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n387), .B1(new_n451), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G952), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n464), .A2(KEYINPUT89), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n464), .A2(KEYINPUT89), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n427), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n467), .B1(G234), .B2(G237), .ZN(new_n468));
  NAND2_X1  g282(.A1(G234), .A2(G237), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(G902), .A3(G953), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT90), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT21), .B(G898), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n468), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(G214), .B1(G237), .B2(G902), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n320), .A2(G125), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT84), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n434), .A2(new_n197), .A3(new_n325), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT84), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n320), .A2(new_n479), .A3(G125), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n477), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G224), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(G953), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT7), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n483), .B1(KEYINPUT85), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(KEYINPUT85), .B2(new_n484), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n273), .A2(G119), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT5), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n265), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n272), .A2(new_n274), .A3(KEYINPUT5), .ZN(new_n490));
  AOI22_X1  g304(.A1(new_n489), .A2(new_n490), .B1(new_n269), .B2(new_n270), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n419), .A2(new_n491), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n272), .A2(new_n274), .A3(KEYINPUT5), .ZN(new_n493));
  OAI21_X1  g307(.A(G113), .B1(new_n272), .B2(KEYINPUT5), .ZN(new_n494));
  OAI22_X1  g308(.A1(new_n493), .A2(new_n494), .B1(new_n275), .B2(new_n276), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n417), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(G110), .B(G122), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(KEYINPUT8), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n481), .A2(new_n486), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n495), .A2(new_n417), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n403), .A2(new_n405), .B1(new_n278), .B2(new_n271), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n501), .B1(new_n402), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n498), .ZN(new_n504));
  INV_X1    g318(.A(new_n480), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n479), .B1(new_n320), .B2(G125), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n483), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n507), .A2(KEYINPUT7), .A3(new_n508), .A4(new_n478), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n500), .A2(new_n504), .A3(new_n509), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n510), .A2(new_n190), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT6), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(new_n503), .B2(new_n498), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n402), .A2(new_n502), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n492), .ZN(new_n515));
  INV_X1    g329(.A(new_n498), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n481), .B(new_n483), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n515), .A2(new_n512), .A3(new_n516), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(G210), .B1(G237), .B2(G902), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n511), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n522), .B1(new_n511), .B2(new_n521), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n474), .B(new_n475), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(G113), .B(G122), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(new_n390), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n337), .A2(G143), .A3(G214), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(G143), .B1(new_n337), .B2(G214), .ZN(new_n530));
  OAI21_X1  g344(.A(G131), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n530), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(new_n305), .A3(new_n528), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n230), .A2(KEYINPUT19), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n199), .A2(new_n200), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n535), .B1(new_n536), .B2(KEYINPUT19), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n205), .B(new_n534), .C1(new_n537), .C2(G146), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n532), .A2(new_n528), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(KEYINPUT18), .A3(G131), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n231), .B1(new_n536), .B2(new_n206), .ZN(new_n541));
  NAND2_X1  g355(.A1(KEYINPUT18), .A2(G131), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n532), .A2(new_n528), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n527), .B1(new_n538), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n544), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n208), .A2(new_n210), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n531), .A2(new_n533), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n539), .A2(KEYINPUT17), .A3(G131), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n546), .B1(new_n547), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n545), .B1(new_n553), .B2(new_n527), .ZN(new_n554));
  NOR2_X1   g368(.A1(G475), .A2(G902), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT20), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n207), .A2(KEYINPUT75), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n206), .B1(new_n201), .B2(new_n203), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n552), .B1(new_n560), .B2(new_n209), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(new_n527), .A3(new_n544), .ZN(new_n562));
  INV_X1    g376(.A(new_n545), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT20), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n565), .A3(new_n555), .ZN(new_n566));
  INV_X1    g380(.A(new_n527), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n551), .B1(new_n208), .B2(new_n210), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n567), .B1(new_n568), .B2(new_n546), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n562), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n190), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n557), .A2(new_n566), .B1(new_n571), .B2(G475), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n288), .A2(KEYINPUT13), .A3(G128), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT13), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(new_n285), .B2(G143), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n285), .A2(G143), .ZN(new_n576));
  OAI211_X1 g390(.A(KEYINPUT86), .B(new_n573), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT86), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n288), .A2(G128), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n288), .A2(G128), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n578), .B(new_n579), .C1(new_n580), .C2(new_n574), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n577), .A2(G134), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT87), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n577), .A2(KEYINPUT87), .A3(G134), .A4(new_n581), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n576), .A2(new_n580), .A3(G134), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  OR2_X1    g402(.A1(new_n273), .A2(G122), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n273), .A2(G122), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n590), .A3(new_n393), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n393), .B1(new_n589), .B2(new_n590), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n588), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n586), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n285), .A2(G143), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n299), .B1(new_n579), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n591), .B1(new_n587), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT14), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(new_n273), .A3(G122), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n600), .B1(new_n273), .B2(G122), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT88), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n602), .A2(KEYINPUT88), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n589), .B(new_n601), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n599), .B1(new_n606), .B2(G107), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n386), .A2(new_n427), .A3(new_n188), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n596), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n594), .B1(new_n584), .B2(new_n585), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n609), .B1(new_n612), .B2(new_n607), .ZN(new_n613));
  AOI21_X1  g427(.A(G902), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(G478), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(KEYINPUT15), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n614), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n572), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n525), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n264), .A2(new_n384), .A3(new_n463), .A4(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G101), .ZN(G3));
  AOI21_X1  g435(.A(new_n565), .B1(new_n564), .B2(new_n555), .ZN(new_n622));
  AOI211_X1 g436(.A(KEYINPUT20), .B(new_n556), .C1(new_n562), .C2(new_n563), .ZN(new_n623));
  INV_X1    g437(.A(G475), .ZN(new_n624));
  AOI21_X1  g438(.A(G902), .B1(new_n562), .B2(new_n569), .ZN(new_n625));
  OAI22_X1  g439(.A1(new_n622), .A2(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n615), .A2(new_n190), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n614), .B2(new_n615), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n611), .A2(new_n613), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT91), .B1(new_n612), .B2(new_n607), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(KEYINPUT33), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n611), .A2(new_n613), .A3(new_n631), .A4(KEYINPUT33), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n615), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n629), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n626), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n525), .A2(new_n637), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n345), .B(new_n190), .C1(new_n352), .C2(new_n361), .ZN(new_n639));
  AOI22_X1  g453(.A1(new_n639), .A2(G472), .B1(new_n376), .B2(new_n346), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n264), .A2(new_n463), .A3(new_n638), .A4(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  INV_X1    g457(.A(KEYINPUT92), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n644), .B1(new_n622), .B2(new_n623), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n571), .A2(G475), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n557), .A2(new_n566), .A3(KEYINPUT92), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n610), .B1(new_n596), .B2(new_n608), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n612), .A2(new_n607), .A3(new_n609), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n190), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n616), .ZN(new_n651));
  INV_X1    g465(.A(new_n616), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n614), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n645), .A2(new_n646), .A3(new_n647), .A4(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n525), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n264), .A2(new_n463), .A3(new_n656), .A4(new_n640), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT94), .B(G107), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT93), .B(KEYINPUT35), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G9));
  NOR2_X1   g475(.A1(new_n244), .A2(KEYINPUT36), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n243), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n250), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n249), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n463), .A2(new_n619), .A3(new_n640), .A4(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT37), .B(G110), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  INV_X1    g482(.A(G900), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n468), .B1(new_n669), .B2(new_n471), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n655), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n664), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n262), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n475), .B1(new_n523), .B2(new_n524), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n384), .A2(new_n463), .A3(new_n671), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  NOR2_X1   g491(.A1(new_n523), .A2(new_n524), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT38), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n557), .A2(new_n566), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n617), .B1(new_n680), .B2(new_n646), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n673), .A2(new_n475), .A3(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT40), .ZN(new_n684));
  INV_X1    g498(.A(new_n448), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n447), .B1(new_n459), .B2(new_n425), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n432), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n433), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n687), .A2(G469), .A3(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n389), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n689), .A2(new_n462), .A3(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n387), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n670), .B(KEYINPUT39), .Z(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n683), .B1(new_n684), .B2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT96), .ZN(new_n699));
  INV_X1    g513(.A(new_n374), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n341), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n350), .A2(new_n371), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n190), .B1(new_n703), .B2(new_n341), .ZN(new_n704));
  OAI21_X1  g518(.A(G472), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n364), .A2(new_n367), .A3(new_n377), .A4(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT95), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n696), .A2(new_n684), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n698), .A2(new_n699), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  OAI21_X1  g527(.A(KEYINPUT96), .B1(new_n713), .B2(new_n697), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(new_n288), .ZN(G45));
  INV_X1    g530(.A(new_n634), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n611), .A2(new_n613), .B1(new_n631), .B2(KEYINPUT33), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n628), .B1(new_n719), .B2(new_n615), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n572), .A2(new_n720), .A3(new_n670), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n384), .A2(new_n463), .A3(new_n675), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G146), .ZN(G48));
  NAND2_X1  g537(.A1(new_n461), .A2(new_n190), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(G469), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n725), .A2(new_n692), .A3(new_n462), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n264), .A2(new_n384), .A3(new_n638), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT41), .B(G113), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(KEYINPUT97), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n727), .B(new_n729), .ZN(G15));
  NAND4_X1  g544(.A1(new_n264), .A2(new_n384), .A3(new_n656), .A4(new_n726), .ZN(new_n731));
  XOR2_X1   g545(.A(KEYINPUT98), .B(G116), .Z(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G18));
  NOR2_X1   g547(.A1(new_n618), .A2(new_n473), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n384), .A2(new_n726), .A3(new_n675), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G119), .ZN(G21));
  NAND2_X1  g550(.A1(new_n626), .A2(new_n654), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n674), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n726), .A2(new_n474), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n262), .A2(new_n255), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n639), .A2(G472), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n346), .B(KEYINPUT99), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n345), .B(new_n742), .C1(new_n352), .C2(new_n361), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT100), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n376), .A2(KEYINPUT100), .A3(new_n742), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n740), .A2(new_n741), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT101), .B1(new_n739), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n475), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n511), .A2(new_n521), .ZN(new_n750));
  INV_X1    g564(.A(new_n522), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n511), .A2(new_n521), .A3(new_n522), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n749), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n681), .A3(new_n474), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n725), .A2(new_n692), .A3(new_n462), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AND4_X1   g571(.A1(new_n740), .A2(new_n741), .A3(new_n745), .A4(new_n746), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT101), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n748), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G122), .ZN(G24));
  AND4_X1   g576(.A1(new_n741), .A2(new_n665), .A3(new_n745), .A4(new_n746), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n756), .A2(new_n674), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n764), .A3(new_n721), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G125), .ZN(G27));
  NOR3_X1   g580(.A1(new_n523), .A2(new_n524), .A3(new_n749), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n383), .A2(new_n362), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT32), .B1(new_n376), .B2(new_n346), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n740), .B(new_n767), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n721), .A2(new_n692), .A3(new_n691), .ZN(new_n771));
  OAI21_X1  g585(.A(KEYINPUT42), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n691), .A2(new_n692), .A3(new_n767), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n637), .A2(KEYINPUT42), .A3(new_n670), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n773), .A2(new_n264), .A3(new_n384), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n305), .ZN(G33));
  NAND4_X1  g591(.A1(new_n773), .A2(new_n264), .A3(new_n384), .A4(new_n671), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G134), .ZN(G36));
  INV_X1    g593(.A(KEYINPUT46), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n389), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n687), .A2(new_n688), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n388), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n687), .A2(KEYINPUT45), .A3(new_n688), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT102), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n431), .B1(new_n446), .B2(new_n448), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n783), .B1(new_n787), .B2(new_n433), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n788), .A2(new_n785), .A3(KEYINPUT102), .A4(G469), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n781), .B1(new_n786), .B2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT103), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n792), .A3(new_n462), .ZN(new_n793));
  INV_X1    g607(.A(new_n781), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n788), .A2(new_n785), .A3(G469), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT102), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n794), .B1(new_n797), .B2(new_n789), .ZN(new_n798));
  INV_X1    g612(.A(new_n462), .ZN(new_n799));
  OAI21_X1  g613(.A(KEYINPUT103), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n690), .B1(new_n786), .B2(new_n790), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n780), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n793), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n692), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n572), .A2(new_n636), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT43), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n805), .B(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n640), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(new_n808), .A3(new_n665), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT44), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n807), .A2(KEYINPUT44), .A3(new_n808), .A4(new_n665), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n767), .A3(new_n812), .ZN(new_n813));
  OR3_X1    g627(.A1(new_n804), .A2(new_n695), .A3(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G137), .ZN(G39));
  NAND2_X1  g629(.A1(new_n721), .A2(new_n767), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n264), .A2(new_n816), .A3(new_n384), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n803), .A2(KEYINPUT47), .A3(new_n692), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT47), .B1(new_n803), .B2(new_n692), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G140), .ZN(G42));
  NAND2_X1  g635(.A1(new_n807), .A2(new_n468), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n747), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n679), .A2(new_n749), .A3(new_n726), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n823), .A2(KEYINPUT50), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT50), .B1(new_n823), .B2(new_n824), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n710), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n264), .A2(new_n468), .A3(new_n726), .A4(new_n767), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n626), .A2(new_n636), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n726), .A2(new_n767), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n822), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n763), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n827), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n725), .A2(new_n462), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n387), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n818), .A2(new_n819), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n823), .A2(new_n767), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n837), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n740), .B1(new_n768), .B2(new_n769), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n822), .A2(new_n844), .A3(new_n832), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n845), .B(KEYINPUT48), .Z(new_n846));
  NAND4_X1  g660(.A1(new_n828), .A2(new_n626), .A3(new_n636), .A4(new_n829), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n467), .B1(new_n823), .B2(new_n764), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n843), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT47), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n804), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n803), .A2(KEYINPUT47), .A3(new_n692), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n839), .B(KEYINPUT114), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n842), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n827), .A2(new_n835), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT51), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT115), .B1(new_n851), .B2(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n384), .A2(new_n675), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n693), .A2(new_n655), .A3(new_n670), .ZN(new_n863));
  INV_X1    g677(.A(new_n771), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT52), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n670), .B(KEYINPUT111), .Z(new_n867));
  NOR2_X1   g681(.A1(new_n665), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n706), .A2(new_n463), .A3(new_n738), .A4(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n865), .A2(new_n866), .A3(new_n765), .A4(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n645), .A2(new_n647), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT109), .ZN(new_n872));
  INV_X1    g686(.A(new_n670), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n651), .A2(new_n653), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n625), .A2(new_n624), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n871), .A2(new_n872), .A3(new_n767), .A4(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n645), .A3(new_n647), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n752), .A2(new_n475), .A3(new_n753), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT109), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n384), .A2(new_n463), .A3(new_n665), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n778), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(new_n776), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n765), .A2(new_n676), .A3(new_n722), .A4(new_n869), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT52), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n763), .A2(new_n773), .A3(new_n721), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT110), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n763), .A2(new_n773), .A3(KEYINPUT110), .A4(new_n721), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AND4_X1   g705(.A1(new_n870), .A2(new_n884), .A3(new_n886), .A4(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n759), .B1(new_n757), .B2(new_n758), .ZN(new_n893));
  NOR4_X1   g707(.A1(new_n747), .A2(new_n755), .A3(new_n756), .A4(KEYINPUT101), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n731), .A2(new_n727), .A3(new_n735), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n895), .A2(KEYINPUT106), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT106), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n731), .A2(new_n727), .A3(new_n735), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n898), .B1(new_n899), .B2(new_n761), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n620), .A2(new_n641), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT107), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT107), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n620), .A2(new_n641), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n572), .A2(new_n654), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n525), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n264), .A2(new_n463), .A3(new_n640), .A4(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n666), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT108), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n909), .A2(KEYINPUT108), .A3(new_n666), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n906), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n892), .A2(new_n901), .A3(KEYINPUT53), .A4(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT53), .ZN(new_n917));
  OAI21_X1  g731(.A(KEYINPUT106), .B1(new_n895), .B2(new_n896), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n899), .A2(new_n761), .A3(new_n898), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n918), .A2(new_n919), .A3(new_n906), .A4(new_n914), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n884), .A2(new_n886), .A3(new_n870), .A4(new_n891), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n916), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT54), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT113), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT112), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n895), .B2(new_n896), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n899), .A2(new_n761), .A3(KEYINPUT112), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n927), .A2(KEYINPUT53), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(new_n892), .A3(new_n915), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT54), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n930), .A2(new_n922), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n924), .A2(new_n925), .A3(new_n932), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n930), .A2(new_n922), .A3(new_n931), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n931), .B1(new_n916), .B2(new_n922), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT113), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n855), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n818), .A2(new_n819), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n859), .B1(new_n938), .B2(new_n842), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n836), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT115), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n853), .A2(new_n854), .A3(new_n839), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n857), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n849), .B1(new_n943), .B2(new_n837), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n940), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n861), .A2(new_n933), .A3(new_n936), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n464), .A2(new_n427), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n740), .A2(new_n692), .A3(new_n475), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n949), .A2(new_n805), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT104), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n828), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT49), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n679), .B1(new_n953), .B2(new_n838), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT105), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n838), .A2(new_n953), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n952), .B(new_n957), .C1(new_n955), .C2(new_n956), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n948), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT116), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n948), .A2(KEYINPUT116), .A3(new_n958), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(G75));
  NOR2_X1   g777(.A1(new_n427), .A2(G952), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n190), .B1(new_n930), .B2(new_n922), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT56), .B1(new_n966), .B2(G210), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n518), .A2(new_n520), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(new_n519), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT55), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n965), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n967), .B2(new_n970), .ZN(G51));
  AOI21_X1  g786(.A(new_n931), .B1(new_n930), .B2(new_n922), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n934), .A2(new_n973), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n389), .B(KEYINPUT57), .Z(new_n975));
  OAI21_X1  g789(.A(new_n461), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n966), .A2(new_n797), .A3(new_n789), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n964), .B1(new_n976), .B2(new_n977), .ZN(G54));
  NAND3_X1  g792(.A1(new_n966), .A2(KEYINPUT58), .A3(G475), .ZN(new_n979));
  OR3_X1    g793(.A1(new_n979), .A2(KEYINPUT117), .A3(new_n554), .ZN(new_n980));
  OAI21_X1  g794(.A(KEYINPUT117), .B1(new_n979), .B2(new_n554), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n964), .B1(new_n979), .B2(new_n554), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(G60));
  XOR2_X1   g797(.A(new_n627), .B(KEYINPUT59), .Z(new_n984));
  NAND2_X1  g798(.A1(new_n719), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n965), .B1(new_n974), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT118), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n933), .A2(new_n936), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n719), .B1(new_n988), .B2(new_n984), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n987), .A2(new_n989), .ZN(G63));
  NAND2_X1  g804(.A1(G217), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT119), .Z(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT60), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n993), .B1(new_n930), .B2(new_n922), .ZN(new_n994));
  INV_X1    g808(.A(new_n253), .ZN(new_n995));
  INV_X1    g809(.A(new_n254), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n965), .B1(new_n994), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n999), .B1(new_n663), .B2(new_n994), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT61), .ZN(G66));
  OAI21_X1  g815(.A(G953), .B1(new_n472), .B2(new_n482), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT120), .ZN(new_n1003));
  INV_X1    g817(.A(new_n920), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1003), .B1(new_n1004), .B2(G953), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n968), .B1(G898), .B2(new_n427), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1005), .B(new_n1006), .ZN(G69));
  XNOR2_X1  g821(.A(new_n348), .B(KEYINPUT121), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(new_n537), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n879), .B1(new_n637), .B2(new_n907), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n696), .A2(new_n384), .A3(new_n264), .A4(new_n1010), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n814), .A2(new_n1011), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n865), .A2(new_n765), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n712), .A2(new_n714), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT62), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n712), .A2(new_n714), .A3(new_n1013), .A4(KEYINPUT62), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1012), .A2(new_n820), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1009), .B1(new_n1019), .B2(new_n427), .ZN(new_n1020));
  OR2_X1    g834(.A1(new_n1020), .A2(KEYINPUT122), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(KEYINPUT122), .ZN(new_n1022));
  NOR3_X1   g836(.A1(new_n844), .A2(new_n674), .A3(new_n737), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n803), .A2(new_n692), .A3(new_n694), .A4(new_n1023), .ZN(new_n1024));
  AND4_X1   g838(.A1(new_n772), .A2(new_n1013), .A3(new_n775), .A4(new_n778), .ZN(new_n1025));
  AND3_X1   g839(.A1(new_n814), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(G953), .B1(new_n1026), .B2(new_n820), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n427), .A2(G900), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1028), .B(KEYINPUT123), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1009), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n1021), .A2(new_n1022), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n427), .B1(G227), .B2(G900), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1031), .B(new_n1032), .ZN(G72));
  NAND4_X1  g847(.A1(new_n1012), .A2(new_n820), .A3(new_n1004), .A4(new_n1018), .ZN(new_n1034));
  XNOR2_X1  g848(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n1035));
  NAND2_X1  g849(.A1(G472), .A2(G902), .ZN(new_n1036));
  XNOR2_X1  g850(.A(new_n1035), .B(new_n1036), .ZN(new_n1037));
  INV_X1    g851(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g853(.A(KEYINPUT125), .B1(new_n1039), .B2(new_n702), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT125), .ZN(new_n1041));
  AOI211_X1 g855(.A(new_n1041), .B(new_n701), .C1(new_n1034), .C2(new_n1038), .ZN(new_n1042));
  OR2_X1    g856(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1026), .A2(new_n820), .A3(new_n1004), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n1044), .A2(KEYINPUT126), .A3(new_n1038), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n700), .A2(new_n341), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g861(.A(KEYINPUT126), .B1(new_n1044), .B2(new_n1038), .ZN(new_n1048));
  OR2_X1    g862(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g863(.A(KEYINPUT127), .ZN(new_n1050));
  NOR3_X1   g864(.A1(new_n702), .A2(new_n1037), .A3(new_n1046), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n964), .B1(new_n923), .B2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g866(.A1(new_n1043), .A2(new_n1049), .A3(new_n1050), .A4(new_n1052), .ZN(new_n1053));
  NOR2_X1   g867(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1054));
  OAI21_X1  g868(.A(new_n1052), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1055));
  OAI21_X1  g869(.A(KEYINPUT127), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n1053), .A2(new_n1056), .ZN(G57));
endmodule


