//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT25), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(G125), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G140), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  OAI211_X1 g009(.A(G146), .B(new_n191), .C1(new_n195), .C2(new_n189), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT73), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G128), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n200), .B(new_n202), .C1(G119), .C2(new_n201), .ZN(new_n203));
  XNOR2_X1  g017(.A(G119), .B(G128), .ZN(new_n204));
  XOR2_X1   g018(.A(KEYINPUT24), .B(G110), .Z(new_n205));
  OAI22_X1  g019(.A1(new_n203), .A2(G110), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G125), .B(G140), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT16), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT73), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G146), .A4(new_n191), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n197), .A2(new_n206), .A3(new_n210), .A4(new_n212), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n203), .A2(G110), .B1(new_n204), .B2(new_n205), .ZN(new_n214));
  INV_X1    g028(.A(new_n196), .ZN(new_n215));
  AOI21_X1  g029(.A(G146), .B1(new_n208), .B2(new_n191), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT22), .B(G137), .ZN(new_n219));
  INV_X1    g033(.A(G953), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(G221), .A3(G234), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n219), .B(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT74), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n218), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n213), .A2(new_n217), .A3(KEYINPUT74), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n222), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n224), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n188), .B1(new_n230), .B2(G902), .ZN(new_n231));
  INV_X1    g045(.A(new_n227), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT74), .B1(new_n213), .B2(new_n217), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n229), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n223), .ZN(new_n235));
  INV_X1    g049(.A(G902), .ZN(new_n236));
  INV_X1    g050(.A(new_n188), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n231), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G217), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(G234), .B2(new_n236), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(G902), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n235), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n211), .A2(G143), .ZN(new_n246));
  INV_X1    g060(.A(G143), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G146), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  OR2_X1    g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n211), .A2(KEYINPUT64), .A3(G143), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n253), .A2(new_n248), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n255), .B1(new_n247), .B2(G146), .ZN(new_n256));
  INV_X1    g070(.A(new_n250), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n254), .A2(KEYINPUT65), .A3(new_n256), .A4(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n256), .A2(new_n253), .A3(new_n248), .A4(new_n257), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT65), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n252), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT11), .ZN(new_n263));
  INV_X1    g077(.A(G134), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(G137), .ZN(new_n265));
  INV_X1    g079(.A(G137), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT11), .A3(G134), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(G137), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n269), .B(G131), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n262), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT1), .B1(new_n247), .B2(G146), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT67), .ZN(new_n273));
  OAI21_X1  g087(.A(G128), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT67), .B1(new_n246), .B2(KEYINPUT1), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n249), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n256), .A2(new_n253), .A3(new_n277), .A4(new_n248), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  OR2_X1    g093(.A1(new_n269), .A2(G131), .ZN(new_n280));
  INV_X1    g094(.A(new_n268), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n264), .A2(G137), .ZN(new_n282));
  OAI21_X1  g096(.A(G131), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n279), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT2), .B(G113), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n199), .A2(G116), .ZN(new_n287));
  INV_X1    g101(.A(G116), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G119), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  OR2_X1    g104(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n286), .A2(new_n290), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n271), .A2(new_n284), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G237), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT69), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT69), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G237), .ZN(new_n299));
  AOI21_X1  g113(.A(G953), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G210), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT27), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT27), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n300), .A2(new_n303), .A3(G210), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT26), .B(G101), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n305), .B1(new_n302), .B2(new_n304), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n295), .A2(KEYINPUT70), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT70), .B1(new_n295), .B2(new_n308), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT68), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n279), .A2(new_n280), .A3(new_n283), .ZN(new_n313));
  INV_X1    g127(.A(G131), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n269), .B(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n252), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n259), .A2(new_n260), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n259), .A2(new_n260), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT66), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n315), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n262), .A2(KEYINPUT66), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n313), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n312), .B1(new_n323), .B2(KEYINPUT30), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n270), .B1(new_n262), .B2(KEYINPUT66), .ZN(new_n325));
  AOI211_X1 g139(.A(new_n320), .B(new_n252), .C1(new_n258), .C2(new_n261), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n284), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT30), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(KEYINPUT68), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n271), .A2(new_n284), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n294), .B1(new_n331), .B2(KEYINPUT30), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n311), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT31), .ZN(new_n334));
  INV_X1    g148(.A(new_n308), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n295), .B(KEYINPUT28), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n327), .A2(new_n293), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n333), .A2(new_n334), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT71), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n327), .A2(KEYINPUT68), .A3(new_n328), .ZN(new_n341));
  AOI21_X1  g155(.A(KEYINPUT68), .B1(new_n327), .B2(new_n328), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n332), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OR2_X1    g157(.A1(new_n309), .A2(new_n310), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n340), .B1(new_n345), .B2(KEYINPUT31), .ZN(new_n346));
  AOI211_X1 g160(.A(KEYINPUT71), .B(new_n334), .C1(new_n343), .C2(new_n344), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n339), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(G472), .A2(G902), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n349), .B(KEYINPUT72), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT32), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OR2_X1    g166(.A1(new_n331), .A2(new_n294), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n336), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n335), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(G902), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n308), .B1(new_n343), .B2(new_n295), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n355), .B1(new_n338), .B2(new_n335), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n348), .A2(new_n352), .B1(G472), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n343), .A2(new_n334), .A3(new_n344), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n338), .A2(new_n335), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT71), .B1(new_n333), .B2(new_n334), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n345), .A2(new_n340), .A3(KEYINPUT31), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n351), .B1(new_n367), .B2(new_n350), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n245), .B1(new_n361), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT9), .B(G234), .ZN(new_n370));
  OAI21_X1  g184(.A(G221), .B1(new_n370), .B2(G902), .ZN(new_n371));
  XNOR2_X1  g185(.A(G110), .B(G140), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(KEYINPUT76), .ZN(new_n373));
  INV_X1    g187(.A(G227), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(G953), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n373), .B(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n377));
  INV_X1    g191(.A(G104), .ZN(new_n378));
  NOR3_X1   g192(.A1(new_n378), .A2(KEYINPUT3), .A3(G107), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  OR2_X1    g194(.A1(KEYINPUT77), .A2(G104), .ZN(new_n381));
  NAND2_X1  g195(.A1(KEYINPUT77), .A2(G104), .ZN(new_n382));
  AOI21_X1  g196(.A(G107), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n380), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n381), .A2(G107), .A3(new_n382), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n377), .B(G101), .C1(new_n385), .C2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G107), .ZN(new_n389));
  AND2_X1   g203(.A1(KEYINPUT77), .A2(G104), .ZN(new_n390));
  NOR2_X1   g204(.A1(KEYINPUT77), .A2(G104), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n379), .B1(new_n392), .B2(KEYINPUT3), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n390), .A2(new_n391), .ZN(new_n394));
  AOI21_X1  g208(.A(G101), .B1(new_n394), .B2(G107), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT4), .ZN(new_n397));
  INV_X1    g211(.A(G101), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n398), .B1(new_n393), .B2(new_n386), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n388), .B(new_n262), .C1(new_n397), .C2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n378), .A2(G107), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n392), .A2(new_n401), .ZN(new_n402));
  AOI22_X1  g216(.A1(new_n393), .A2(new_n395), .B1(new_n402), .B2(G101), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(new_n279), .A3(KEYINPUT10), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT78), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n256), .A2(new_n253), .A3(new_n248), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n272), .A2(G128), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n278), .ZN(new_n409));
  AOI211_X1 g223(.A(new_n405), .B(KEYINPUT10), .C1(new_n403), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n402), .A2(G101), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n396), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT10), .ZN(new_n413));
  AOI21_X1  g227(.A(KEYINPUT78), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n400), .B(new_n404), .C1(new_n410), .C2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n376), .B1(new_n415), .B2(new_n270), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT80), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT80), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n418), .B(new_n376), .C1(new_n415), .C2(new_n270), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT12), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n386), .A2(new_n398), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n411), .B1(new_n385), .B2(new_n421), .ZN(new_n422));
  AND4_X1   g236(.A1(new_n256), .A2(new_n253), .A3(new_n277), .A4(new_n248), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n272), .A2(new_n273), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n246), .A2(KEYINPUT67), .A3(KEYINPUT1), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(G128), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n423), .B1(new_n426), .B2(new_n249), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n428), .A2(KEYINPUT79), .A3(new_n412), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n270), .B1(new_n428), .B2(KEYINPUT79), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n420), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n403), .A2(new_n279), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT79), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n315), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n428), .A2(KEYINPUT79), .A3(new_n412), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(KEYINPUT12), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n431), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n417), .A2(new_n419), .A3(new_n437), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n400), .A2(new_n404), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n439), .B(new_n315), .C1(new_n414), .C2(new_n410), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n415), .A2(new_n270), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n376), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI211_X1 g258(.A(G469), .B(G902), .C1(new_n438), .C2(new_n444), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n429), .A2(new_n430), .A3(new_n420), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT12), .B1(new_n434), .B2(new_n435), .ZN(new_n447));
  OAI22_X1  g261(.A1(new_n446), .A2(new_n447), .B1(new_n415), .B2(new_n270), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n443), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n440), .A2(new_n441), .A3(new_n376), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(G469), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(G469), .A2(G902), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n371), .B1(new_n445), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT87), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n298), .A2(G237), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n296), .A2(KEYINPUT69), .ZN(new_n457));
  OAI211_X1 g271(.A(G214), .B(new_n220), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n247), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n300), .A2(G143), .A3(G214), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n455), .B1(new_n461), .B2(G131), .ZN(new_n462));
  AOI211_X1 g276(.A(KEYINPUT87), .B(new_n314), .C1(new_n459), .C2(new_n460), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT17), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OR3_X1    g278(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT89), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT89), .B1(new_n215), .B2(new_n216), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n458), .A2(new_n247), .ZN(new_n468));
  AOI21_X1  g282(.A(G143), .B1(new_n300), .B2(G214), .ZN(new_n469));
  OAI21_X1  g283(.A(G131), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT87), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n461), .A2(new_n455), .A3(G131), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n459), .A2(new_n314), .A3(new_n460), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT86), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n459), .A2(KEYINPUT86), .A3(new_n460), .A4(new_n314), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n471), .A2(new_n472), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n464), .B(new_n467), .C1(new_n477), .C2(KEYINPUT17), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT85), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT84), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n459), .A2(new_n480), .A3(new_n460), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n480), .B1(new_n459), .B2(new_n460), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(KEYINPUT18), .A2(G131), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n479), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT84), .B1(new_n468), .B2(new_n469), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n459), .A2(new_n480), .A3(new_n460), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT85), .ZN(new_n489));
  INV_X1    g303(.A(new_n461), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n195), .A2(G146), .ZN(new_n491));
  AOI22_X1  g305(.A1(new_n490), .A2(new_n484), .B1(new_n212), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n485), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(G113), .B(G122), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(new_n378), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n478), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n495), .B1(new_n478), .B2(new_n493), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n236), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT90), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g314(.A(KEYINPUT90), .B(new_n236), .C1(new_n496), .C2(new_n497), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(G475), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(G475), .A2(G902), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n197), .A2(new_n210), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n207), .B(KEYINPUT19), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n211), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT88), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT88), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n505), .A2(new_n508), .A3(new_n211), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n504), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n477), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n495), .B1(new_n493), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n503), .B1(new_n496), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT20), .ZN(new_n514));
  INV_X1    g328(.A(new_n495), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n492), .B1(new_n488), .B2(KEYINPUT85), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n483), .A2(new_n479), .A3(new_n484), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n477), .A2(new_n510), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n478), .A2(new_n493), .A3(new_n495), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT20), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n523), .A3(new_n503), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n514), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n247), .A2(G128), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n247), .A2(G128), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT13), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT92), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(new_n528), .B2(new_n526), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n529), .A2(KEYINPUT92), .ZN(new_n532));
  OAI21_X1  g346(.A(G134), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(G122), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT91), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT91), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G122), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n288), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n534), .A2(G116), .ZN(new_n539));
  OR3_X1    g353(.A1(new_n538), .A2(G107), .A3(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(G107), .B1(new_n538), .B2(new_n539), .ZN(new_n541));
  INV_X1    g355(.A(new_n526), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(new_n527), .ZN(new_n543));
  AOI22_X1  g357(.A1(new_n540), .A2(new_n541), .B1(new_n264), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n533), .A2(new_n544), .ZN(new_n545));
  XOR2_X1   g359(.A(new_n539), .B(KEYINPUT14), .Z(new_n546));
  OAI21_X1  g360(.A(G107), .B1(new_n546), .B2(new_n538), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n543), .B(new_n264), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n540), .A3(new_n548), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n370), .A2(new_n240), .A3(G953), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n545), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n545), .B2(new_n549), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n236), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(G478), .ZN(new_n555));
  NOR2_X1   g369(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n555), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  XOR2_X1   g373(.A(new_n554), .B(new_n559), .Z(new_n560));
  NAND3_X1  g374(.A1(new_n502), .A2(new_n525), .A3(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(G210), .B1(G237), .B2(G902), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n388), .B(new_n293), .C1(new_n397), .C2(new_n399), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n290), .A2(KEYINPUT5), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n287), .A2(KEYINPUT5), .ZN(new_n566));
  INV_X1    g380(.A(G113), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n565), .A2(new_n568), .B1(new_n286), .B2(new_n290), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n403), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(G110), .B(G122), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n564), .A2(new_n570), .A3(new_n572), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(KEYINPUT6), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT6), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n571), .A2(new_n577), .A3(new_n573), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n427), .A2(new_n193), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n193), .B2(new_n262), .ZN(new_n580));
  INV_X1    g394(.A(G224), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(G953), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(KEYINPUT81), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n580), .B(new_n583), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n576), .A2(new_n578), .A3(new_n584), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n572), .B(KEYINPUT8), .Z(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n565), .A2(new_n568), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n292), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n422), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n403), .A2(new_n569), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n587), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT82), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT7), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n583), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n580), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n422), .A2(new_n589), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n570), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT82), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n600), .A3(new_n587), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n579), .B(new_n595), .C1(new_n193), .C2(new_n262), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n593), .A2(new_n597), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n575), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n236), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n563), .B1(new_n585), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n576), .A2(new_n578), .A3(new_n584), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n597), .A2(new_n602), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n609), .A2(new_n575), .A3(new_n593), .A4(new_n601), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n607), .A2(new_n610), .A3(new_n236), .A4(new_n562), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n606), .A2(KEYINPUT83), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT83), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n613), .B(new_n563), .C1(new_n585), .C2(new_n605), .ZN(new_n614));
  NAND2_X1  g428(.A1(G234), .A2(G237), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n615), .A2(G952), .A3(new_n220), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT21), .B(G898), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT94), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n615), .A2(G902), .A3(G953), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(G214), .B1(G237), .B2(G902), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n612), .A2(new_n614), .A3(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n454), .A2(new_n561), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n369), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G101), .ZN(G3));
  OAI21_X1  g441(.A(G472), .B1(new_n367), .B2(G902), .ZN(new_n628));
  INV_X1    g442(.A(new_n350), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n348), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n631), .A2(new_n245), .A3(new_n454), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n545), .A2(new_n549), .ZN(new_n634));
  INV_X1    g448(.A(new_n550), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT96), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n551), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n545), .A2(KEYINPUT96), .A3(new_n549), .A4(new_n550), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT97), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n633), .B1(new_n552), .B2(new_n553), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT97), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n636), .A2(new_n638), .A3(new_n643), .A4(new_n639), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n555), .A2(G902), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n641), .A2(new_n642), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n554), .A2(new_n555), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n502), .B2(new_n525), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n606), .A2(KEYINPUT95), .A3(new_n611), .ZN(new_n651));
  INV_X1    g465(.A(new_n620), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT95), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n653), .B(new_n563), .C1(new_n585), .C2(new_n605), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n651), .A2(new_n652), .A3(new_n621), .A4(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n632), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT34), .B(G104), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G6));
  INV_X1    g473(.A(KEYINPUT98), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n523), .B1(new_n522), .B2(new_n503), .ZN(new_n661));
  INV_X1    g475(.A(new_n503), .ZN(new_n662));
  AOI211_X1 g476(.A(KEYINPUT20), .B(new_n662), .C1(new_n520), .C2(new_n521), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n660), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n514), .A2(KEYINPUT98), .A3(new_n524), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n501), .A2(G475), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n560), .B1(new_n667), .B2(new_n500), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n655), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n632), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT35), .B(G107), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  NOR2_X1   g487(.A1(new_n229), .A2(KEYINPUT36), .ZN(new_n674));
  OR2_X1    g488(.A1(new_n228), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n228), .A2(new_n674), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n675), .A2(new_n243), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n239), .B2(new_n241), .ZN(new_n678));
  NOR4_X1   g492(.A1(new_n454), .A2(new_n561), .A3(new_n624), .A4(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n631), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT37), .B(G110), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT99), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n681), .B(new_n683), .ZN(G12));
  INV_X1    g498(.A(new_n371), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n438), .A2(new_n444), .ZN(new_n686));
  INV_X1    g500(.A(G469), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n686), .A2(new_n687), .A3(new_n236), .ZN(new_n688));
  INV_X1    g502(.A(new_n416), .ZN(new_n689));
  AOI22_X1  g503(.A1(new_n689), .A2(new_n441), .B1(new_n448), .B2(new_n443), .ZN(new_n690));
  OAI21_X1  g504(.A(G469), .B1(new_n690), .B2(G902), .ZN(new_n691));
  AOI211_X1 g505(.A(new_n685), .B(new_n678), .C1(new_n688), .C2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(KEYINPUT32), .B1(new_n348), .B2(new_n629), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n360), .A2(G472), .ZN(new_n694));
  INV_X1    g508(.A(new_n352), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n694), .B1(new_n367), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n692), .B1(new_n693), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n611), .A2(KEYINPUT95), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n600), .B1(new_n599), .B2(new_n587), .ZN(new_n699));
  AOI211_X1 g513(.A(KEYINPUT82), .B(new_n586), .C1(new_n598), .C2(new_n570), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n608), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(G902), .B1(new_n701), .B2(new_n575), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n562), .B1(new_n702), .B2(new_n607), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n654), .A2(new_n621), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT100), .B(G900), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n616), .B1(new_n619), .B2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n706), .A2(new_n666), .A3(new_n668), .A4(new_n709), .ZN(new_n710));
  OAI21_X1  g524(.A(KEYINPUT101), .B1(new_n697), .B2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n678), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n371), .B(new_n712), .C1(new_n445), .C2(new_n453), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n713), .B1(new_n361), .B2(new_n368), .ZN(new_n714));
  AND4_X1   g528(.A1(new_n706), .A2(new_n666), .A3(new_n668), .A4(new_n709), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT101), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n711), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G128), .ZN(G30));
  AND2_X1   g533(.A1(new_n353), .A2(new_n295), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n345), .B1(new_n308), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n236), .ZN(new_n722));
  AOI22_X1  g536(.A1(new_n348), .A2(new_n352), .B1(G472), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n368), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(KEYINPUT102), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n560), .B1(new_n502), .B2(new_n525), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n621), .A3(new_n678), .ZN(new_n727));
  XOR2_X1   g541(.A(new_n727), .B(KEYINPUT103), .Z(new_n728));
  AOI21_X1  g542(.A(new_n685), .B1(new_n688), .B2(new_n691), .ZN(new_n729));
  XOR2_X1   g543(.A(new_n708), .B(KEYINPUT39), .Z(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(KEYINPUT40), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n612), .A2(new_n614), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT38), .ZN(new_n734));
  OR4_X1    g548(.A1(new_n725), .A2(new_n728), .A3(new_n732), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G143), .ZN(G45));
  AND3_X1   g550(.A1(new_n649), .A2(new_n706), .A3(new_n709), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n714), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G146), .ZN(G48));
  AOI21_X1  g553(.A(G902), .B1(new_n438), .B2(new_n444), .ZN(new_n740));
  OAI21_X1  g554(.A(KEYINPUT104), .B1(new_n740), .B2(new_n687), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT104), .ZN(new_n742));
  AOI22_X1  g556(.A1(new_n416), .A2(KEYINPUT80), .B1(new_n436), .B2(new_n431), .ZN(new_n743));
  AOI22_X1  g557(.A1(new_n743), .A2(new_n419), .B1(new_n442), .B2(new_n443), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n742), .B(G469), .C1(new_n744), .C2(G902), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n445), .A2(new_n685), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n369), .A2(new_n656), .A3(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(KEYINPUT41), .B(G113), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G15));
  NAND3_X1  g565(.A1(new_n369), .A2(new_n670), .A3(new_n748), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G116), .ZN(G18));
  INV_X1    g567(.A(KEYINPUT105), .ZN(new_n754));
  INV_X1    g568(.A(new_n561), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n678), .A2(new_n620), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n755), .B(new_n756), .C1(new_n693), .C2(new_n696), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n746), .A2(new_n747), .A3(new_n706), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n754), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n758), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n361), .A2(new_n368), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n561), .A2(new_n620), .A3(new_n678), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n760), .A2(KEYINPUT105), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G119), .ZN(G21));
  NAND2_X1  g579(.A1(new_n331), .A2(KEYINPUT30), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n293), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n767), .B1(new_n324), .B2(new_n329), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT31), .B1(new_n768), .B2(new_n311), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n336), .A2(new_n353), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n335), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n769), .A2(new_n362), .A3(new_n771), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n772), .A2(KEYINPUT106), .A3(new_n629), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT106), .B1(new_n772), .B2(new_n629), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n245), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n776), .A3(new_n628), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n704), .A2(new_n705), .A3(new_n620), .ZN(new_n779));
  AND4_X1   g593(.A1(new_n779), .A2(new_n746), .A3(new_n726), .A4(new_n747), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G122), .ZN(G24));
  NAND2_X1  g596(.A1(new_n501), .A2(G475), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n478), .A2(new_n493), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n515), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n521), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT90), .B1(new_n786), .B2(new_n236), .ZN(new_n787));
  OAI22_X1  g601(.A1(new_n783), .A2(new_n787), .B1(new_n661), .B2(new_n663), .ZN(new_n788));
  INV_X1    g602(.A(new_n648), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n789), .A3(new_n709), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n758), .A2(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n775), .A2(new_n628), .A3(new_n712), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G125), .ZN(G27));
  INV_X1    g608(.A(KEYINPUT42), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n776), .B1(new_n693), .B2(new_n696), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n622), .B1(new_n612), .B2(new_n614), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n649), .A2(new_n729), .A3(new_n797), .A4(new_n709), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n795), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n729), .A2(new_n649), .A3(new_n709), .A4(new_n797), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n369), .A3(KEYINPUT42), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G131), .ZN(G33));
  NOR3_X1   g617(.A1(new_n669), .A2(new_n454), .A3(new_n708), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n369), .A3(new_n797), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G134), .ZN(G36));
  INV_X1    g620(.A(new_n788), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n789), .ZN(new_n808));
  XOR2_X1   g622(.A(new_n808), .B(KEYINPUT43), .Z(new_n809));
  AND3_X1   g623(.A1(new_n809), .A2(new_n631), .A3(new_n712), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n810), .A2(KEYINPUT44), .ZN(new_n811));
  OAI21_X1  g625(.A(G469), .B1(new_n690), .B2(KEYINPUT45), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n812), .A2(KEYINPUT107), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n690), .A2(KEYINPUT45), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n812), .A2(KEYINPUT107), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT46), .B1(new_n816), .B2(new_n452), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n817), .B1(new_n687), .B2(new_n740), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(KEYINPUT46), .A3(new_n452), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n685), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n820), .A2(new_n730), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n810), .A2(KEYINPUT44), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n811), .A2(new_n821), .A3(new_n797), .A4(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G137), .ZN(G39));
  NAND2_X1  g638(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n820), .A2(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n788), .A2(new_n789), .A3(new_n709), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n245), .A3(new_n797), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n761), .ZN(new_n829));
  XOR2_X1   g643(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n830));
  OAI211_X1 g644(.A(new_n826), .B(new_n829), .C1(new_n820), .C2(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G140), .ZN(G42));
  INV_X1    g646(.A(G952), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n220), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT117), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n734), .A2(new_n748), .A3(new_n622), .ZN(new_n837));
  AND4_X1   g651(.A1(new_n616), .A2(new_n809), .A3(new_n778), .A4(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT50), .ZN(new_n840));
  OR3_X1    g654(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n840), .B1(new_n838), .B2(new_n839), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n809), .A2(new_n616), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n748), .A2(new_n797), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n616), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n844), .A2(new_n245), .A3(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n847), .A2(new_n725), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n788), .A2(new_n789), .ZN(new_n849));
  AOI22_X1  g663(.A1(new_n845), .A2(new_n792), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n841), .A2(new_n842), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n843), .A2(new_n777), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n797), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n826), .B1(new_n820), .B2(new_n830), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n746), .A2(new_n688), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n371), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n858), .B1(new_n857), .B2(new_n856), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n853), .B1(new_n854), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n836), .B1(new_n851), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n848), .A2(new_n649), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n845), .A2(new_n369), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT48), .ZN(new_n864));
  AOI211_X1 g678(.A(new_n833), .B(G953), .C1(new_n852), .C2(new_n760), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n861), .A2(new_n862), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  OR3_X1    g680(.A1(new_n851), .A2(new_n860), .A3(new_n836), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n867), .A2(KEYINPUT116), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(KEYINPUT116), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT113), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n726), .A2(new_n706), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n678), .A2(new_n709), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n454), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n724), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n775), .A2(new_n628), .A3(new_n712), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n827), .A2(new_n706), .A3(new_n746), .A4(new_n747), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n738), .B(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT52), .B1(new_n879), .B2(new_n718), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n697), .A2(KEYINPUT101), .A3(new_n710), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n716), .B1(new_n714), .B2(new_n715), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT52), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n883), .A2(new_n878), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n871), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n884), .B1(new_n883), .B2(new_n878), .ZN(new_n887));
  AOI22_X1  g701(.A1(new_n791), .A2(new_n792), .B1(new_n714), .B2(new_n737), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n718), .A2(KEYINPUT52), .A3(new_n888), .A4(new_n875), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n887), .A2(KEYINPUT113), .A3(new_n889), .ZN(new_n890));
  AOI22_X1  g704(.A1(new_n679), .A2(new_n680), .B1(new_n369), .B2(new_n625), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n369), .B(new_n748), .C1(new_n656), .C2(new_n670), .ZN(new_n892));
  INV_X1    g706(.A(new_n560), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n502), .A2(new_n525), .A3(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT109), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n502), .A2(new_n525), .A3(KEYINPUT109), .A4(new_n893), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n896), .A2(new_n650), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n624), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n454), .A2(new_n245), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n898), .A2(new_n680), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n891), .A2(new_n892), .A3(new_n901), .A4(new_n781), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n759), .A2(new_n763), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n792), .A2(new_n800), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n502), .A2(new_n560), .A3(new_n709), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n666), .A3(new_n797), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT110), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n906), .A2(KEYINPUT110), .A3(new_n797), .A4(new_n666), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n909), .A2(new_n714), .A3(new_n910), .ZN(new_n911));
  AND4_X1   g725(.A1(new_n802), .A2(new_n805), .A3(new_n905), .A4(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT111), .B1(new_n904), .B2(new_n912), .ZN(new_n913));
  AOI22_X1  g727(.A1(new_n894), .A2(new_n895), .B1(new_n788), .B2(new_n789), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n624), .B1(new_n914), .B2(new_n897), .ZN(new_n915));
  AOI22_X1  g729(.A1(new_n632), .A2(new_n915), .B1(new_n778), .B2(new_n780), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n764), .A2(new_n916), .A3(new_n891), .A4(new_n892), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n802), .A2(new_n805), .A3(new_n905), .A4(new_n911), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT111), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n886), .B(new_n890), .C1(new_n913), .C2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(KEYINPUT53), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n904), .A2(new_n912), .A3(KEYINPUT111), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n919), .B1(new_n917), .B2(new_n918), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT53), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT112), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n880), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n887), .A2(KEYINPUT112), .A3(new_n889), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n925), .A2(new_n926), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n922), .A2(KEYINPUT54), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n921), .A2(new_n926), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT54), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n917), .A2(new_n918), .A3(new_n926), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n934), .A2(new_n928), .A3(new_n929), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n932), .A2(new_n933), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n931), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n835), .B1(new_n870), .B2(new_n938), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n245), .A2(new_n622), .A3(new_n685), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n734), .A2(new_n807), .A3(new_n789), .A4(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(KEYINPUT49), .B2(new_n855), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n942), .B(new_n725), .C1(KEYINPUT49), .C2(new_n855), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n939), .A2(new_n943), .ZN(G75));
  NOR2_X1   g758(.A1(new_n220), .A2(G952), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n935), .B1(new_n921), .B2(new_n926), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n947), .A2(new_n236), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT56), .B1(new_n948), .B2(G210), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n576), .A2(new_n578), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(new_n584), .Z(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT55), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n946), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(new_n949), .B2(new_n953), .ZN(G51));
  XOR2_X1   g769(.A(new_n452), .B(KEYINPUT57), .Z(new_n956));
  AND3_X1   g770(.A1(new_n887), .A2(KEYINPUT113), .A3(new_n889), .ZN(new_n957));
  AOI21_X1  g771(.A(KEYINPUT113), .B1(new_n887), .B2(new_n889), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(KEYINPUT53), .B1(new_n959), .B2(new_n925), .ZN(new_n960));
  OAI21_X1  g774(.A(KEYINPUT54), .B1(new_n960), .B2(new_n935), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n937), .B2(KEYINPUT118), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT118), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(new_n947), .B2(new_n933), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n956), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n744), .B(KEYINPUT119), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(G902), .B1(new_n960), .B2(new_n935), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n968), .A2(new_n816), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n945), .B1(new_n967), .B2(new_n969), .ZN(G54));
  NAND4_X1  g784(.A1(new_n948), .A2(KEYINPUT58), .A3(G475), .A4(new_n522), .ZN(new_n971));
  NAND2_X1  g785(.A1(KEYINPUT58), .A2(G475), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n521), .B(new_n520), .C1(new_n968), .C2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n971), .A2(new_n973), .A3(new_n946), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT120), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n971), .A2(new_n973), .A3(KEYINPUT120), .A4(new_n946), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(G60));
  NAND2_X1  g792(.A1(G478), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT59), .Z(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n922), .A2(KEYINPUT54), .A3(new_n930), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n960), .A2(KEYINPUT54), .A3(new_n935), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT121), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n980), .B1(new_n931), .B2(new_n937), .ZN(new_n988));
  INV_X1    g802(.A(new_n986), .ZN(new_n989));
  OAI21_X1  g803(.A(KEYINPUT121), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n986), .A2(new_n980), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n991), .B1(new_n962), .B2(new_n964), .ZN(new_n992));
  AND4_X1   g806(.A1(new_n946), .A2(new_n987), .A3(new_n990), .A4(new_n992), .ZN(G63));
  INV_X1    g807(.A(KEYINPUT61), .ZN(new_n994));
  NAND2_X1  g808(.A1(G217), .A2(G902), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT60), .ZN(new_n996));
  OAI21_X1  g810(.A(KEYINPUT122), .B1(new_n947), .B2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT122), .ZN(new_n998));
  INV_X1    g812(.A(new_n996), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n998), .B(new_n999), .C1(new_n960), .C2(new_n935), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n997), .A2(new_n230), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n946), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n675), .A2(new_n676), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1004), .B1(new_n997), .B2(new_n1000), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n994), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n997), .A2(new_n1000), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n1003), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1008), .A2(KEYINPUT61), .A3(new_n946), .A4(new_n1001), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1006), .A2(new_n1009), .ZN(G66));
  OAI21_X1  g824(.A(G953), .B1(new_n618), .B2(new_n581), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1011), .B1(new_n904), .B2(G953), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT123), .Z(new_n1013));
  OAI21_X1  g827(.A(new_n950), .B1(G898), .B2(new_n220), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1013), .B(new_n1014), .ZN(G69));
  NAND3_X1  g829(.A1(new_n821), .A2(new_n369), .A3(new_n872), .ZN(new_n1016));
  AND2_X1   g830(.A1(new_n823), .A2(new_n1016), .ZN(new_n1017));
  AND3_X1   g831(.A1(new_n831), .A2(new_n802), .A3(new_n805), .ZN(new_n1018));
  AND2_X1   g832(.A1(new_n718), .A2(new_n888), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1017), .A2(new_n1018), .A3(new_n220), .A4(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n330), .A2(new_n766), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1021), .B(new_n505), .Z(new_n1022));
  INV_X1    g836(.A(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1023), .B1(G900), .B2(G953), .ZN(new_n1024));
  AND3_X1   g838(.A1(new_n1020), .A2(KEYINPUT125), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n731), .ZN(new_n1026));
  NAND4_X1  g840(.A1(new_n898), .A2(new_n369), .A3(new_n1026), .A4(new_n797), .ZN(new_n1027));
  AND3_X1   g841(.A1(new_n823), .A2(new_n831), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n735), .A2(new_n1019), .ZN(new_n1029));
  OR2_X1    g843(.A1(new_n1029), .A2(KEYINPUT62), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1029), .A2(KEYINPUT62), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1028), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1022), .B1(new_n1032), .B2(new_n220), .ZN(new_n1033));
  AOI21_X1  g847(.A(KEYINPUT125), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1034));
  NOR3_X1   g848(.A1(new_n1025), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g849(.A(G900), .ZN(new_n1036));
  OAI21_X1  g850(.A(G953), .B1(new_n374), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1038));
  XOR2_X1   g852(.A(new_n1037), .B(KEYINPUT124), .Z(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI22_X1  g854(.A1(new_n1035), .A2(new_n1037), .B1(new_n1033), .B2(new_n1040), .ZN(G72));
  AND2_X1   g855(.A1(new_n343), .A2(new_n295), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n1042), .A2(new_n335), .ZN(new_n1043));
  NAND4_X1  g857(.A1(new_n1028), .A2(new_n904), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1044));
  INV_X1    g858(.A(KEYINPUT126), .ZN(new_n1045));
  NAND2_X1  g859(.A1(G472), .A2(G902), .ZN(new_n1046));
  XOR2_X1   g860(.A(new_n1046), .B(KEYINPUT63), .Z(new_n1047));
  AND3_X1   g861(.A1(new_n1044), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1045), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1043), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n345), .B1(new_n1042), .B2(new_n308), .ZN(new_n1051));
  NAND4_X1  g865(.A1(new_n922), .A2(new_n930), .A3(new_n1047), .A4(new_n1051), .ZN(new_n1052));
  NAND3_X1  g866(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n1047), .B1(new_n1053), .B2(new_n917), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1042), .A2(new_n335), .ZN(new_n1055));
  XOR2_X1   g869(.A(new_n1055), .B(KEYINPUT127), .Z(new_n1056));
  AOI21_X1  g870(.A(new_n945), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  AND3_X1   g871(.A1(new_n1050), .A2(new_n1052), .A3(new_n1057), .ZN(G57));
endmodule


