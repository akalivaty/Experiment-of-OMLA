

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582;

  NOR2_X1 U321 ( .A1(n525), .A2(n453), .ZN(n467) );
  XOR2_X1 U322 ( .A(G211GAT), .B(KEYINPUT21), .Z(n289) );
  XOR2_X1 U323 ( .A(n397), .B(n358), .Z(n290) );
  XOR2_X1 U324 ( .A(G218GAT), .B(G106GAT), .Z(n291) );
  XOR2_X1 U325 ( .A(KEYINPUT40), .B(n493), .Z(n292) );
  XNOR2_X1 U326 ( .A(n382), .B(KEYINPUT48), .ZN(n383) );
  XNOR2_X1 U327 ( .A(n314), .B(n291), .ZN(n315) );
  INV_X1 U328 ( .A(KEYINPUT120), .ZN(n427) );
  XNOR2_X1 U329 ( .A(n384), .B(n383), .ZN(n522) );
  XNOR2_X1 U330 ( .A(n316), .B(n315), .ZN(n321) );
  XNOR2_X1 U331 ( .A(n427), .B(KEYINPUT55), .ZN(n428) );
  XNOR2_X1 U332 ( .A(n335), .B(n334), .ZN(n377) );
  XNOR2_X1 U333 ( .A(n429), .B(n428), .ZN(n443) );
  NOR2_X1 U334 ( .A1(n508), .A2(n484), .ZN(n485) );
  XOR2_X1 U335 ( .A(n452), .B(KEYINPUT28), .Z(n517) );
  XNOR2_X1 U336 ( .A(n444), .B(KEYINPUT122), .ZN(n445) );
  XNOR2_X1 U337 ( .A(n446), .B(n445), .ZN(G1350GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT77), .B(G211GAT), .Z(n294) );
  XNOR2_X1 U339 ( .A(G127GAT), .B(G78GAT), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U341 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n296) );
  XNOR2_X1 U342 ( .A(KEYINPUT78), .B(KEYINPUT12), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n298), .B(n297), .ZN(n307) );
  XNOR2_X1 U345 ( .A(G8GAT), .B(G183GAT), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n299), .B(KEYINPUT76), .ZN(n389) );
  XNOR2_X1 U347 ( .A(G71GAT), .B(G57GAT), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n300), .B(KEYINPUT13), .ZN(n333) );
  XOR2_X1 U349 ( .A(G64GAT), .B(n333), .Z(n302) );
  NAND2_X1 U350 ( .A1(G231GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U351 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U352 ( .A(n389), .B(n303), .Z(n305) );
  XOR2_X1 U353 ( .A(G15GAT), .B(G1GAT), .Z(n338) );
  XOR2_X1 U354 ( .A(G22GAT), .B(G155GAT), .Z(n310) );
  XNOR2_X1 U355 ( .A(n338), .B(n310), .ZN(n304) );
  XNOR2_X1 U356 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U357 ( .A(n307), .B(n306), .Z(n448) );
  XOR2_X1 U358 ( .A(n448), .B(KEYINPUT111), .Z(n531) );
  XNOR2_X1 U359 ( .A(G197GAT), .B(KEYINPUT82), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n289), .B(n308), .ZN(n397) );
  XOR2_X1 U361 ( .A(G50GAT), .B(G162GAT), .Z(n358) );
  NAND2_X1 U362 ( .A1(G228GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n290), .B(n309), .ZN(n311) );
  XOR2_X1 U364 ( .A(n311), .B(n310), .Z(n316) );
  XOR2_X1 U365 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n313) );
  XNOR2_X1 U366 ( .A(KEYINPUT24), .B(KEYINPUT81), .ZN(n312) );
  XNOR2_X1 U367 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U368 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n317), .B(KEYINPUT2), .ZN(n408) );
  XOR2_X1 U370 ( .A(G78GAT), .B(G148GAT), .Z(n319) );
  XNOR2_X1 U371 ( .A(KEYINPUT69), .B(G204GAT), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n328) );
  XNOR2_X1 U373 ( .A(n408), .B(n328), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n459) );
  XOR2_X1 U375 ( .A(KEYINPUT70), .B(KEYINPUT32), .Z(n323) );
  NAND2_X1 U376 ( .A1(G230GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U377 ( .A(n323), .B(n322), .ZN(n325) );
  INV_X1 U378 ( .A(KEYINPUT31), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n325), .B(n324), .ZN(n330) );
  XNOR2_X1 U380 ( .A(G99GAT), .B(G106GAT), .ZN(n327) );
  XOR2_X1 U381 ( .A(G92GAT), .B(G85GAT), .Z(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n367) );
  XNOR2_X1 U383 ( .A(n328), .B(n367), .ZN(n329) );
  XOR2_X1 U384 ( .A(n330), .B(n329), .Z(n331) );
  XOR2_X1 U385 ( .A(G176GAT), .B(G64GAT), .Z(n388) );
  XNOR2_X1 U386 ( .A(n331), .B(n388), .ZN(n335) );
  XNOR2_X1 U387 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U389 ( .A(KEYINPUT41), .B(n377), .ZN(n541) );
  XOR2_X1 U390 ( .A(G22GAT), .B(G141GAT), .Z(n337) );
  XNOR2_X1 U391 ( .A(G169GAT), .B(G113GAT), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n337), .B(n336), .ZN(n353) );
  XOR2_X1 U393 ( .A(n338), .B(G50GAT), .Z(n342) );
  XOR2_X1 U394 ( .A(G29GAT), .B(G43GAT), .Z(n340) );
  XNOR2_X1 U395 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n339) );
  XNOR2_X1 U396 ( .A(n340), .B(n339), .ZN(n368) );
  XNOR2_X1 U397 ( .A(G36GAT), .B(n368), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U399 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n344) );
  NAND2_X1 U400 ( .A1(G229GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U401 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U402 ( .A(n346), .B(n345), .Z(n351) );
  XOR2_X1 U403 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n348) );
  XNOR2_X1 U404 ( .A(G197GAT), .B(G8GAT), .ZN(n347) );
  XNOR2_X1 U405 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n349), .B(KEYINPUT29), .ZN(n350) );
  XNOR2_X1 U407 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U408 ( .A(n353), .B(n352), .Z(n567) );
  NAND2_X1 U409 ( .A1(n541), .A2(n567), .ZN(n355) );
  XNOR2_X1 U410 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n354) );
  XNOR2_X1 U411 ( .A(n355), .B(n354), .ZN(n356) );
  NAND2_X1 U412 ( .A1(n356), .A2(n531), .ZN(n357) );
  XNOR2_X1 U413 ( .A(n357), .B(KEYINPUT113), .ZN(n373) );
  XNOR2_X1 U414 ( .A(n358), .B(KEYINPUT11), .ZN(n359) );
  XNOR2_X1 U415 ( .A(n359), .B(KEYINPUT9), .ZN(n372) );
  XNOR2_X1 U416 ( .A(G36GAT), .B(G190GAT), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n360), .B(G218GAT), .ZN(n396) );
  XOR2_X1 U418 ( .A(n396), .B(KEYINPUT74), .Z(n362) );
  NAND2_X1 U419 ( .A1(G232GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U421 ( .A(KEYINPUT10), .B(KEYINPUT72), .Z(n364) );
  XNOR2_X1 U422 ( .A(G134GAT), .B(KEYINPUT73), .ZN(n363) );
  XNOR2_X1 U423 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U425 ( .A(n368), .B(n367), .Z(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n372), .B(n371), .ZN(n550) );
  NAND2_X1 U428 ( .A1(n373), .A2(n550), .ZN(n374) );
  XNOR2_X1 U429 ( .A(n374), .B(KEYINPUT47), .ZN(n381) );
  XOR2_X1 U430 ( .A(KEYINPUT45), .B(KEYINPUT114), .Z(n376) );
  INV_X1 U431 ( .A(n448), .ZN(n575) );
  XNOR2_X1 U432 ( .A(KEYINPUT75), .B(n550), .ZN(n560) );
  XNOR2_X1 U433 ( .A(KEYINPUT36), .B(n560), .ZN(n578) );
  NAND2_X1 U434 ( .A1(n575), .A2(n578), .ZN(n375) );
  XNOR2_X1 U435 ( .A(n376), .B(n375), .ZN(n378) );
  NAND2_X1 U436 ( .A1(n378), .A2(n377), .ZN(n379) );
  NOR2_X1 U437 ( .A1(n379), .A2(n567), .ZN(n380) );
  NOR2_X1 U438 ( .A1(n381), .A2(n380), .ZN(n384) );
  XOR2_X1 U439 ( .A(KEYINPUT115), .B(KEYINPUT64), .Z(n382) );
  XOR2_X1 U440 ( .A(KEYINPUT79), .B(KEYINPUT17), .Z(n386) );
  XNOR2_X1 U441 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U443 ( .A(G169GAT), .B(n387), .Z(n440) );
  XOR2_X1 U444 ( .A(n389), .B(n388), .Z(n391) );
  NAND2_X1 U445 ( .A1(G226GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U446 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U447 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n393) );
  XNOR2_X1 U448 ( .A(G204GAT), .B(G92GAT), .ZN(n392) );
  XNOR2_X1 U449 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U450 ( .A(n395), .B(n394), .Z(n399) );
  XNOR2_X1 U451 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U452 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U453 ( .A(n440), .B(n400), .Z(n514) );
  INV_X1 U454 ( .A(n514), .ZN(n490) );
  NOR2_X1 U455 ( .A1(n522), .A2(n490), .ZN(n401) );
  XNOR2_X1 U456 ( .A(n401), .B(KEYINPUT54), .ZN(n426) );
  XOR2_X1 U457 ( .A(KEYINPUT89), .B(KEYINPUT5), .Z(n403) );
  XNOR2_X1 U458 ( .A(KEYINPUT86), .B(KEYINPUT85), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U460 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n405) );
  XNOR2_X1 U461 ( .A(KEYINPUT4), .B(KEYINPUT83), .ZN(n404) );
  XNOR2_X1 U462 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U463 ( .A(n407), .B(n406), .Z(n413) );
  XOR2_X1 U464 ( .A(G85GAT), .B(n408), .Z(n410) );
  NAND2_X1 U465 ( .A1(G225GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U467 ( .A(G29GAT), .B(n411), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U469 ( .A(G57GAT), .B(G162GAT), .Z(n415) );
  XNOR2_X1 U470 ( .A(G148GAT), .B(G155GAT), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U472 ( .A(n417), .B(n416), .Z(n425) );
  XOR2_X1 U473 ( .A(G127GAT), .B(G134GAT), .Z(n419) );
  XNOR2_X1 U474 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U476 ( .A(G113GAT), .B(n420), .Z(n439) );
  XOR2_X1 U477 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n422) );
  XNOR2_X1 U478 ( .A(G1GAT), .B(KEYINPUT84), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n439), .B(n423), .ZN(n424) );
  XOR2_X1 U481 ( .A(n425), .B(n424), .Z(n511) );
  INV_X1 U482 ( .A(n511), .ZN(n486) );
  NAND2_X1 U483 ( .A1(n426), .A2(n486), .ZN(n565) );
  NOR2_X1 U484 ( .A1(n459), .A2(n565), .ZN(n429) );
  XOR2_X1 U485 ( .A(G71GAT), .B(G99GAT), .Z(n431) );
  XNOR2_X1 U486 ( .A(G43GAT), .B(G190GAT), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U488 ( .A(G183GAT), .B(n432), .Z(n434) );
  NAND2_X1 U489 ( .A1(G227GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U490 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U491 ( .A(KEYINPUT80), .B(G176GAT), .Z(n436) );
  XNOR2_X1 U492 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n435) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U494 ( .A(n438), .B(n437), .Z(n442) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U496 ( .A(n442), .B(n441), .Z(n492) );
  INV_X1 U497 ( .A(n492), .ZN(n525) );
  NAND2_X1 U498 ( .A1(n443), .A2(n525), .ZN(n559) );
  NOR2_X1 U499 ( .A1(n531), .A2(n559), .ZN(n446) );
  INV_X1 U500 ( .A(G183GAT), .ZN(n444) );
  INV_X1 U501 ( .A(n567), .ZN(n552) );
  INV_X1 U502 ( .A(n377), .ZN(n572) );
  NOR2_X1 U503 ( .A1(n552), .A2(n572), .ZN(n447) );
  XNOR2_X1 U504 ( .A(n447), .B(KEYINPUT71), .ZN(n484) );
  NOR2_X1 U505 ( .A1(n560), .A2(n448), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n449), .B(KEYINPUT16), .ZN(n469) );
  XNOR2_X1 U507 ( .A(KEYINPUT27), .B(KEYINPUT92), .ZN(n450) );
  XOR2_X1 U508 ( .A(n450), .B(n514), .Z(n462) );
  NOR2_X1 U509 ( .A1(n486), .A2(n462), .ZN(n451) );
  XOR2_X1 U510 ( .A(KEYINPUT93), .B(n451), .Z(n539) );
  XNOR2_X1 U511 ( .A(n459), .B(KEYINPUT65), .ZN(n452) );
  INV_X1 U512 ( .A(n517), .ZN(n495) );
  NAND2_X1 U513 ( .A1(n539), .A2(n495), .ZN(n523) );
  XNOR2_X1 U514 ( .A(KEYINPUT94), .B(n523), .ZN(n453) );
  XNOR2_X1 U515 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n454) );
  XNOR2_X1 U516 ( .A(n454), .B(KEYINPUT25), .ZN(n458) );
  NOR2_X1 U517 ( .A1(n492), .A2(n490), .ZN(n455) );
  XNOR2_X1 U518 ( .A(n455), .B(KEYINPUT96), .ZN(n456) );
  NOR2_X1 U519 ( .A1(n459), .A2(n456), .ZN(n457) );
  XNOR2_X1 U520 ( .A(n458), .B(n457), .ZN(n464) );
  XOR2_X1 U521 ( .A(KEYINPUT26), .B(KEYINPUT95), .Z(n461) );
  NAND2_X1 U522 ( .A1(n459), .A2(n492), .ZN(n460) );
  XNOR2_X1 U523 ( .A(n461), .B(n460), .ZN(n566) );
  NOR2_X1 U524 ( .A1(n462), .A2(n566), .ZN(n463) );
  NOR2_X1 U525 ( .A1(n464), .A2(n463), .ZN(n465) );
  NOR2_X1 U526 ( .A1(n465), .A2(n511), .ZN(n466) );
  NOR2_X1 U527 ( .A1(n467), .A2(n466), .ZN(n480) );
  INV_X1 U528 ( .A(n480), .ZN(n468) );
  NAND2_X1 U529 ( .A1(n469), .A2(n468), .ZN(n497) );
  NOR2_X1 U530 ( .A1(n484), .A2(n497), .ZN(n477) );
  NAND2_X1 U531 ( .A1(n511), .A2(n477), .ZN(n470) );
  XNOR2_X1 U532 ( .A(n470), .B(KEYINPUT34), .ZN(n471) );
  XNOR2_X1 U533 ( .A(G1GAT), .B(n471), .ZN(G1324GAT) );
  XOR2_X1 U534 ( .A(G8GAT), .B(KEYINPUT99), .Z(n473) );
  NAND2_X1 U535 ( .A1(n477), .A2(n514), .ZN(n472) );
  XNOR2_X1 U536 ( .A(n473), .B(n472), .ZN(G1325GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT35), .B(KEYINPUT100), .Z(n475) );
  NAND2_X1 U538 ( .A1(n477), .A2(n525), .ZN(n474) );
  XNOR2_X1 U539 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U540 ( .A(G15GAT), .B(n476), .ZN(G1326GAT) );
  XOR2_X1 U541 ( .A(G22GAT), .B(KEYINPUT101), .Z(n479) );
  NAND2_X1 U542 ( .A1(n477), .A2(n517), .ZN(n478) );
  XNOR2_X1 U543 ( .A(n479), .B(n478), .ZN(G1327GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT37), .B(KEYINPUT102), .Z(n483) );
  NOR2_X1 U545 ( .A1(n575), .A2(n480), .ZN(n481) );
  NAND2_X1 U546 ( .A1(n481), .A2(n578), .ZN(n482) );
  XNOR2_X1 U547 ( .A(n483), .B(n482), .ZN(n508) );
  XOR2_X1 U548 ( .A(KEYINPUT38), .B(n485), .Z(n494) );
  NOR2_X1 U549 ( .A1(n494), .A2(n486), .ZN(n489) );
  XOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT39), .Z(n487) );
  XNOR2_X1 U551 ( .A(KEYINPUT103), .B(n487), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n489), .B(n488), .ZN(G1328GAT) );
  NOR2_X1 U553 ( .A1(n494), .A2(n490), .ZN(n491) );
  XOR2_X1 U554 ( .A(G36GAT), .B(n491), .Z(G1329GAT) );
  NOR2_X1 U555 ( .A1(n494), .A2(n492), .ZN(n493) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n292), .ZN(G1330GAT) );
  NOR2_X1 U557 ( .A1(n495), .A2(n494), .ZN(n496) );
  XOR2_X1 U558 ( .A(G50GAT), .B(n496), .Z(G1331GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT107), .B(KEYINPUT106), .Z(n499) );
  XNOR2_X1 U560 ( .A(n541), .B(KEYINPUT105), .ZN(n555) );
  OR2_X1 U561 ( .A1(n555), .A2(n567), .ZN(n509) );
  NOR2_X1 U562 ( .A1(n509), .A2(n497), .ZN(n505) );
  NAND2_X1 U563 ( .A1(n505), .A2(n511), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n499), .B(n498), .ZN(n501) );
  XOR2_X1 U565 ( .A(G57GAT), .B(KEYINPUT42), .Z(n500) );
  XNOR2_X1 U566 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U567 ( .A(KEYINPUT104), .B(n502), .Z(G1332GAT) );
  NAND2_X1 U568 ( .A1(n505), .A2(n514), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n503), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U570 ( .A1(n505), .A2(n525), .ZN(n504) );
  XNOR2_X1 U571 ( .A(n504), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U572 ( .A(G78GAT), .B(KEYINPUT43), .Z(n507) );
  NAND2_X1 U573 ( .A1(n505), .A2(n517), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n507), .B(n506), .ZN(G1335GAT) );
  XOR2_X1 U575 ( .A(G85GAT), .B(KEYINPUT109), .Z(n513) );
  NOR2_X1 U576 ( .A1(n509), .A2(n508), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n510), .B(KEYINPUT108), .ZN(n518) );
  NAND2_X1 U578 ( .A1(n518), .A2(n511), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(G1336GAT) );
  NAND2_X1 U580 ( .A1(n514), .A2(n518), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G92GAT), .B(n515), .ZN(G1337GAT) );
  NAND2_X1 U582 ( .A1(n518), .A2(n525), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n516), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT110), .B(KEYINPUT44), .Z(n520) );
  NAND2_X1 U585 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U587 ( .A(G106GAT), .B(n521), .Z(G1339GAT) );
  NOR2_X1 U588 ( .A1(n522), .A2(n523), .ZN(n524) );
  NAND2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n534) );
  NOR2_X1 U590 ( .A1(n552), .A2(n534), .ZN(n527) );
  XNOR2_X1 U591 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G113GAT), .B(n528), .ZN(G1340GAT) );
  NOR2_X1 U594 ( .A1(n555), .A2(n534), .ZN(n530) );
  XNOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n530), .B(n529), .ZN(G1341GAT) );
  NOR2_X1 U597 ( .A1(n531), .A2(n534), .ZN(n532) );
  XOR2_X1 U598 ( .A(KEYINPUT50), .B(n532), .Z(n533) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(n533), .ZN(G1342GAT) );
  XOR2_X1 U600 ( .A(G134GAT), .B(KEYINPUT51), .Z(n537) );
  INV_X1 U601 ( .A(n534), .ZN(n535) );
  NAND2_X1 U602 ( .A1(n535), .A2(n560), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(G1343GAT) );
  NOR2_X1 U604 ( .A1(n522), .A2(n566), .ZN(n538) );
  NAND2_X1 U605 ( .A1(n539), .A2(n538), .ZN(n549) );
  NOR2_X1 U606 ( .A1(n552), .A2(n549), .ZN(n540) );
  XOR2_X1 U607 ( .A(G141GAT), .B(n540), .Z(G1344GAT) );
  INV_X1 U608 ( .A(n549), .ZN(n546) );
  NAND2_X1 U609 ( .A1(n546), .A2(n541), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n542), .B(KEYINPUT118), .ZN(n543) );
  XOR2_X1 U611 ( .A(n543), .B(KEYINPUT53), .Z(n545) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(G1345GAT) );
  XOR2_X1 U614 ( .A(G155GAT), .B(KEYINPUT119), .Z(n548) );
  NAND2_X1 U615 ( .A1(n546), .A2(n575), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(G1346GAT) );
  NOR2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U618 ( .A(G162GAT), .B(n551), .Z(G1347GAT) );
  NOR2_X1 U619 ( .A1(n552), .A2(n559), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(G169GAT), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(KEYINPUT121), .ZN(G1348GAT) );
  NOR2_X1 U622 ( .A1(n559), .A2(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(G176GAT), .B(n558), .ZN(G1349GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n563) );
  INV_X1 U627 ( .A(n559), .ZN(n561) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(n564), .ZN(G1351GAT) );
  NOR2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n579) );
  NAND2_X1 U632 ( .A1(n579), .A2(n567), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n568), .B(KEYINPUT60), .ZN(n569) );
  XOR2_X1 U634 ( .A(n569), .B(KEYINPUT124), .Z(n571) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n574) );
  NAND2_X1 U638 ( .A1(n579), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  XOR2_X1 U640 ( .A(G211GAT), .B(KEYINPUT125), .Z(n577) );
  NAND2_X1 U641 ( .A1(n579), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1354GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n581) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XOR2_X1 U646 ( .A(G218GAT), .B(n582), .Z(G1355GAT) );
endmodule

