//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945;
  XOR2_X1   g000(.A(G197gat), .B(G204gat), .Z(new_n202));
  XOR2_X1   g001(.A(KEYINPUT76), .B(G211gat), .Z(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G218gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT22), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n202), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G211gat), .B(G218gat), .Z(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G226gat), .A2(G233gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT64), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(G169gat), .A3(G176gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT26), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT68), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT68), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n219), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n215), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT69), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n216), .A2(new_n217), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT69), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n215), .A2(new_n218), .A3(new_n224), .A4(new_n220), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n222), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT28), .ZN(new_n229));
  AND3_X1   g028(.A1(KEYINPUT65), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT27), .ZN(new_n231));
  NOR2_X1   g030(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n232));
  NOR3_X1   g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n234));
  INV_X1    g033(.A(G190gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n229), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT27), .B(G183gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(KEYINPUT28), .A3(new_n235), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n228), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n226), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n242));
  INV_X1    g041(.A(G183gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(new_n235), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AND3_X1   g047(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n244), .A2(KEYINPUT66), .A3(new_n235), .A4(new_n245), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n248), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  OR2_X1    g052(.A1(new_n216), .A2(KEYINPUT23), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n216), .A2(KEYINPUT23), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n254), .A2(new_n215), .A3(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n253), .A2(KEYINPUT25), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT25), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n254), .A2(new_n215), .A3(new_n255), .ZN(new_n259));
  NOR2_X1   g058(.A1(G183gat), .A2(G190gat), .ZN(new_n260));
  NOR3_X1   g059(.A1(new_n249), .A2(new_n250), .A3(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n258), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n241), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT29), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n210), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT77), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n241), .A2(new_n263), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n267), .B1(new_n241), .B2(new_n263), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n210), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT79), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI211_X1 g071(.A(KEYINPUT79), .B(new_n210), .C1(new_n268), .C2(new_n269), .ZN(new_n273));
  AOI211_X1 g072(.A(new_n208), .B(new_n266), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n264), .A2(KEYINPUT77), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n241), .A2(new_n263), .A3(new_n267), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT29), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT78), .B1(new_n277), .B2(new_n210), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n264), .A2(new_n210), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n265), .B1(new_n268), .B2(new_n269), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT78), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(new_n281), .A3(new_n209), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n278), .A2(new_n279), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n274), .B1(new_n208), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G8gat), .B(G36gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(G64gat), .B(G92gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n284), .A2(KEYINPUT30), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n283), .A2(new_n208), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n266), .B1(new_n272), .B2(new_n273), .ZN(new_n291));
  INV_X1    g090(.A(new_n208), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n290), .A2(new_n293), .A3(new_n288), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT30), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G1gat), .B(G29gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n298), .B(G85gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT0), .B(G57gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G225gat), .A2(G233gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G120gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G113gat), .ZN(new_n305));
  INV_X1    g104(.A(G113gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G120gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT1), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(G127gat), .A2(G134gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G127gat), .A2(G134gat), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n312), .A2(new_n313), .B1(KEYINPUT70), .B2(new_n309), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n309), .A2(KEYINPUT70), .ZN(new_n316));
  INV_X1    g115(.A(new_n313), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n316), .B1(new_n317), .B2(new_n311), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n318), .A2(new_n309), .A3(new_n308), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G155gat), .B(G162gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G148gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G141gat), .ZN(new_n324));
  INV_X1    g123(.A(G141gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G148gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT80), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT2), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT80), .B1(new_n324), .B2(new_n326), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n322), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n324), .A2(new_n326), .ZN(new_n332));
  INV_X1    g131(.A(G162gat), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT2), .B1(new_n333), .B2(KEYINPUT81), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n332), .A2(new_n321), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n331), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT80), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n340), .A2(new_n328), .A3(new_n327), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n335), .B1(new_n341), .B2(new_n322), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n342), .A2(new_n320), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n303), .B1(new_n338), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT5), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n337), .A2(KEYINPUT82), .A3(KEYINPUT4), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n342), .A2(new_n348), .A3(new_n320), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n348), .B1(new_n342), .B2(new_n320), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n349), .B1(new_n350), .B2(KEYINPUT82), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n303), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n331), .A2(new_n336), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT3), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT3), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n342), .A2(new_n355), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n315), .A2(new_n319), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n354), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n345), .B1(new_n352), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n337), .A2(KEYINPUT4), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n349), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n358), .ZN(new_n362));
  OR2_X1    g161(.A1(new_n303), .A2(KEYINPUT5), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n301), .B1(new_n359), .B2(new_n364), .ZN(new_n365));
  OR2_X1    g164(.A1(new_n365), .A2(KEYINPUT83), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(KEYINPUT83), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n347), .A2(new_n351), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n368), .A2(new_n302), .A3(new_n358), .ZN(new_n369));
  INV_X1    g168(.A(new_n345), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n364), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n301), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT6), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n366), .A2(new_n367), .A3(new_n373), .ZN(new_n374));
  OAI211_X1 g173(.A(KEYINPUT6), .B(new_n301), .C1(new_n359), .C2(new_n364), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n290), .A2(new_n293), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n287), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n297), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n355), .B1(new_n208), .B2(KEYINPUT29), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(new_n353), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n356), .A2(new_n265), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n208), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(G50gat), .ZN(new_n385));
  INV_X1    g184(.A(G50gat), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n381), .A2(new_n386), .A3(new_n383), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT31), .B(G22gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(G228gat), .A2(G233gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n391), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n385), .A2(new_n387), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G78gat), .B(G106gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n392), .A2(new_n396), .A3(new_n394), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n379), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n264), .A2(new_n320), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n241), .A2(new_n263), .A3(new_n357), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(G227gat), .ZN(new_n406));
  INV_X1    g205(.A(G233gat), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT74), .ZN(new_n409));
  OR3_X1    g208(.A1(new_n408), .A2(new_n409), .A3(KEYINPUT34), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(KEYINPUT34), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n409), .B1(new_n408), .B2(KEYINPUT34), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n406), .A2(new_n407), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n403), .A2(new_n415), .A3(new_n404), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT71), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n403), .A2(KEYINPUT71), .A3(new_n415), .A4(new_n404), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT32), .ZN(new_n421));
  XNOR2_X1  g220(.A(G71gat), .B(G99gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(G43gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT72), .B(G15gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  AOI21_X1  g224(.A(new_n421), .B1(KEYINPUT33), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT33), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n420), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n421), .A2(new_n428), .A3(new_n425), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT73), .ZN(new_n430));
  INV_X1    g229(.A(new_n425), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n431), .B1(new_n420), .B2(KEYINPUT32), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT73), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n428), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n426), .B1(new_n430), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n414), .B1(new_n435), .B2(KEYINPUT75), .ZN(new_n436));
  INV_X1    g235(.A(new_n426), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n432), .A2(new_n433), .A3(new_n428), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n433), .B1(new_n432), .B2(new_n428), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT75), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n441), .A3(new_n413), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n436), .A2(KEYINPUT36), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n440), .A2(new_n414), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT36), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n437), .B(new_n413), .C1(new_n438), .C2(new_n439), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n301), .B(KEYINPUT84), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT88), .B1(new_n371), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT88), .ZN(new_n451));
  INV_X1    g250(.A(new_n449), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n451), .B(new_n452), .C1(new_n359), .C2(new_n364), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n373), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n455), .A2(new_n375), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n294), .ZN(new_n457));
  AOI211_X1 g256(.A(new_n292), .B(new_n266), .C1(new_n272), .C2(new_n273), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n458), .B1(new_n292), .B2(new_n283), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n288), .B1(new_n459), .B2(KEYINPUT37), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT37), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT89), .B1(new_n284), .B2(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n290), .A2(KEYINPUT89), .A3(new_n461), .A4(new_n293), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n460), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT38), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT89), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n468), .B1(new_n377), .B2(KEYINPUT37), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n463), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n461), .B1(new_n290), .B2(new_n293), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT90), .B1(new_n471), .B2(new_n288), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT90), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n473), .B(new_n287), .C1(new_n284), .C2(new_n461), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n470), .A2(KEYINPUT38), .A3(new_n472), .A4(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n457), .B1(new_n467), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n289), .A2(new_n296), .A3(new_n378), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n362), .A2(new_n303), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n449), .B1(new_n478), .B2(KEYINPUT39), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT85), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n338), .A2(new_n343), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT39), .B1(new_n482), .B2(new_n303), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT86), .ZN(new_n484));
  OR2_X1    g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n484), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(new_n478), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n479), .A2(new_n480), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n481), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT40), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n450), .B2(new_n453), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n490), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n493), .A2(KEYINPUT87), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(KEYINPUT87), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n477), .B(new_n492), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n400), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n402), .B(new_n448), .C1(new_n476), .C2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n436), .A2(new_n400), .A3(new_n442), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT35), .B1(new_n499), .B2(new_n379), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT91), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n455), .A2(new_n375), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n297), .A2(new_n501), .A3(new_n502), .A4(new_n378), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n401), .B1(new_n444), .B2(new_n446), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT91), .B1(new_n477), .B2(new_n456), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT35), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n503), .A2(new_n504), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n500), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n498), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G43gat), .B(G50gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n510), .A2(KEYINPUT15), .ZN(new_n511));
  XNOR2_X1  g310(.A(KEYINPUT94), .B(G36gat), .ZN(new_n512));
  INV_X1    g311(.A(G29gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(G29gat), .A2(G36gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT14), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n511), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n510), .A2(KEYINPUT15), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n518), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT17), .ZN(new_n522));
  INV_X1    g321(.A(G8gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT16), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n524), .B1(new_n525), .B2(G1gat), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n523), .B1(new_n526), .B2(KEYINPUT95), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n526), .B1(G1gat), .B2(new_n524), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI221_X1 g328(.A(new_n526), .B1(KEYINPUT95), .B2(new_n523), .C1(G1gat), .C2(new_n524), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n519), .A2(new_n520), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n522), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n521), .A2(new_n531), .ZN(new_n536));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n535), .A2(KEYINPUT18), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n538), .B(KEYINPUT97), .Z(new_n539));
  XOR2_X1   g338(.A(G169gat), .B(G197gat), .Z(new_n540));
  XNOR2_X1  g339(.A(G113gat), .B(G141gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(KEYINPUT92), .B(KEYINPUT11), .Z(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT93), .B(KEYINPUT12), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n521), .B(new_n531), .ZN(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT98), .B(KEYINPUT13), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(new_n537), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT96), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT18), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n535), .A2(KEYINPUT96), .A3(new_n536), .A4(new_n537), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n539), .A2(new_n547), .A3(new_n551), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n551), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n538), .B(KEYINPUT97), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n546), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n558), .A2(new_n561), .A3(KEYINPUT99), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT99), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n563), .B(new_n546), .C1(new_n559), .C2(new_n560), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT21), .ZN(new_n567));
  XNOR2_X1  g366(.A(G57gat), .B(G64gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT9), .ZN(new_n569));
  INV_X1    g368(.A(G71gat), .ZN(new_n570));
  INV_X1    g369(.A(G78gat), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n568), .B1(KEYINPUT100), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G71gat), .B(G78gat), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n573), .B(new_n574), .C1(KEYINPUT100), .C2(new_n572), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n568), .A2(new_n569), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n576), .A2(new_n574), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n531), .B1(new_n567), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(G183gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n578), .A2(new_n567), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n583), .B(KEYINPUT101), .Z(new_n584));
  XNOR2_X1  g383(.A(new_n582), .B(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G127gat), .B(G155gat), .Z(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT102), .B(KEYINPUT20), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(G211gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT19), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n585), .A2(new_n586), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n585), .A2(new_n586), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n590), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G85gat), .A2(G92gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT7), .ZN(new_n598));
  INV_X1    g397(.A(G99gat), .ZN(new_n599));
  INV_X1    g398(.A(G106gat), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT8), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n598), .B(new_n601), .C1(G85gat), .C2(G92gat), .ZN(new_n602));
  XOR2_X1   g401(.A(G99gat), .B(G106gat), .Z(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT105), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n602), .A2(new_n603), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n606), .A2(KEYINPUT104), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(KEYINPUT104), .ZN(new_n608));
  OR3_X1    g407(.A1(new_n605), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(new_n522), .A3(new_n534), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n606), .B(KEYINPUT104), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(new_n605), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n532), .ZN(new_n613));
  XOR2_X1   g412(.A(G190gat), .B(G218gat), .Z(new_n614));
  NAND2_X1  g413(.A1(G232gat), .A2(G233gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n615), .B(KEYINPUT103), .Z(new_n616));
  INV_X1    g415(.A(KEYINPUT41), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n610), .A2(new_n613), .A3(new_n614), .A4(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT106), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n616), .A2(new_n617), .ZN(new_n622));
  XOR2_X1   g421(.A(G134gat), .B(G162gat), .Z(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n610), .A2(new_n613), .A3(new_n618), .ZN(new_n626));
  INV_X1    g425(.A(new_n614), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n619), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n625), .B(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n578), .B1(new_n611), .B2(new_n605), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT10), .ZN(new_n632));
  INV_X1    g431(.A(new_n578), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n633), .A2(new_n606), .A3(new_n604), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n612), .A2(KEYINPUT10), .A3(new_n633), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(G230gat), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n407), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G120gat), .B(G148gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(G176gat), .B(G204gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n631), .A2(new_n634), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n641), .B(new_n645), .C1(new_n640), .C2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT107), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n646), .A2(new_n640), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n639), .B1(new_n635), .B2(new_n636), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n644), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n649), .B(new_n652), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n596), .A2(new_n630), .A3(new_n653), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n509), .A2(new_n566), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n376), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n477), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT16), .B(G8gat), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n661), .B(KEYINPUT42), .Z(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(G8gat), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(G1325gat));
  NAND2_X1  g463(.A1(new_n444), .A2(new_n446), .ZN(new_n665));
  AOI21_X1  g464(.A(G15gat), .B1(new_n655), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n448), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(G15gat), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(KEYINPUT108), .Z(new_n669));
  AOI21_X1  g468(.A(new_n666), .B1(new_n655), .B2(new_n669), .ZN(G1326gat));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n401), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT43), .B(G22gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1327gat));
  INV_X1    g472(.A(new_n630), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n674), .B1(new_n498), .B2(new_n508), .ZN(new_n675));
  INV_X1    g474(.A(new_n596), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n676), .A2(new_n565), .A3(new_n653), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n678), .A2(new_n513), .A3(new_n656), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT45), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n681), .B1(new_n509), .B2(new_n630), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n630), .B(KEYINPUT110), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n685));
  AOI211_X1 g484(.A(new_n684), .B(new_n685), .C1(new_n498), .C2(new_n508), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n677), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n687), .A2(new_n376), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n680), .B1(new_n689), .B2(new_n513), .ZN(G1328gat));
  NAND3_X1  g489(.A1(new_n678), .A2(new_n512), .A3(new_n477), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n691), .B(KEYINPUT46), .Z(new_n692));
  INV_X1    g491(.A(new_n477), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n687), .A2(new_n693), .A3(new_n688), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n512), .B2(new_n694), .ZN(G1329gat));
  INV_X1    g494(.A(G43gat), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n678), .A2(new_n696), .A3(new_n665), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n687), .A2(new_n688), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n667), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n697), .B1(new_n699), .B2(G43gat), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT47), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT111), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n697), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n700), .B(new_n703), .ZN(G1330gat));
  AND4_X1   g503(.A1(new_n386), .A2(new_n675), .A3(new_n401), .A4(new_n677), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n401), .B(new_n677), .C1(new_n682), .C2(new_n686), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n705), .B1(new_n706), .B2(G50gat), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT48), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT112), .ZN(new_n709));
  AOI211_X1 g508(.A(new_n709), .B(new_n705), .C1(new_n706), .C2(G50gat), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n706), .A2(new_n709), .A3(G50gat), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT48), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n708), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(KEYINPUT113), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT113), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n716), .B(new_n708), .C1(new_n710), .C2(new_n713), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(G1331gat));
  NOR2_X1   g517(.A1(new_n596), .A2(new_n630), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n509), .A2(new_n565), .A3(new_n719), .A4(new_n653), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n720), .A2(KEYINPUT114), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(KEYINPUT114), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n656), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g525(.A1(new_n723), .A2(new_n693), .ZN(new_n727));
  NOR2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  AND2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n727), .B2(new_n728), .ZN(G1333gat));
  NAND3_X1  g530(.A1(new_n724), .A2(G71gat), .A3(new_n667), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n665), .B(KEYINPUT115), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n570), .B1(new_n723), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n732), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n735), .B1(new_n732), .B2(new_n734), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(G1334gat));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n400), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(new_n571), .ZN(G1335gat));
  NOR2_X1   g539(.A1(new_n676), .A2(new_n566), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n653), .B(new_n741), .C1(new_n682), .C2(new_n686), .ZN(new_n742));
  INV_X1    g541(.A(G85gat), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n742), .A2(new_n743), .A3(new_n376), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n509), .A2(new_n630), .A3(new_n741), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(KEYINPUT51), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n675), .B2(new_n741), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n653), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n656), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n744), .B1(new_n752), .B2(new_n743), .ZN(G1336gat));
  OAI21_X1  g552(.A(G92gat), .B1(new_n742), .B2(new_n693), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT52), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n693), .A2(G92gat), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n754), .B(new_n755), .C1(new_n750), .C2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT118), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n745), .A2(KEYINPUT117), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(new_n746), .B2(new_n748), .ZN(new_n760));
  INV_X1    g559(.A(new_n653), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n745), .A2(KEYINPUT117), .A3(new_n747), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n760), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n754), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n758), .B1(new_n765), .B2(KEYINPUT52), .ZN(new_n766));
  AOI211_X1 g565(.A(KEYINPUT118), .B(new_n755), .C1(new_n764), .C2(new_n754), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n757), .B1(new_n766), .B2(new_n767), .ZN(G1337gat));
  NAND3_X1  g567(.A1(new_n751), .A2(new_n599), .A3(new_n665), .ZN(new_n769));
  OAI21_X1  g568(.A(G99gat), .B1(new_n742), .B2(new_n448), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1338gat));
  NOR2_X1   g570(.A1(new_n742), .A2(new_n400), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n600), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n761), .A2(G106gat), .A3(new_n400), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n760), .A2(new_n763), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT53), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n749), .A2(new_n774), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n776), .B1(new_n773), .B2(new_n779), .ZN(G1339gat));
  NAND3_X1  g579(.A1(new_n635), .A2(new_n639), .A3(new_n636), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n641), .A2(KEYINPUT54), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n645), .B1(new_n651), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n782), .A2(KEYINPUT55), .A3(new_n784), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(new_n647), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT119), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT119), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n787), .A2(new_n791), .A3(new_n647), .A4(new_n788), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n565), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n548), .A2(new_n550), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n537), .B1(new_n535), .B2(new_n536), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n544), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n558), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n653), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n684), .B1(new_n793), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n790), .A2(new_n792), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n683), .A2(new_n802), .A3(new_n798), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n676), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  NOR4_X1   g603(.A1(new_n596), .A2(new_n566), .A3(new_n630), .A4(new_n653), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n806), .A2(new_n376), .A3(new_n499), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n807), .A2(new_n693), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n808), .A2(new_n306), .A3(new_n566), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n802), .A2(new_n566), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n683), .B1(new_n810), .B2(new_n799), .ZN(new_n811));
  INV_X1    g610(.A(new_n803), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n596), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n805), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n815), .A2(new_n656), .A3(new_n693), .A4(new_n504), .ZN(new_n816));
  OAI21_X1  g615(.A(G113gat), .B1(new_n816), .B2(new_n565), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n809), .A2(new_n817), .ZN(G1340gat));
  NAND3_X1  g617(.A1(new_n808), .A2(new_n304), .A3(new_n653), .ZN(new_n819));
  OAI21_X1  g618(.A(G120gat), .B1(new_n816), .B2(new_n761), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(G1341gat));
  INV_X1    g620(.A(G127gat), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n816), .A2(new_n822), .A3(new_n596), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n676), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n823), .B1(new_n824), .B2(new_n822), .ZN(G1342gat));
  INV_X1    g624(.A(G134gat), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n674), .A2(new_n477), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n807), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n828), .A2(KEYINPUT56), .ZN(new_n829));
  OAI21_X1  g628(.A(G134gat), .B1(new_n816), .B2(new_n674), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(KEYINPUT56), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(G1343gat));
  AND2_X1   g631(.A1(new_n787), .A2(new_n788), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n833), .A2(new_n562), .A3(new_n564), .A4(new_n647), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n630), .B1(new_n834), .B2(new_n799), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n596), .B1(new_n812), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n814), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT57), .B1(new_n837), .B2(new_n400), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n815), .A2(new_n839), .A3(new_n401), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n667), .A2(new_n376), .A3(new_n477), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G141gat), .B1(new_n842), .B2(new_n565), .ZN(new_n843));
  NOR4_X1   g642(.A1(new_n806), .A2(new_n376), .A3(new_n400), .A4(new_n667), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n565), .A2(G141gat), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT120), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n693), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT58), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n843), .A2(new_n850), .A3(new_n847), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(G1344gat));
  AND2_X1   g651(.A1(new_n844), .A2(new_n693), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n853), .A2(KEYINPUT121), .A3(new_n323), .A4(new_n653), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n844), .A2(new_n653), .A3(new_n693), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(G148gat), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(new_n859));
  AOI211_X1 g658(.A(KEYINPUT59), .B(new_n323), .C1(new_n859), .C2(new_n653), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861));
  OAI211_X1 g660(.A(KEYINPUT57), .B(new_n401), .C1(new_n804), .C2(new_n805), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n815), .A2(KEYINPUT122), .A3(KEYINPUT57), .A4(new_n401), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n674), .A2(new_n789), .A3(new_n797), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n835), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n805), .B1(new_n596), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n839), .B1(new_n868), .B2(new_n400), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n864), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n653), .A3(new_n841), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n861), .B1(new_n871), .B2(G148gat), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n858), .B1(new_n860), .B2(new_n872), .ZN(G1345gat));
  AOI21_X1  g672(.A(G155gat), .B1(new_n853), .B2(new_n676), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n676), .A2(G155gat), .ZN(new_n875));
  XOR2_X1   g674(.A(new_n875), .B(KEYINPUT123), .Z(new_n876));
  AOI21_X1  g675(.A(new_n874), .B1(new_n859), .B2(new_n876), .ZN(G1346gat));
  XOR2_X1   g676(.A(KEYINPUT81), .B(G162gat), .Z(new_n878));
  OAI21_X1  g677(.A(new_n878), .B1(new_n842), .B2(new_n684), .ZN(new_n879));
  INV_X1    g678(.A(new_n878), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n844), .A2(new_n880), .A3(new_n827), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(G1347gat));
  NOR2_X1   g681(.A1(new_n693), .A2(new_n656), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n813), .B2(new_n814), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n436), .A2(new_n442), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n885), .A2(new_n400), .A3(new_n887), .ZN(new_n888));
  OR3_X1    g687(.A1(new_n888), .A2(G169gat), .A3(new_n565), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n400), .B(new_n883), .C1(new_n804), .C2(new_n805), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n733), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(G169gat), .B1(new_n893), .B2(new_n565), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n889), .A2(new_n894), .ZN(G1348gat));
  NAND4_X1  g694(.A1(new_n891), .A2(G176gat), .A3(new_n653), .A4(new_n892), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT124), .ZN(new_n897));
  INV_X1    g696(.A(new_n888), .ZN(new_n898));
  AOI21_X1  g697(.A(G176gat), .B1(new_n898), .B2(new_n653), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n897), .A2(new_n899), .ZN(G1349gat));
  NAND2_X1  g699(.A1(new_n244), .A2(new_n245), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n901), .B1(new_n893), .B2(new_n596), .ZN(new_n902));
  INV_X1    g701(.A(new_n238), .ZN(new_n903));
  NOR4_X1   g702(.A1(new_n888), .A2(KEYINPUT125), .A3(new_n596), .A4(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n890), .A2(new_n903), .A3(new_n886), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n905), .B1(new_n906), .B2(new_n676), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n902), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT60), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT60), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n910), .B(new_n902), .C1(new_n904), .C2(new_n907), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(G1350gat));
  NAND3_X1  g711(.A1(new_n898), .A2(new_n235), .A3(new_n683), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n885), .A2(new_n630), .A3(new_n400), .A4(new_n892), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n914), .A2(new_n915), .A3(G190gat), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n914), .B2(G190gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT126), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g719(.A(KEYINPUT126), .B(new_n913), .C1(new_n916), .C2(new_n917), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1351gat));
  NOR2_X1   g721(.A1(new_n667), .A2(new_n884), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n870), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(G197gat), .B1(new_n924), .B2(new_n565), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n806), .A2(new_n400), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n923), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n927), .A2(G197gat), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n925), .B1(new_n565), .B2(new_n928), .ZN(G1352gat));
  NOR3_X1   g728(.A1(new_n927), .A2(G204gat), .A3(new_n761), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT62), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n870), .A2(new_n653), .A3(new_n923), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(G204gat), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1353gat));
  NAND3_X1  g733(.A1(new_n870), .A2(new_n676), .A3(new_n923), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G211gat), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT63), .ZN(new_n937));
  INV_X1    g736(.A(new_n203), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n926), .A2(new_n676), .A3(new_n938), .A4(new_n923), .ZN(new_n939));
  XOR2_X1   g738(.A(new_n939), .B(KEYINPUT127), .Z(new_n940));
  INV_X1    g739(.A(KEYINPUT63), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n935), .A2(new_n941), .A3(G211gat), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n937), .A2(new_n940), .A3(new_n942), .ZN(G1354gat));
  OAI21_X1  g742(.A(G218gat), .B1(new_n924), .B2(new_n674), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n927), .A2(G218gat), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n684), .B2(new_n945), .ZN(G1355gat));
endmodule


