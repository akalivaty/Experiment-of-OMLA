//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n541, new_n542, new_n543, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n610, new_n612,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160,
    new_n1161, new_n1163, new_n1164;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT68), .ZN(G261));
  AOI22_X1  g032(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G137), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT69), .B(G2105), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n461), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  XOR2_X1   g042(.A(KEYINPUT3), .B(G2104), .Z(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n466), .B1(new_n470), .B2(new_n465), .ZN(G160));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n462), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n468), .A2(new_n464), .ZN(new_n475));
  AOI22_X1  g050(.A1(G136), .A2(new_n474), .B1(new_n475), .B2(G124), .ZN(new_n476));
  OAI221_X1 g051(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n464), .C2(G112), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(G162));
  NAND3_X1  g053(.A1(new_n462), .A2(new_n464), .A3(G138), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n482));
  INV_X1    g057(.A(G114), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  NOR3_X1   g059(.A1(new_n472), .A2(KEYINPUT70), .A3(G114), .ZN(new_n485));
  OAI221_X1 g060(.A(G2104), .B1(G102), .B2(G2105), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n462), .A2(new_n464), .A3(KEYINPUT4), .A4(G138), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n462), .A2(G126), .A3(G2105), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n481), .A2(new_n486), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G164));
  NAND2_X1  g065(.A1(G75), .A2(G543), .ZN(new_n491));
  AND2_X1   g066(.A1(KEYINPUT5), .A2(G543), .ZN(new_n492));
  NOR2_X1   g067(.A1(KEYINPUT5), .A2(G543), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G62), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  OR2_X1    g072(.A1(KEYINPUT6), .A2(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT6), .A2(G651), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n496), .A2(G651), .B1(G50), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  OAI22_X1  g078(.A1(new_n502), .A2(new_n503), .B1(new_n492), .B2(new_n493), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT71), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n498), .A2(new_n499), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT5), .B(G543), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n505), .A2(G88), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n501), .A2(new_n510), .ZN(G303));
  INV_X1    g086(.A(G303), .ZN(G166));
  XOR2_X1   g087(.A(KEYINPUT72), .B(KEYINPUT7), .Z(new_n513));
  NAND3_X1  g088(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n514), .A2(new_n515), .ZN(new_n517));
  OR3_X1    g092(.A1(new_n513), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n500), .A2(G51), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n518), .A2(new_n519), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n505), .A2(G89), .A3(new_n509), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(G168));
  NAND2_X1  g099(.A1(G77), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G64), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n494), .B2(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n527), .A2(G651), .B1(G52), .B2(new_n500), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n505), .A2(G90), .A3(new_n509), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(G301));
  INV_X1    g105(.A(G301), .ZN(G171));
  NAND2_X1  g106(.A1(G68), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G56), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n494), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n534), .A2(G651), .B1(G43), .B2(new_n500), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n505), .A2(G81), .A3(new_n509), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G860), .ZN(G153));
  NAND4_X1  g114(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g115(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n541));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NAND4_X1  g118(.A1(G319), .A2(G483), .A3(G661), .A4(new_n543), .ZN(G188));
  AND3_X1   g119(.A1(new_n505), .A2(G91), .A3(new_n509), .ZN(new_n545));
  INV_X1    g120(.A(G65), .ZN(new_n546));
  OR2_X1    g121(.A1(KEYINPUT5), .A2(G543), .ZN(new_n547));
  NAND2_X1  g122(.A1(KEYINPUT5), .A2(G543), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g124(.A1(G78), .A2(G543), .ZN(new_n550));
  OAI21_X1  g125(.A(G651), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  XOR2_X1   g126(.A(KEYINPUT75), .B(KEYINPUT9), .Z(new_n552));
  NAND3_X1  g127(.A1(new_n500), .A2(new_n552), .A3(G53), .ZN(new_n553));
  NOR2_X1   g128(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n554));
  OAI21_X1  g129(.A(G543), .B1(new_n503), .B2(new_n502), .ZN(new_n555));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n551), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n545), .A2(new_n558), .ZN(G299));
  INV_X1    g134(.A(G168), .ZN(G286));
  NAND3_X1  g135(.A1(new_n505), .A2(G87), .A3(new_n509), .ZN(new_n561));
  INV_X1    g136(.A(G74), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n494), .A2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n563), .A2(G651), .B1(new_n500), .B2(G49), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT76), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n565), .B(new_n566), .ZN(G288));
  NAND2_X1  g142(.A1(G73), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G61), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n494), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n570), .A2(G651), .B1(G48), .B2(new_n500), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n505), .A2(G86), .A3(new_n509), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n573), .B1(new_n571), .B2(new_n572), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(G305));
  INV_X1    g152(.A(G651), .ZN(new_n578));
  OAI21_X1  g153(.A(G60), .B1(new_n492), .B2(new_n493), .ZN(new_n579));
  NAND2_X1  g154(.A1(G72), .A2(G543), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT78), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n581), .A2(new_n582), .B1(G47), .B2(new_n500), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n505), .A2(G85), .A3(new_n509), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G290));
  INV_X1    g161(.A(G868), .ZN(new_n587));
  NOR2_X1   g162(.A1(G301), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n505), .A2(G92), .A3(new_n509), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(KEYINPUT10), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n500), .A2(G54), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n547), .B2(new_n548), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n592), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  OAI211_X1 g172(.A(KEYINPUT79), .B(new_n595), .C1(new_n494), .C2(new_n593), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n597), .A2(G651), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n505), .A2(new_n600), .A3(G92), .A4(new_n509), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n590), .A2(new_n591), .A3(new_n599), .A4(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT80), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n588), .B1(new_n604), .B2(new_n587), .ZN(G284));
  XNOR2_X1  g180(.A(G284), .B(KEYINPUT81), .ZN(G321));
  NAND2_X1  g181(.A1(G299), .A2(new_n587), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(new_n587), .B2(G168), .ZN(G297));
  OAI21_X1  g183(.A(new_n607), .B1(new_n587), .B2(G168), .ZN(G280));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n604), .B1(new_n610), .B2(G860), .ZN(G148));
  NOR2_X1   g186(.A1(new_n538), .A2(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n604), .A2(new_n610), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT82), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g191(.A1(G135), .A2(new_n474), .B1(new_n475), .B2(G123), .ZN(new_n617));
  OAI221_X1 g192(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n464), .C2(G111), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(G2096), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n462), .A2(new_n460), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  INV_X1    g198(.A(G2100), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n620), .A2(new_n625), .A3(new_n626), .ZN(G156));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2427), .B(G2430), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(KEYINPUT14), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT83), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n629), .A2(new_n630), .ZN(new_n634));
  XOR2_X1   g209(.A(G2443), .B(G2446), .Z(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n636), .B1(new_n633), .B2(new_n634), .ZN(new_n642));
  OR3_X1    g217(.A1(new_n638), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT84), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n641), .B1(new_n638), .B2(new_n642), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n643), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  AND2_X1   g222(.A1(new_n647), .A2(G14), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n645), .B1(new_n646), .B2(new_n643), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT85), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI211_X1 g226(.A(KEYINPUT85), .B(new_n645), .C1(new_n643), .C2(new_n646), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n648), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(G2067), .B(G2678), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT86), .ZN(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  XNOR2_X1  g232(.A(G2084), .B(G2090), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT18), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT87), .B(KEYINPUT17), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n657), .B(new_n662), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n661), .B(new_n658), .C1(new_n656), .C2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n658), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n663), .A2(new_n656), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n660), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(new_n624), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT88), .B(G2096), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G227));
  XOR2_X1   g245(.A(G1971), .B(G1976), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  AND2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n673), .A2(new_n674), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n672), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n672), .B2(new_n678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT89), .Z(new_n682));
  XOR2_X1   g257(.A(G1981), .B(G1986), .Z(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n682), .B(new_n687), .ZN(G229));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G32), .ZN(new_n690));
  NAND3_X1  g265(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT26), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n465), .A2(new_n462), .ZN(new_n693));
  INV_X1    g268(.A(G129), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n472), .A2(G105), .A3(G2104), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT95), .ZN(new_n697));
  INV_X1    g272(.A(G141), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(new_n473), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n690), .B1(new_n701), .B2(new_n689), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT27), .ZN(new_n703));
  INV_X1    g278(.A(G1996), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G35), .ZN(new_n706));
  OR3_X1    g281(.A1(new_n706), .A2(KEYINPUT98), .A3(G29), .ZN(new_n707));
  OAI21_X1  g282(.A(KEYINPUT98), .B1(new_n706), .B2(G29), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n707), .B(new_n708), .C1(G162), .C2(new_n689), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT29), .B(G2090), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G5), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G171), .B2(new_n712), .ZN(new_n714));
  INV_X1    g289(.A(G1961), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(G16), .A2(G19), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n538), .B2(G16), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n711), .B(new_n716), .C1(G1341), .C2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT24), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n720), .A2(G34), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(G34), .ZN(new_n722));
  AOI21_X1  g297(.A(G29), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G160), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(G29), .ZN(new_n725));
  INV_X1    g300(.A(G2084), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT31), .B(G11), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT30), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n729), .A2(G28), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n689), .B1(new_n729), .B2(G28), .ZN(new_n731));
  OAI221_X1 g306(.A(new_n728), .B1(new_n730), .B2(new_n731), .C1(new_n619), .C2(new_n689), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n689), .A2(G26), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT28), .Z(new_n735));
  AOI22_X1  g310(.A1(G140), .A2(new_n474), .B1(new_n475), .B2(G128), .ZN(new_n736));
  OAI221_X1 g311(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n464), .C2(G116), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n735), .B1(new_n738), .B2(G29), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G2067), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n718), .A2(G1341), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n733), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT99), .B(KEYINPUT23), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n712), .A2(G20), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G299), .B2(G16), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(G1956), .Z(new_n747));
  NOR4_X1   g322(.A1(new_n705), .A2(new_n719), .A3(new_n742), .A4(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(G4), .A2(G16), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n604), .B2(G16), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT93), .B(G1348), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n712), .A2(G21), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G168), .B2(new_n712), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT96), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT97), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n756), .B2(G1966), .ZN(new_n757));
  INV_X1    g332(.A(G1966), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n758), .A2(KEYINPUT97), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n757), .B(new_n759), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n689), .A2(G33), .ZN(new_n761));
  NAND2_X1  g336(.A1(G115), .A2(G2104), .ZN(new_n762));
  INV_X1    g337(.A(G127), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n468), .B2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT94), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n464), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n765), .B2(new_n764), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n474), .A2(G139), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT25), .Z(new_n770));
  NAND3_X1  g345(.A1(new_n767), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n761), .B1(new_n771), .B2(G29), .ZN(new_n772));
  INV_X1    g347(.A(G2072), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n689), .A2(G27), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G164), .B2(new_n689), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G2078), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n774), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n748), .A2(new_n752), .A3(new_n760), .A4(new_n779), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n712), .A2(G6), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G305), .B2(G16), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT32), .B(G1981), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  MUX2_X1   g360(.A(G23), .B(new_n565), .S(G16), .Z(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT33), .B(G1976), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n782), .A2(new_n784), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n712), .A2(G22), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G166), .B2(new_n712), .ZN(new_n791));
  INV_X1    g366(.A(G1971), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n785), .A2(new_n788), .A3(new_n789), .A4(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT91), .B(KEYINPUT34), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  NOR2_X1   g372(.A1(G25), .A2(G29), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n474), .A2(G131), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n475), .A2(G119), .ZN(new_n800));
  OAI221_X1 g375(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n464), .C2(G107), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n798), .B1(new_n803), .B2(G29), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT35), .B(G1991), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT90), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n804), .B(new_n806), .Z(new_n807));
  OR2_X1    g382(.A1(G16), .A2(G24), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G290), .B2(new_n712), .ZN(new_n809));
  INV_X1    g384(.A(G1986), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  NOR4_X1   g387(.A1(new_n807), .A2(new_n811), .A3(new_n812), .A4(KEYINPUT92), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n796), .A2(new_n797), .A3(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT36), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n780), .A2(new_n816), .A3(new_n817), .ZN(G311));
  INV_X1    g393(.A(G311), .ZN(G150));
  NAND2_X1  g394(.A1(new_n604), .A2(G559), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT38), .Z(new_n821));
  NAND2_X1  g396(.A1(new_n537), .A2(KEYINPUT102), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT102), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n535), .A2(new_n536), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT100), .B1(new_n826), .B2(new_n578), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT101), .B(G93), .Z(new_n828));
  NAND3_X1  g403(.A1(new_n505), .A2(new_n509), .A3(new_n828), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n507), .A2(G67), .ZN(new_n831));
  NAND2_X1  g406(.A1(G80), .A2(G543), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n578), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT100), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n833), .A2(new_n834), .B1(G55), .B2(new_n500), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n830), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n825), .A2(new_n836), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n822), .A2(new_n824), .B1(new_n830), .B2(new_n835), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n821), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n842));
  AOI21_X1  g417(.A(G860), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n841), .A2(KEYINPUT103), .A3(new_n842), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT103), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n821), .B(new_n839), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n845), .B1(new_n846), .B2(KEYINPUT39), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n843), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n836), .A2(G860), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT104), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT37), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n851), .ZN(G145));
  INV_X1    g427(.A(KEYINPUT108), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n700), .B(new_n489), .ZN(new_n854));
  INV_X1    g429(.A(G118), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT107), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n465), .A2(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n856), .B2(new_n857), .ZN(new_n859));
  INV_X1    g434(.A(G130), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n859), .B1(new_n693), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n474), .A2(G142), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT106), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n862), .A2(KEYINPUT106), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n854), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n854), .A2(new_n865), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n738), .A2(KEYINPUT105), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT105), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n736), .A2(new_n870), .A3(new_n737), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(new_n771), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n872), .A2(new_n771), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n802), .B(new_n622), .ZN(new_n876));
  NOR3_X1   g451(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n876), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n872), .A2(new_n771), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n878), .B1(new_n879), .B2(new_n873), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n868), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n724), .B(new_n619), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(G162), .Z(new_n883));
  OAI21_X1  g458(.A(new_n876), .B1(new_n874), .B2(new_n875), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n879), .A2(new_n873), .A3(new_n878), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n884), .A2(new_n885), .A3(new_n866), .A4(new_n867), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n881), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n883), .B1(new_n881), .B2(new_n886), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n853), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n890), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n892), .A2(KEYINPUT108), .A3(new_n888), .A4(new_n887), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g469(.A(KEYINPUT109), .B(KEYINPUT40), .Z(new_n895));
  XNOR2_X1  g470(.A(new_n894), .B(new_n895), .ZN(G395));
  NAND2_X1  g471(.A1(new_n602), .A2(G299), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n545), .A2(new_n558), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n596), .B1(new_n507), .B2(G66), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n578), .B1(new_n899), .B2(KEYINPUT79), .ZN(new_n900));
  AOI22_X1  g475(.A1(new_n900), .A2(new_n597), .B1(G54), .B2(new_n500), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n898), .A2(new_n901), .A3(new_n590), .A4(new_n601), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n613), .A2(new_n839), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n613), .A2(new_n839), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n897), .A2(new_n902), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT111), .B1(new_n908), .B2(KEYINPUT41), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(KEYINPUT41), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n897), .A2(new_n902), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n909), .B1(new_n913), .B2(KEYINPUT111), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n906), .B(KEYINPUT110), .C1(new_n907), .C2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n576), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT112), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n501), .A2(new_n510), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n917), .B1(new_n501), .B2(new_n510), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n916), .B(new_n574), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n920), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n922), .B(new_n918), .C1(new_n575), .C2(new_n576), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT113), .ZN(new_n925));
  AND2_X1   g500(.A1(G290), .A2(new_n565), .ZN(new_n926));
  NOR2_X1   g501(.A1(G290), .A2(new_n565), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OR2_X1    g503(.A1(G290), .A2(new_n565), .ZN(new_n929));
  NAND2_X1  g504(.A1(G290), .A2(new_n565), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(KEYINPUT113), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n924), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT113), .B1(new_n929), .B2(new_n930), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(new_n921), .A3(new_n923), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT42), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n906), .A2(KEYINPUT110), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n915), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n936), .B1(new_n915), .B2(new_n937), .ZN(new_n939));
  OAI21_X1  g514(.A(G868), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n835), .A2(new_n827), .A3(new_n829), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n940), .B1(G868), .B2(new_n941), .ZN(G295));
  OAI21_X1  g517(.A(new_n940), .B1(G868), .B2(new_n941), .ZN(G331));
  AND3_X1   g518(.A1(new_n897), .A2(new_n911), .A3(new_n902), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n911), .B1(new_n897), .B2(new_n902), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT111), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT111), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(new_n903), .B2(new_n911), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n825), .A2(new_n836), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n941), .A2(new_n822), .A3(new_n824), .ZN(new_n950));
  NAND2_X1  g525(.A1(G168), .A2(G301), .ZN(new_n951));
  OAI21_X1  g526(.A(G171), .B1(new_n523), .B2(new_n522), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n949), .A2(new_n950), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(new_n837), .B2(new_n838), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n946), .A2(new_n948), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n953), .A3(new_n903), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n935), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n932), .A2(new_n934), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n955), .A2(new_n953), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n960), .B(new_n957), .C1(new_n914), .C2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n959), .A2(new_n963), .A3(new_n888), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n961), .A2(new_n913), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n935), .B1(new_n967), .B2(new_n958), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n968), .A2(new_n963), .A3(new_n888), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n969), .A2(new_n965), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT44), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT114), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n964), .A2(new_n972), .A3(KEYINPUT43), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n972), .B1(new_n964), .B2(KEYINPUT43), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n971), .B1(new_n976), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g552(.A(new_n466), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n470), .A2(new_n465), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n978), .A2(G40), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G1384), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n489), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n700), .B(new_n704), .ZN(new_n986));
  INV_X1    g561(.A(G2067), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n738), .B(new_n987), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n803), .A2(new_n806), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n803), .A2(new_n806), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(G290), .B(G1986), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n985), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n982), .A2(new_n983), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n489), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n995), .A2(new_n980), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n758), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n978), .A2(new_n979), .A3(G40), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n999), .B1(new_n982), .B2(KEYINPUT50), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n489), .A2(new_n1001), .A3(new_n981), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1000), .A2(new_n726), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n998), .A2(G168), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(G8), .ZN(new_n1005));
  AOI21_X1  g580(.A(G168), .B1(new_n998), .B2(new_n1003), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT51), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1004), .A2(new_n1008), .A3(G8), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT62), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n999), .B1(new_n982), .B2(new_n983), .ZN(new_n1012));
  INV_X1    g587(.A(G2078), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(new_n1013), .A3(new_n996), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n1014), .A2(new_n1015), .B1(new_n1016), .B2(new_n715), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1012), .A2(KEYINPUT53), .A3(new_n1013), .A4(new_n996), .ZN(new_n1018));
  AOI21_X1  g593(.A(G301), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(G303), .A2(G8), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1020), .B(KEYINPUT55), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1016), .A2(G2090), .ZN(new_n1023));
  AOI21_X1  g598(.A(G1971), .B1(new_n1012), .B2(new_n996), .ZN(new_n1024));
  OAI211_X1 g599(.A(G8), .B(new_n1022), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G8), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1024), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT120), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1002), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n489), .A2(KEYINPUT120), .A3(new_n1001), .A4(new_n981), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G2090), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(new_n1032), .A3(new_n1000), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1026), .B1(new_n1027), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1025), .B1(new_n1034), .B2(new_n1022), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n561), .A2(G1976), .A3(new_n564), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1036), .B(KEYINPUT116), .ZN(new_n1037));
  NAND4_X1  g612(.A1(G160), .A2(new_n489), .A3(G40), .A4(new_n981), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(new_n1039), .A3(G8), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1039), .B1(new_n1038), .B2(G8), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1037), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT52), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n982), .A2(new_n999), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT115), .B1(new_n1045), .B2(new_n1026), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n1040), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n571), .A2(new_n572), .ZN(new_n1048));
  INV_X1    g623(.A(G1981), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n570), .A2(G651), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1048), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n571), .A2(new_n572), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT118), .B1(new_n570), .B2(G651), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1054), .B1(new_n1049), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1053), .A2(new_n1056), .A3(KEYINPUT119), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT49), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1047), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT117), .B(G1976), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT52), .B1(G288), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1047), .A2(new_n1037), .A3(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1044), .A2(new_n1061), .A3(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1035), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT62), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1007), .A2(new_n1067), .A3(new_n1009), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1011), .A2(new_n1019), .A3(new_n1066), .A4(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1023), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1026), .B1(new_n1070), .B2(new_n1027), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1071), .A2(KEYINPUT121), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1021), .B1(new_n1071), .B2(KEYINPUT121), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1044), .A2(new_n1061), .A3(new_n1064), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n998), .A2(new_n1003), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1075), .A2(G8), .A3(G168), .A4(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT63), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1034), .A2(new_n1022), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT63), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1076), .A2(new_n1080), .A3(G8), .A4(G168), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1025), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(G288), .A2(G1976), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1061), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(G1981), .B2(new_n1054), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1082), .A2(new_n1075), .B1(new_n1085), .B2(new_n1047), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1069), .A2(new_n1078), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1016), .A2(new_n715), .ZN(new_n1089));
  OR2_X1    g664(.A1(new_n1013), .A2(KEYINPUT125), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1013), .A2(KEYINPUT125), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1015), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1012), .A2(new_n996), .A3(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1088), .A2(new_n1089), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT126), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1017), .A2(KEYINPUT126), .A3(new_n1093), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(G171), .A3(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1088), .A2(new_n1089), .A3(G301), .A4(new_n1018), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1099), .A2(KEYINPUT54), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1094), .A2(G171), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1102), .B1(new_n1103), .B2(new_n1019), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1101), .A2(new_n1066), .A3(new_n1010), .A4(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(G1956), .B1(new_n1031), .B2(new_n1000), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT56), .B(G2072), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1012), .A2(new_n996), .A3(new_n1107), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT122), .B(KEYINPUT57), .Z(new_n1109));
  XNOR2_X1  g684(.A(new_n898), .B(new_n1109), .ZN(new_n1110));
  OR3_X1    g685(.A1(new_n1106), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1110), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n604), .A2(KEYINPUT60), .ZN(new_n1115));
  INV_X1    g690(.A(G1348), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1016), .A2(new_n1116), .B1(new_n987), .B2(new_n1045), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n604), .A2(KEYINPUT60), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1115), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1117), .A2(KEYINPUT60), .A3(new_n604), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1113), .A2(new_n1114), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  OR3_X1    g697(.A1(new_n1106), .A2(new_n1108), .A3(KEYINPUT123), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT123), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(new_n1110), .A3(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1125), .A2(KEYINPUT61), .A3(new_n1111), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT124), .B1(new_n997), .B2(G1996), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1012), .A2(new_n1128), .A3(new_n704), .A4(new_n996), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT58), .B(G1341), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1127), .B(new_n1129), .C1(new_n1045), .C2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n538), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(KEYINPUT59), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1131), .A2(new_n1134), .A3(new_n538), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1122), .A2(new_n1126), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1111), .A2(new_n604), .A3(new_n1118), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1125), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1105), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n994), .B1(new_n1087), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n984), .B1(new_n988), .B2(new_n701), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT46), .B1(new_n984), .B2(G1996), .ZN(new_n1143));
  OR3_X1    g718(.A1(new_n984), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT47), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n984), .A2(G1986), .A3(G290), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT127), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1147), .B(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT48), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1152));
  AOI211_X1 g727(.A(new_n1151), .B(new_n1152), .C1(new_n985), .C2(new_n992), .ZN(new_n1153));
  INV_X1    g728(.A(new_n989), .ZN(new_n1154));
  OAI22_X1  g729(.A1(new_n1154), .A2(new_n990), .B1(G2067), .B2(new_n738), .ZN(new_n1155));
  AOI211_X1 g730(.A(new_n1146), .B(new_n1153), .C1(new_n985), .C2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1141), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g732(.A(G319), .ZN(new_n1159));
  NOR3_X1   g733(.A1(G227), .A2(G229), .A3(new_n1159), .ZN(new_n1160));
  NAND3_X1  g734(.A1(new_n894), .A2(new_n653), .A3(new_n1160), .ZN(new_n1161));
  NOR2_X1   g735(.A1(new_n1161), .A2(new_n976), .ZN(G308));
  AND2_X1   g736(.A1(new_n653), .A2(new_n1160), .ZN(new_n1163));
  OR2_X1    g737(.A1(new_n974), .A2(new_n975), .ZN(new_n1164));
  OAI211_X1 g738(.A(new_n894), .B(new_n1163), .C1(new_n1164), .C2(new_n973), .ZN(G225));
endmodule


