//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n557, new_n559, new_n560,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1151, new_n1152;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(new_n455), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n453), .A2(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT68), .Z(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AND3_X1   g041(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT69), .ZN(new_n467));
  AOI21_X1  g042(.A(KEYINPUT69), .B1(new_n464), .B2(new_n466), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  XOR2_X1   g045(.A(new_n470), .B(KEYINPUT70), .Z(new_n471));
  AOI21_X1  g046(.A(new_n462), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n462), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT72), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n473), .B(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  OAI21_X1  g051(.A(KEYINPUT71), .B1(new_n465), .B2(G2104), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT71), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(new_n463), .A3(KEYINPUT3), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n477), .A2(new_n479), .A3(new_n466), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n462), .A2(G137), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n472), .A2(new_n483), .ZN(G160));
  NAND3_X1  g059(.A1(new_n477), .A2(new_n479), .A3(new_n466), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT73), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n485), .B(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n487), .A2(new_n462), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n487), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  OR2_X1    g066(.A1(G100), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n489), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  INV_X1    g070(.A(KEYINPUT74), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G114), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(KEYINPUT74), .ZN(new_n499));
  OAI21_X1  g074(.A(G2105), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(G126), .A2(G2105), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n485), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G138), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n506), .A2(G2105), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n480), .A2(KEYINPUT75), .A3(new_n507), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n477), .A2(new_n479), .A3(new_n466), .A4(new_n507), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT75), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n508), .A2(KEYINPUT4), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT4), .ZN(new_n513));
  OAI211_X1 g088(.A(new_n513), .B(new_n507), .C1(new_n467), .C2(new_n468), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n505), .B1(new_n512), .B2(new_n514), .ZN(G164));
  INV_X1    g090(.A(KEYINPUT76), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n516), .B1(KEYINPUT6), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  NOR3_X1   g094(.A1(new_n519), .A2(KEYINPUT76), .A3(G651), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(G543), .A3(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G50), .ZN(new_n525));
  OR2_X1    g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n528), .B(new_n522), .C1(new_n518), .C2(new_n520), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G88), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n528), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(new_n517), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n525), .A2(new_n531), .A3(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  NAND2_X1  g110(.A1(new_n524), .A2(G51), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n528), .A2(G63), .A3(G651), .ZN(new_n537));
  XOR2_X1   g112(.A(new_n537), .B(KEYINPUT77), .Z(new_n538));
  NAND2_X1  g113(.A1(new_n530), .A2(G89), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n536), .A2(new_n538), .A3(new_n539), .A4(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  NAND2_X1  g118(.A1(new_n524), .A2(G52), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n530), .A2(G90), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n528), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n517), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(new_n524), .A2(G43), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n530), .A2(G81), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n528), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n517), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  NAND4_X1  g136(.A1(new_n521), .A2(G53), .A3(G543), .A4(new_n522), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT78), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n521), .A2(new_n564), .A3(new_n522), .A4(new_n528), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n529), .A2(KEYINPUT78), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n565), .A2(G91), .A3(new_n566), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n528), .A2(G65), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  XOR2_X1   g144(.A(new_n569), .B(KEYINPUT79), .Z(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n563), .A2(new_n567), .A3(new_n571), .ZN(G299));
  INV_X1    g147(.A(new_n528), .ZN(new_n573));
  INV_X1    g148(.A(G74), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n517), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(new_n524), .B2(G49), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n565), .A2(G87), .A3(new_n566), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(G288));
  NAND3_X1  g153(.A1(new_n565), .A2(G86), .A3(new_n566), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(KEYINPUT80), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT80), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n565), .A2(new_n566), .A3(new_n581), .A4(G86), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n573), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n524), .A2(G48), .B1(G651), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(new_n524), .A2(G47), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n530), .A2(G85), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n591), .A2(new_n517), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  INV_X1    g169(.A(G54), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n528), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n523), .A2(new_n595), .B1(new_n517), .B2(new_n596), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT81), .Z(new_n598));
  NAND2_X1  g173(.A1(new_n565), .A2(new_n566), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  OR3_X1    g175(.A1(new_n599), .A2(KEYINPUT10), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(KEYINPUT10), .B1(new_n599), .B2(new_n600), .ZN(new_n602));
  AND3_X1   g177(.A1(new_n598), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n594), .B1(new_n603), .B2(G868), .ZN(G284));
  OAI21_X1  g179(.A(new_n594), .B1(new_n603), .B2(G868), .ZN(G321));
  NAND2_X1  g180(.A1(G286), .A2(G868), .ZN(new_n606));
  INV_X1    g181(.A(G299), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(G297));
  OAI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(G280));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n603), .B1(new_n610), .B2(G860), .ZN(G148));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n554), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n598), .A2(new_n601), .A3(new_n602), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n614), .A2(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n613), .B1(new_n615), .B2(new_n612), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT82), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g193(.A(new_n475), .B1(new_n467), .B2(new_n468), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n488), .A2(G135), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n490), .A2(G123), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n462), .A2(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(G2096), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(G2096), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n622), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT83), .ZN(G156));
  XOR2_X1   g206(.A(G2451), .B(G2454), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT84), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n633), .B(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT14), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n640), .B2(new_n639), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n636), .B(new_n642), .Z(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  AND3_X1   g221(.A1(new_n645), .A2(G14), .A3(new_n646), .ZN(G401));
  NOR2_X1   g222(.A1(G2072), .A2(G2078), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n442), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT17), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT86), .ZN(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  NAND3_X1  g228(.A1(new_n650), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT87), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n653), .B(new_n651), .C1(new_n442), .C2(new_n648), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n653), .B1(new_n652), .B2(new_n649), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n652), .B2(new_n650), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n655), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT88), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  NAND3_X1  g244(.A1(new_n666), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT20), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n666), .B1(new_n668), .B2(new_n669), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n668), .A2(new_n669), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n671), .B(new_n674), .C1(new_n665), .C2(new_n673), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G229));
  INV_X1    g256(.A(G29), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G25), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n488), .A2(G131), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n490), .A2(G119), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n462), .A2(G107), .ZN(new_n686));
  OAI21_X1  g261(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n684), .B(new_n685), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT89), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n683), .B1(new_n690), .B2(new_n682), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT35), .B(G1991), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G6), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n583), .A2(new_n587), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n694), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT32), .B(G1981), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n694), .A2(G22), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G166), .B2(new_n694), .ZN(new_n701));
  INV_X1    g276(.A(G1971), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  MUX2_X1   g278(.A(G23), .B(G288), .S(G16), .Z(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT33), .B(G1976), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n699), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n707), .A2(KEYINPUT34), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(KEYINPUT34), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n694), .A2(G24), .ZN(new_n710));
  INV_X1    g285(.A(G290), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(new_n694), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(G1986), .Z(new_n713));
  NAND4_X1  g288(.A1(new_n693), .A2(new_n708), .A3(new_n709), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT36), .ZN(new_n715));
  NAND3_X1  g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT26), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n475), .A2(G105), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT95), .Z(new_n719));
  AOI211_X1 g294(.A(new_n717), .B(new_n719), .C1(G141), .C2(new_n488), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n490), .A2(G129), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT94), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n724), .A2(new_n682), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n682), .B2(G32), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT27), .B(G1996), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n682), .A2(G26), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT28), .Z(new_n731));
  OR2_X1    g306(.A1(G104), .A2(G2105), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n732), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT91), .Z(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n488), .B2(G140), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n490), .A2(G128), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n731), .B1(new_n737), .B2(G29), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G2067), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n728), .A2(new_n729), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n694), .A2(G21), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G168), .B2(new_n694), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1966), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n694), .A2(G5), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G171), .B2(new_n694), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1961), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n694), .A2(G19), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n555), .B2(new_n694), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1341), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT31), .B(G11), .Z(new_n750));
  INV_X1    g325(.A(KEYINPUT30), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n682), .B1(new_n751), .B2(G28), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(KEYINPUT96), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n753), .A2(KEYINPUT96), .B1(new_n751), .B2(G28), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n750), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n627), .B2(new_n682), .ZN(new_n757));
  NOR4_X1   g332(.A1(new_n743), .A2(new_n746), .A3(new_n749), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n682), .A2(G33), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n488), .A2(G139), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT25), .Z(new_n762));
  OAI21_X1  g337(.A(G127), .B1(new_n467), .B2(new_n468), .ZN(new_n763));
  NAND2_X1  g338(.A1(G115), .A2(G2104), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n760), .B(new_n762), .C1(new_n462), .C2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n759), .B1(new_n767), .B2(new_n682), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(G2072), .Z(new_n769));
  AND2_X1   g344(.A1(KEYINPUT24), .A2(G34), .ZN(new_n770));
  NOR2_X1   g345(.A1(KEYINPUT24), .A2(G34), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n682), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT92), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G160), .B2(G29), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n774), .A2(G2084), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT97), .Z(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(G2084), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT93), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n694), .A2(G20), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT23), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n607), .B2(new_n694), .ZN(new_n782));
  INV_X1    g357(.A(G1956), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n758), .A2(new_n769), .A3(new_n779), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(G4), .A2(G16), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT90), .Z(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n614), .B2(new_n694), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1348), .ZN(new_n789));
  INV_X1    g364(.A(G2078), .ZN(new_n790));
  NOR2_X1   g365(.A1(G27), .A2(G29), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G164), .B2(G29), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT98), .Z(new_n793));
  NAND2_X1  g368(.A1(new_n682), .A2(G35), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G162), .B2(new_n682), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT29), .Z(new_n796));
  INV_X1    g371(.A(G2090), .ZN(new_n797));
  OAI221_X1 g372(.A(new_n789), .B1(new_n790), .B2(new_n793), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n793), .A2(new_n790), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR4_X1   g376(.A1(new_n740), .A2(new_n785), .A3(new_n798), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n715), .A2(new_n802), .ZN(G150));
  INV_X1    g378(.A(G150), .ZN(G311));
  NOR2_X1   g379(.A1(new_n614), .A2(new_n610), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT38), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT99), .B(G55), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n524), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n530), .A2(G93), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n528), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(new_n517), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n554), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n554), .A2(new_n812), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n806), .B(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT39), .ZN(new_n818));
  AOI21_X1  g393(.A(G860), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n818), .B2(new_n817), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n812), .A2(G860), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT100), .B(KEYINPUT37), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(KEYINPUT101), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT101), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n820), .A2(new_n826), .A3(new_n823), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(G145));
  XOR2_X1   g403(.A(new_n627), .B(G160), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n494), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n737), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G164), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n509), .A2(new_n510), .ZN(new_n834));
  OAI21_X1  g409(.A(KEYINPUT4), .B1(new_n509), .B2(new_n510), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n514), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n505), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n737), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n833), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n724), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n723), .A2(new_n839), .A3(new_n833), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT102), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n767), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n841), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n767), .A2(new_n843), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n848));
  INV_X1    g423(.A(G118), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n848), .B1(new_n849), .B2(G2105), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(new_n488), .B2(G142), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT103), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n490), .A2(new_n852), .A3(G130), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n852), .B1(new_n490), .B2(G130), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n851), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n620), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n690), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n846), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n841), .A2(new_n858), .A3(new_n842), .A4(new_n844), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n847), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n857), .B1(new_n847), .B2(new_n859), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n831), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G37), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n847), .A2(new_n859), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n856), .B(new_n689), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n867), .A2(new_n830), .A3(new_n860), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n863), .A2(new_n864), .A3(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g445(.A(G305), .B(new_n711), .ZN(new_n871));
  XNOR2_X1  g446(.A(G166), .B(G288), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  AND2_X1   g448(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n874));
  OR3_X1    g449(.A1(new_n873), .A2(KEYINPUT105), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT105), .B1(new_n873), .B2(new_n874), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n603), .A2(new_n607), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n614), .A2(G299), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n615), .A2(new_n815), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n816), .B1(new_n614), .B2(G559), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n614), .B(new_n607), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT41), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n880), .A2(KEYINPUT41), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n881), .A2(new_n882), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n877), .A2(new_n883), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n883), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(new_n875), .A3(new_n876), .ZN(new_n892));
  NOR2_X1   g467(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n890), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n893), .B1(new_n890), .B2(new_n892), .ZN(new_n895));
  OAI21_X1  g470(.A(G868), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n812), .A2(new_n612), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(G295));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n897), .ZN(G331));
  XOR2_X1   g474(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n900));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n901));
  NOR2_X1   g476(.A1(G286), .A2(G301), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(G286), .A2(G301), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n903), .A2(new_n814), .A3(new_n813), .A4(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n904), .ZN(new_n906));
  INV_X1    g481(.A(new_n814), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n554), .A2(new_n812), .ZN(new_n908));
  OAI22_X1  g483(.A1(new_n906), .A2(new_n902), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(new_n909), .A3(KEYINPUT108), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n903), .A2(new_n904), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT108), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(new_n815), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n884), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT109), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n909), .A2(KEYINPUT107), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT107), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n911), .A2(new_n815), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(new_n919), .A3(new_n905), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n878), .A2(new_n885), .A3(new_n879), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n885), .B1(new_n878), .B2(new_n879), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n914), .A2(new_n924), .A3(new_n884), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n916), .A2(new_n923), .A3(new_n873), .A4(new_n925), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n926), .A2(new_n864), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT110), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n873), .B(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n916), .A2(new_n923), .A3(new_n925), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n901), .B1(new_n927), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n920), .A2(new_n880), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT111), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n886), .A2(new_n887), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n914), .B1(KEYINPUT111), .B2(new_n922), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n926), .B(new_n864), .C1(new_n938), .C2(new_n929), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n900), .B1(new_n933), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n927), .A2(new_n901), .A3(new_n932), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(new_n943), .A3(KEYINPUT44), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n944), .ZN(G397));
  INV_X1    g520(.A(KEYINPUT45), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(G164), .B2(G1384), .ZN(new_n947));
  NAND2_X1  g522(.A1(G160), .A2(G40), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G1996), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n723), .B(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G2067), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n737), .B(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n692), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n689), .B(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n949), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(G290), .A2(G1986), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT112), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n949), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n949), .A2(G1986), .A3(G290), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OR2_X1    g537(.A1(new_n962), .A2(KEYINPUT113), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(KEYINPUT113), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n957), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT114), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n965), .B(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(G303), .A2(G8), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT55), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G40), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n472), .A2(new_n483), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(G1384), .B1(new_n836), .B2(new_n837), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n972), .B1(new_n973), .B2(KEYINPUT45), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT115), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(new_n973), .B2(KEYINPUT45), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n973), .A2(new_n975), .A3(KEYINPUT45), .ZN(new_n978));
  AOI21_X1  g553(.A(G1971), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n981));
  INV_X1    g556(.A(G1384), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n838), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n980), .A2(new_n972), .A3(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n984), .A2(G2090), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n970), .B(G8), .C1(new_n979), .C2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1976), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT52), .B1(G288), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n973), .A2(new_n972), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n576), .A2(G1976), .A3(new_n577), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n989), .A2(new_n990), .A3(G8), .A4(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(G8), .A3(new_n991), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT52), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n990), .A2(G8), .ZN(new_n996));
  INV_X1    g571(.A(G1981), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n530), .A2(G86), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n997), .B1(new_n587), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(G305), .B2(G1981), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT49), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n996), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n696), .A2(new_n997), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(KEYINPUT49), .A3(new_n1000), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n995), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n987), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1008));
  NOR2_X1   g583(.A1(G288), .A2(G1976), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n996), .B1(new_n1010), .B2(new_n1004), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n838), .A2(new_n982), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n948), .B1(new_n1013), .B2(new_n946), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n838), .A2(KEYINPUT45), .A3(new_n982), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT115), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1014), .A2(new_n978), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n972), .B1(new_n973), .B2(new_n981), .ZN(new_n1018));
  NOR3_X1   g593(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI22_X1  g595(.A1(new_n1017), .A2(new_n702), .B1(new_n1020), .B2(new_n797), .ZN(new_n1021));
  INV_X1    g596(.A(G8), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n969), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G2084), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n947), .A2(new_n972), .A3(new_n1015), .ZN(new_n1025));
  INV_X1    g600(.A(G1966), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1020), .A2(new_n1024), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1027), .A2(new_n1022), .A3(G286), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1023), .A2(new_n986), .A3(new_n1006), .A4(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT63), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1012), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1012), .B(KEYINPUT116), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT51), .ZN(new_n1038));
  NOR2_X1   g613(.A1(G168), .A2(new_n1022), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1038), .B1(new_n1039), .B2(KEYINPUT123), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1042), .B1(G2084), .B2(new_n984), .ZN(new_n1043));
  OAI211_X1 g618(.A(G8), .B(new_n1041), .C1(new_n1043), .C2(G286), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1039), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1045), .B(new_n1040), .C1(new_n1027), .C2(new_n1022), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1043), .A2(new_n1039), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1044), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT62), .ZN(new_n1049));
  OR2_X1    g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1023), .A2(new_n986), .A3(new_n1006), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1014), .A2(new_n790), .A3(new_n1016), .A4(new_n978), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n1054));
  INV_X1    g629(.A(G1961), .ZN(new_n1055));
  AOI22_X1  g630(.A1(new_n1053), .A2(new_n1054), .B1(new_n1055), .B2(new_n984), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT124), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n1025), .B2(G2078), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1014), .A2(KEYINPUT124), .A3(new_n790), .A4(new_n1015), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(KEYINPUT53), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G171), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1052), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1050), .A2(new_n1051), .A3(new_n1063), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n1065));
  NAND2_X1  g640(.A1(G299), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT119), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n1068));
  NAND3_X1  g643(.A1(G299), .A2(new_n1068), .A3(new_n1065), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1067), .B(new_n1069), .C1(new_n1070), .C2(G299), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT56), .B(G2072), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n977), .A2(new_n978), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT117), .B1(new_n984), .B2(new_n783), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n984), .A2(KEYINPUT117), .A3(new_n783), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1071), .B(new_n1073), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G1348), .ZN(new_n1078));
  INV_X1    g653(.A(new_n990), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n984), .A2(new_n1078), .B1(new_n1079), .B2(new_n952), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1080), .A2(new_n614), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n1081), .B(KEYINPUT120), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1073), .B1(new_n1075), .B2(new_n1074), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1071), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1077), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT61), .B1(new_n1085), .B2(new_n1076), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1078), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1079), .A2(new_n952), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT60), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT122), .B1(new_n1090), .B2(new_n614), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1080), .A2(KEYINPUT60), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT122), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1093), .B(new_n603), .C1(new_n1080), .C2(KEYINPUT60), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1091), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1092), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1087), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT58), .B(G1341), .Z(new_n1100));
  NAND3_X1  g675(.A1(new_n990), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1099), .B1(new_n990), .B2(new_n1100), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n977), .A2(new_n950), .A3(new_n978), .ZN(new_n1105));
  AOI211_X1 g680(.A(new_n1098), .B(new_n554), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1103), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1107), .B(new_n1101), .C1(new_n1017), .C2(G1996), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT59), .B1(new_n1108), .B2(new_n555), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1085), .A2(new_n1076), .A3(KEYINPUT61), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1086), .B1(new_n1097), .B2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n977), .A2(KEYINPUT53), .A3(new_n790), .A4(new_n978), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1056), .A2(G301), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT125), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT125), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1056), .A2(new_n1117), .A3(G301), .A4(new_n1114), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1116), .A2(new_n1118), .A3(new_n1062), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1056), .A2(new_n1114), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1120), .B1(new_n1122), .B2(G171), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(G171), .B2(new_n1061), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1048), .A2(new_n1052), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1121), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1064), .B1(new_n1113), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n967), .B1(new_n1037), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n954), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n689), .A2(new_n955), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1129), .A2(new_n1130), .B1(new_n952), .B2(new_n832), .ZN(new_n1131));
  INV_X1    g706(.A(new_n949), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT127), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n949), .A2(KEYINPUT46), .A3(new_n950), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT46), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1132), .B2(G1996), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n724), .A2(new_n953), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1135), .B(new_n1137), .C1(new_n1138), .C2(new_n1132), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT47), .ZN(new_n1140));
  XOR2_X1   g715(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1141));
  XNOR2_X1  g716(.A(new_n960), .B(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n957), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1133), .A2(new_n1134), .A3(new_n1140), .A4(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1143), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1140), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT127), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1128), .A2(new_n1148), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g724(.A(G319), .ZN(new_n1151));
  NOR4_X1   g725(.A1(G229), .A2(new_n1151), .A3(G401), .A4(G227), .ZN(new_n1152));
  OAI211_X1 g726(.A(new_n869), .B(new_n1152), .C1(new_n933), .C2(new_n940), .ZN(G225));
  INV_X1    g727(.A(G225), .ZN(G308));
endmodule


