//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n852, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT73), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n209), .A2(new_n210), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n207), .B(new_n208), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT74), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n207), .B1(new_n211), .B2(new_n212), .ZN(new_n215));
  INV_X1    g014(.A(new_n208), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n216), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(KEYINPUT74), .A3(new_n213), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G226gat), .ZN(new_n221));
  INV_X1    g020(.A(G233gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n227), .A2(KEYINPUT26), .ZN(new_n228));
  NAND2_X1  g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n227), .B1(new_n230), .B2(KEYINPUT26), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n225), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT66), .B(G190gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT27), .B(G183gat), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n233), .A2(new_n234), .B1(KEYINPUT67), .B2(KEYINPUT28), .ZN(new_n235));
  NOR2_X1   g034(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI211_X1 g036(.A(KEYINPUT67), .B(KEYINPUT28), .C1(new_n233), .C2(new_n234), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n232), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G183gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n233), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n225), .B1(new_n242), .B2(KEYINPUT24), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT24), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n224), .A2(KEYINPUT65), .A3(new_n244), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n241), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n226), .B1(KEYINPUT23), .B2(new_n229), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n226), .A2(KEYINPUT23), .ZN(new_n248));
  OR2_X1    g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT25), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  NOR3_X1   g049(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT25), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n225), .A2(KEYINPUT24), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n224), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT64), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n255), .B1(new_n252), .B2(new_n254), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n251), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n239), .A2(new_n250), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT29), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n223), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n259), .A2(new_n223), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n220), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n263), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n214), .B(new_n218), .ZN(new_n266));
  NOR3_X1   g065(.A1(new_n265), .A2(new_n261), .A3(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n206), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT30), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(KEYINPUT75), .A3(new_n269), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n259), .A2(new_n260), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n263), .B(new_n220), .C1(new_n271), .C2(new_n223), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n266), .B1(new_n265), .B2(new_n261), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n205), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT75), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT30), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n272), .A2(new_n273), .A3(new_n205), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n270), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G1gat), .B(G29gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT0), .ZN(new_n281));
  XNOR2_X1  g080(.A(G57gat), .B(G85gat), .ZN(new_n282));
  XOR2_X1   g081(.A(new_n281), .B(new_n282), .Z(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  XOR2_X1   g083(.A(KEYINPUT79), .B(G155gat), .Z(new_n285));
  INV_X1    g084(.A(G162gat), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT2), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G141gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G148gat), .ZN(new_n289));
  XOR2_X1   g088(.A(KEYINPUT78), .B(G148gat), .Z(new_n290));
  OAI21_X1  g089(.A(new_n289), .B1(new_n290), .B2(new_n288), .ZN(new_n291));
  XNOR2_X1  g090(.A(G155gat), .B(G162gat), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n287), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT76), .B1(G155gat), .B2(G162gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NOR3_X1   g095(.A1(KEYINPUT76), .A2(G155gat), .A3(G162gat), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT77), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT76), .ZN(new_n301));
  INV_X1    g100(.A(G155gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n302), .A3(new_n286), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n303), .A2(new_n295), .B1(G155gat), .B2(G162gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT77), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n294), .A2(KEYINPUT2), .ZN(new_n306));
  XOR2_X1   g105(.A(G141gat), .B(G148gat), .Z(new_n307));
  AOI22_X1  g106(.A1(new_n300), .A2(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT3), .B1(new_n293), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n306), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n298), .A2(new_n299), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n304), .A2(KEYINPUT77), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT3), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n287), .A2(new_n291), .A3(new_n292), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G120gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G113gat), .ZN(new_n318));
  INV_X1    g117(.A(G113gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G120gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT1), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G127gat), .B(G134gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n323), .A2(KEYINPUT68), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT68), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT1), .B1(new_n318), .B2(new_n320), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n327), .B1(new_n328), .B2(new_n324), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n325), .A2(KEYINPUT1), .ZN(new_n331));
  OR3_X1    g130(.A1(new_n319), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT69), .B1(new_n319), .B2(G120gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n318), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n330), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n309), .A2(new_n316), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n293), .A2(new_n308), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n326), .A2(new_n329), .B1(new_n331), .B2(new_n335), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(KEYINPUT4), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n313), .A2(new_n341), .A3(new_n315), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT4), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n338), .A2(new_n339), .A3(new_n342), .A4(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT5), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n337), .B1(new_n293), .B2(new_n308), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n343), .ZN(new_n350));
  INV_X1    g149(.A(new_n339), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n346), .A2(new_n352), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n284), .B(new_n348), .C1(new_n353), .C2(new_n347), .ZN(new_n354));
  INV_X1    g153(.A(new_n348), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n347), .B1(new_n346), .B2(new_n352), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n283), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT6), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n354), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n355), .A2(new_n356), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(KEYINPUT6), .A3(new_n284), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n279), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n259), .A2(new_n341), .ZN(new_n364));
  AND2_X1   g163(.A1(G227gat), .A2(G233gat), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n239), .A2(new_n337), .A3(new_n250), .A4(new_n258), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(G15gat), .B(G43gat), .Z(new_n368));
  XNOR2_X1  g167(.A(G71gat), .B(G99gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT33), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(KEYINPUT32), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT70), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n367), .A2(KEYINPUT70), .A3(KEYINPUT32), .A4(new_n371), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n365), .B1(new_n364), .B2(new_n366), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT34), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n377), .A2(new_n378), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n370), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n382), .B1(new_n367), .B2(KEYINPUT32), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT33), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n376), .A2(new_n381), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT72), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AND2_X1   g188(.A1(G228gat), .A2(G233gat), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT3), .B1(new_n266), .B2(new_n260), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n316), .A2(new_n260), .B1(new_n217), .B2(new_n219), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT80), .ZN(new_n393));
  OAI22_X1  g192(.A1(new_n391), .A2(new_n340), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n316), .A2(new_n260), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n220), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n396), .A2(KEYINPUT80), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n390), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n390), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n218), .A2(new_n213), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT3), .B1(new_n400), .B2(new_n260), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n396), .B(new_n399), .C1(new_n340), .C2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G78gat), .B(G106gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT31), .B(G50gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n403), .B(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(G22gat), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n398), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n406), .B1(new_n398), .B2(new_n402), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n376), .A2(new_n386), .ZN(new_n410));
  INV_X1    g209(.A(new_n381), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n376), .A2(new_n381), .A3(KEYINPUT72), .A4(new_n386), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n389), .A2(new_n409), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n202), .B1(new_n363), .B2(new_n414), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n409), .A2(new_n412), .A3(new_n387), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n416), .A2(KEYINPUT35), .A3(new_n362), .A4(new_n279), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n409), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n279), .A2(new_n419), .A3(new_n362), .ZN(new_n420));
  INV_X1    g219(.A(new_n362), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT37), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n272), .A2(new_n273), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n422), .B1(new_n272), .B2(new_n273), .ZN(new_n424));
  OAI211_X1 g223(.A(KEYINPUT38), .B(new_n205), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT37), .B1(new_n264), .B2(new_n267), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n272), .A2(new_n273), .A3(new_n422), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n206), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OR2_X1    g227(.A1(new_n274), .A2(KEYINPUT38), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n425), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n338), .A2(new_n345), .A3(new_n342), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n351), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n349), .A2(new_n339), .A3(new_n343), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT39), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT81), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT81), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(new_n436), .A3(KEYINPUT39), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n432), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT39), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n431), .A2(new_n439), .A3(new_n351), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n283), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT40), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n438), .A2(KEYINPUT40), .A3(new_n283), .A4(new_n440), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n443), .A2(new_n354), .A3(new_n444), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n421), .A2(new_n430), .B1(new_n445), .B2(new_n278), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n420), .B1(new_n446), .B2(new_n419), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT36), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n412), .A2(new_n413), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n374), .A2(new_n375), .B1(new_n385), .B2(new_n383), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT72), .B1(new_n450), .B2(new_n381), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n448), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n412), .A2(KEYINPUT36), .A3(new_n387), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT71), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n412), .A2(KEYINPUT71), .A3(KEYINPUT36), .A4(new_n387), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n452), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n418), .B1(new_n447), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(G113gat), .B(G141gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT11), .ZN(new_n460));
  INV_X1    g259(.A(G169gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n462), .B(G197gat), .ZN(new_n463));
  XOR2_X1   g262(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n464));
  XNOR2_X1  g263(.A(new_n463), .B(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(G22gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(G15gat), .ZN(new_n467));
  INV_X1    g266(.A(G15gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(G22gat), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT16), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n467), .B(new_n469), .C1(new_n470), .C2(G1gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(G15gat), .B(G22gat), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n471), .B1(G1gat), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G8gat), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT86), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n475), .B1(new_n472), .B2(G1gat), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  OAI221_X1 g276(.A(new_n471), .B1(new_n475), .B2(G8gat), .C1(G1gat), .C2(new_n472), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT83), .ZN(new_n481));
  NAND2_X1  g280(.A1(G29gat), .A2(G36gat), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NOR3_X1   g283(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n481), .B(new_n482), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(G50gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(G43gat), .ZN(new_n488));
  INV_X1    g287(.A(G43gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(G50gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n490), .A3(KEYINPUT15), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n488), .A2(new_n490), .A3(KEYINPUT15), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT14), .ZN(new_n494));
  INV_X1    g293(.A(G29gat), .ZN(new_n495));
  INV_X1    g294(.A(G36gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n483), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n493), .A2(new_n481), .A3(new_n498), .A4(new_n482), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n492), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n488), .ZN(new_n501));
  AND2_X1   g300(.A1(KEYINPUT84), .A2(G50gat), .ZN(new_n502));
  NOR2_X1   g301(.A1(KEYINPUT84), .A2(G50gat), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n489), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT85), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(KEYINPUT85), .B(new_n489), .C1(new_n502), .C2(new_n503), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT15), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n509), .B(new_n482), .C1(new_n484), .C2(new_n485), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n500), .A2(new_n512), .A3(KEYINPUT17), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT17), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n492), .A2(new_n499), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n510), .B1(new_n506), .B2(new_n507), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n480), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n500), .A2(new_n512), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(new_n479), .ZN(new_n520));
  NAND2_X1  g319(.A1(G229gat), .A2(G233gat), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n518), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT18), .B1(new_n523), .B2(KEYINPUT87), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT17), .B1(new_n500), .B2(new_n512), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n515), .A2(new_n516), .A3(new_n514), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n479), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n515), .A2(new_n516), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n480), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n527), .A2(new_n521), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT87), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT18), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n519), .A2(new_n479), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n529), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n521), .B(KEYINPUT13), .Z(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n465), .A2(new_n524), .A3(new_n533), .A4(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n464), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n463), .B(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n533), .A2(new_n537), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n532), .B1(new_n530), .B2(new_n531), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT88), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n524), .A2(new_n533), .A3(new_n537), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT88), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(new_n547), .A3(new_n541), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n539), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n458), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT97), .ZN(new_n551));
  XOR2_X1   g350(.A(G183gat), .B(G211gat), .Z(new_n552));
  XNOR2_X1  g351(.A(G127gat), .B(G155gat), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(KEYINPUT20), .Z(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT90), .ZN(new_n556));
  INV_X1    g355(.A(G64gat), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n557), .A2(G57gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT89), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n557), .A2(G57gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n561), .A2(KEYINPUT89), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n560), .B1(new_n562), .B2(new_n558), .ZN(new_n563));
  NAND2_X1  g362(.A1(G71gat), .A2(G78gat), .ZN(new_n564));
  OR2_X1    g363(.A1(G71gat), .A2(G78gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT9), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT9), .B1(new_n558), .B2(new_n561), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n569), .A2(new_n564), .A3(new_n565), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT21), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n556), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n571), .A2(new_n556), .A3(new_n572), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n574), .A2(G231gat), .A3(G233gat), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577));
  INV_X1    g376(.A(new_n575), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n577), .B1(new_n578), .B2(new_n573), .ZN(new_n579));
  XOR2_X1   g378(.A(KEYINPUT91), .B(KEYINPUT19), .Z(new_n580));
  NAND3_X1  g379(.A1(new_n576), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n580), .B1(new_n576), .B2(new_n579), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n555), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n583), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(new_n554), .A3(new_n581), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n568), .A2(new_n570), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n480), .B1(KEYINPUT21), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n584), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n589), .B1(new_n584), .B2(new_n586), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n552), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n584), .A2(new_n586), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(new_n588), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n584), .A2(new_n586), .A3(new_n589), .ZN(new_n595));
  INV_X1    g394(.A(new_n552), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(G99gat), .A2(G106gat), .ZN(new_n599));
  INV_X1    g398(.A(G85gat), .ZN(new_n600));
  INV_X1    g399(.A(G92gat), .ZN(new_n601));
  AOI22_X1  g400(.A1(KEYINPUT8), .A2(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT7), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n603), .B1(new_n600), .B2(new_n601), .ZN(new_n604));
  NAND3_X1  g403(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n602), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G99gat), .B(G106gat), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n608), .B1(new_n525), .B2(new_n526), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT41), .ZN(new_n610));
  NAND2_X1  g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n611), .B(KEYINPUT92), .Z(new_n612));
  OAI22_X1  g411(.A1(new_n519), .A2(new_n608), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n613), .A2(KEYINPUT94), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n613), .A2(KEYINPUT94), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n609), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G190gat), .B(G218gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n617), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n609), .B(new_n619), .C1(new_n614), .C2(new_n615), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n612), .A2(new_n610), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT93), .ZN(new_n623));
  XNOR2_X1  g422(.A(G134gat), .B(G162gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n625), .B1(new_n620), .B2(KEYINPUT95), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n618), .B(new_n620), .C1(KEYINPUT95), .C2(new_n625), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n598), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n608), .A2(new_n571), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n606), .A2(new_n607), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n606), .A2(new_n607), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n635), .A2(new_n568), .A3(new_n570), .A4(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(G230gat), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n639), .A2(new_n222), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n634), .A2(new_n643), .A3(new_n637), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n587), .A2(KEYINPUT10), .A3(new_n635), .A4(new_n636), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT96), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n633), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n633), .ZN(new_n650));
  OAI211_X1 g449(.A(KEYINPUT96), .B(new_n650), .C1(new_n642), .C2(new_n646), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n630), .A2(new_n653), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n550), .A2(new_n551), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n551), .B1(new_n550), .B2(new_n654), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n421), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT98), .B(G1gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1324gat));
  XNOR2_X1  g460(.A(KEYINPUT16), .B(G8gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT99), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n278), .B(new_n663), .C1(new_n655), .C2(new_n656), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(KEYINPUT42), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT42), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n278), .B1(new_n655), .B2(new_n656), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n666), .B1(new_n667), .B2(G8gat), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n665), .B1(new_n664), .B2(new_n668), .ZN(G1325gat));
  OAI21_X1  g468(.A(G15gat), .B1(new_n657), .B2(new_n457), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n449), .A2(new_n451), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n468), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n657), .B2(new_n672), .ZN(G1326gat));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n409), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT43), .B(G22gat), .Z(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1327gat));
  NOR3_X1   g475(.A1(new_n598), .A2(new_n629), .A3(new_n653), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT100), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n550), .A2(new_n495), .A3(new_n421), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT101), .B(KEYINPUT45), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n598), .A2(KEYINPUT102), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n592), .A2(new_n597), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n549), .A2(new_n653), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n685), .A2(KEYINPUT103), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT103), .B1(new_n685), .B2(new_n686), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n629), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n691));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n430), .A2(new_n361), .A3(new_n359), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n278), .A2(new_n354), .A3(new_n444), .A4(new_n443), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n419), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n420), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n457), .B(new_n692), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n415), .A2(new_n417), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n692), .B1(new_n447), .B2(new_n457), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n690), .B(new_n691), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT44), .B1(new_n458), .B2(new_n629), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n689), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n495), .B1(new_n703), .B2(new_n421), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT106), .ZN(new_n705));
  OR3_X1    g504(.A1(new_n681), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n705), .B1(new_n681), .B2(new_n704), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(G1328gat));
  AND2_X1   g507(.A1(new_n550), .A2(new_n678), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n709), .A2(new_n496), .A3(new_n278), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT46), .Z(new_n711));
  INV_X1    g510(.A(new_n703), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n279), .ZN(new_n713));
  OAI21_X1  g512(.A(G36gat), .B1(new_n713), .B2(KEYINPUT107), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n713), .A2(KEYINPUT107), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n711), .B1(new_n714), .B2(new_n715), .ZN(G1329gat));
  AND2_X1   g515(.A1(new_n709), .A2(new_n671), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(G43gat), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n457), .A2(new_n489), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n712), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT47), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722));
  OAI221_X1 g521(.A(new_n722), .B1(new_n712), .B2(new_n719), .C1(new_n717), .C2(G43gat), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(G1330gat));
  NOR2_X1   g523(.A1(new_n502), .A2(new_n503), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n709), .A2(new_n419), .A3(new_n725), .ZN(new_n726));
  AOI211_X1 g525(.A(new_n409), .B(new_n689), .C1(new_n701), .C2(new_n702), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(new_n725), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT108), .B1(new_n727), .B2(new_n725), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n728), .A2(new_n729), .A3(KEYINPUT48), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n731));
  OAI221_X1 g530(.A(new_n726), .B1(KEYINPUT108), .B2(new_n731), .C1(new_n727), .C2(new_n725), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n730), .A2(new_n732), .ZN(G1331gat));
  OR2_X1    g532(.A1(new_n699), .A2(new_n700), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n546), .A2(new_n547), .A3(new_n541), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n547), .B1(new_n546), .B2(new_n541), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n538), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n630), .A2(new_n737), .A3(new_n652), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n421), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g541(.A(new_n279), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT109), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n744), .B(new_n746), .ZN(G1333gat));
  OAI21_X1  g546(.A(G71gat), .B1(new_n739), .B2(new_n457), .ZN(new_n748));
  INV_X1    g547(.A(G71gat), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n671), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n748), .B1(new_n739), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1334gat));
  NAND2_X1  g552(.A1(new_n740), .A2(new_n419), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g554(.A1(new_n598), .A2(new_n737), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n690), .B(new_n756), .C1(new_n699), .C2(new_n700), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n759), .A2(new_n600), .A3(new_n421), .A4(new_n653), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n756), .A2(new_n653), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT110), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n762), .B1(new_n701), .B2(new_n702), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(G85gat), .B1(new_n764), .B2(new_n362), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n760), .A2(new_n765), .ZN(G1336gat));
  AND3_X1   g565(.A1(new_n757), .A2(KEYINPUT111), .A3(KEYINPUT51), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT51), .B1(new_n757), .B2(KEYINPUT111), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n279), .A2(G92gat), .A3(new_n652), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n767), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n601), .B1(new_n763), .B2(new_n278), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT52), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(KEYINPUT112), .B1(new_n764), .B2(new_n279), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n763), .A2(new_n775), .A3(new_n278), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n601), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n759), .A2(new_n769), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n773), .B1(new_n777), .B2(new_n780), .ZN(G1337gat));
  NOR2_X1   g580(.A1(new_n652), .A2(G99gat), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n759), .A2(new_n671), .A3(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(G99gat), .B1(new_n764), .B2(new_n457), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1338gat));
  NOR3_X1   g584(.A1(new_n409), .A2(G106gat), .A3(new_n652), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT53), .B1(new_n759), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(KEYINPUT113), .B(G106gat), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n789), .B1(new_n763), .B2(new_n419), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n786), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n767), .A2(new_n768), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT53), .B1(new_n794), .B2(new_n790), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n792), .A2(new_n795), .ZN(G1339gat));
  NAND4_X1  g595(.A1(new_n598), .A2(new_n549), .A3(new_n629), .A4(new_n652), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n646), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n644), .A2(new_n645), .A3(new_n640), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI211_X1 g600(.A(KEYINPUT54), .B(new_n640), .C1(new_n644), .C2(new_n645), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n802), .A2(new_n803), .A3(new_n650), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n644), .A2(new_n645), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n805), .A2(new_n798), .A3(new_n641), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT114), .B1(new_n806), .B2(new_n633), .ZN(new_n807));
  OAI211_X1 g606(.A(KEYINPUT55), .B(new_n801), .C1(new_n804), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n647), .A2(new_n650), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n803), .B1(new_n802), .B2(new_n650), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n806), .A2(KEYINPUT114), .A3(new_n633), .ZN(new_n812));
  AOI22_X1  g611(.A1(new_n811), .A2(new_n812), .B1(new_n800), .B2(new_n799), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(KEYINPUT55), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n521), .B1(new_n527), .B2(new_n529), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n535), .A2(new_n536), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n463), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n538), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n690), .A2(new_n815), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n819), .A2(new_n652), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n822), .B1(new_n737), .B2(new_n815), .ZN(new_n823));
  OAI211_X1 g622(.A(KEYINPUT115), .B(new_n821), .C1(new_n823), .C2(new_n690), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n685), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n820), .A2(new_n653), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n801), .B1(new_n804), .B2(new_n807), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n829), .A2(new_n809), .A3(new_n808), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n826), .B1(new_n549), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n629), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT115), .B1(new_n832), .B2(new_n821), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n797), .B1(new_n825), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n362), .A2(new_n278), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n416), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n549), .A2(G113gat), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT118), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  OR3_X1    g640(.A1(new_n836), .A2(KEYINPUT116), .A3(new_n414), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT116), .B1(new_n836), .B2(new_n414), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n737), .A3(new_n843), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n844), .A2(KEYINPUT117), .A3(G113gat), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT117), .B1(new_n844), .B2(G113gat), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n841), .B1(new_n845), .B2(new_n846), .ZN(G1340gat));
  AOI21_X1  g646(.A(G120gat), .B1(new_n838), .B2(new_n653), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n842), .A2(new_n843), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n652), .A2(new_n317), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(G1341gat));
  INV_X1    g650(.A(G127gat), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n838), .A2(new_n852), .A3(new_n598), .ZN(new_n853));
  INV_X1    g652(.A(new_n685), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n853), .B1(new_n855), .B2(new_n852), .ZN(G1342gat));
  NAND2_X1  g655(.A1(new_n849), .A2(new_n690), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(G134gat), .ZN(new_n858));
  NOR4_X1   g657(.A1(new_n836), .A2(G134gat), .A3(new_n837), .A4(new_n629), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT56), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(G1343gat));
  NAND2_X1  g660(.A1(new_n457), .A2(new_n419), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n737), .A2(new_n288), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n836), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n457), .A2(new_n835), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  XNOR2_X1  g665(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n868), .B1(new_n834), .B2(new_n419), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n419), .A2(KEYINPUT57), .ZN(new_n870));
  INV_X1    g669(.A(new_n598), .ZN(new_n871));
  XOR2_X1   g670(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n872));
  NOR2_X1   g671(.A1(new_n813), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n874), .A2(KEYINPUT121), .A3(new_n809), .A4(new_n808), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n876), .B1(new_n810), .B2(new_n873), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n877), .A3(new_n737), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n690), .B1(new_n878), .B2(new_n826), .ZN(new_n879));
  INV_X1    g678(.A(new_n821), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n871), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n870), .B1(new_n881), .B2(new_n797), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n737), .B(new_n866), .C1(new_n869), .C2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n864), .B1(new_n883), .B2(G141gat), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT58), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n883), .A2(G141gat), .ZN(new_n887));
  INV_X1    g686(.A(new_n864), .ZN(new_n888));
  AND4_X1   g687(.A1(KEYINPUT122), .A2(new_n887), .A3(new_n885), .A4(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT122), .B1(new_n884), .B2(new_n885), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(G1344gat));
  NOR2_X1   g690(.A1(new_n836), .A2(new_n862), .ZN(new_n892));
  INV_X1    g691(.A(new_n290), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n893), .A3(new_n653), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n797), .B(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n881), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n419), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n834), .A2(new_n419), .A3(new_n868), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n653), .A3(new_n866), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n895), .B1(new_n904), .B2(G148gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n866), .B1(new_n869), .B2(new_n882), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  AOI211_X1 g706(.A(KEYINPUT59), .B(new_n893), .C1(new_n907), .C2(new_n653), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n894), .B1(new_n905), .B2(new_n908), .ZN(G1345gat));
  INV_X1    g708(.A(new_n285), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(new_n906), .B2(new_n685), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n892), .A2(new_n285), .A3(new_n598), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1346gat));
  OAI21_X1  g712(.A(G162gat), .B1(new_n906), .B2(new_n629), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n892), .A2(new_n286), .A3(new_n690), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1347gat));
  NOR2_X1   g715(.A1(new_n421), .A2(new_n279), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n821), .B1(new_n823), .B2(new_n690), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT115), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n685), .A3(new_n824), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n918), .B1(new_n922), .B2(new_n797), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n924), .A2(new_n837), .ZN(new_n925));
  AOI21_X1  g724(.A(G169gat), .B1(new_n925), .B2(new_n737), .ZN(new_n926));
  INV_X1    g725(.A(new_n414), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n834), .A2(new_n927), .A3(new_n917), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT124), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n923), .A2(new_n930), .A3(new_n927), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n549), .A2(new_n461), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n926), .B1(new_n932), .B2(new_n933), .ZN(G1348gat));
  AOI21_X1  g733(.A(G176gat), .B1(new_n925), .B2(new_n653), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n932), .A2(G176gat), .A3(new_n653), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n932), .A2(KEYINPUT125), .A3(G176gat), .A4(new_n653), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(G1349gat));
  AND2_X1   g739(.A1(new_n598), .A2(new_n234), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n834), .A2(new_n416), .A3(new_n917), .A4(new_n941), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n942), .A2(KEYINPUT126), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n942), .A2(KEYINPUT126), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT60), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n945), .A2(KEYINPUT127), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n929), .A2(new_n931), .A3(new_n854), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(G183gat), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n945), .A2(KEYINPUT127), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(new_n947), .B2(new_n949), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(G1350gat));
  NAND3_X1  g752(.A1(new_n925), .A2(new_n233), .A3(new_n690), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n929), .A2(new_n931), .A3(new_n690), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n955), .A2(new_n956), .A3(G190gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n956), .B1(new_n955), .B2(G190gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n954), .B1(new_n957), .B2(new_n958), .ZN(G1351gat));
  NOR2_X1   g758(.A1(new_n924), .A2(new_n862), .ZN(new_n960));
  AOI21_X1  g759(.A(G197gat), .B1(new_n960), .B2(new_n737), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n457), .A2(new_n917), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n962), .B1(new_n901), .B2(new_n902), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n737), .A2(G197gat), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1352gat));
  NOR4_X1   g764(.A1(new_n924), .A2(G204gat), .A3(new_n652), .A4(new_n862), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT62), .ZN(new_n967));
  AOI211_X1 g766(.A(new_n652), .B(new_n962), .C1(new_n901), .C2(new_n902), .ZN(new_n968));
  INV_X1    g767(.A(G204gat), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(G1353gat));
  INV_X1    g769(.A(G211gat), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n960), .A2(new_n971), .A3(new_n598), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n963), .A2(new_n598), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT63), .B1(new_n973), .B2(G211gat), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT63), .ZN(new_n975));
  AOI211_X1 g774(.A(new_n975), .B(new_n971), .C1(new_n963), .C2(new_n598), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n972), .B1(new_n974), .B2(new_n976), .ZN(G1354gat));
  INV_X1    g776(.A(G218gat), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n960), .A2(new_n978), .A3(new_n690), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n963), .A2(new_n690), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n979), .B1(new_n980), .B2(new_n978), .ZN(G1355gat));
endmodule


