//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1187, new_n1188, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  AOI211_X1 g0011(.A(new_n206), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  OAI22_X1  g0017(.A1(new_n212), .A2(KEYINPUT0), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n219), .B1(new_n202), .B2(new_n220), .C1(new_n221), .C2(new_n206), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  INV_X1    g0025(.A(G68), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n207), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n218), .B(new_n230), .C1(KEYINPUT0), .C2(new_n212), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT64), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  INV_X1    g0041(.A(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT65), .B(G107), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n202), .A2(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n226), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n245), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(G222), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G77), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(G1698), .ZN(new_n261));
  INV_X1    g0061(.A(G223), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n259), .B1(new_n260), .B2(new_n257), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n267));
  INV_X1    g0067(.A(G274), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n264), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n267), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n269), .B1(new_n272), .B2(G226), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n265), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G200), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT68), .ZN(new_n276));
  INV_X1    g0076(.A(G190), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n275), .B(new_n276), .C1(new_n277), .C2(new_n274), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n213), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n280), .B1(new_n266), .B2(G20), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G50), .ZN(new_n282));
  INV_X1    g0082(.A(G13), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n283), .A2(new_n214), .A3(G1), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n282), .B1(G50), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n280), .ZN(new_n287));
  XOR2_X1   g0087(.A(KEYINPUT8), .B(G58), .Z(new_n288));
  NAND2_X1  g0088(.A1(new_n214), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n288), .A2(new_n290), .B1(G20), .B2(new_n203), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n214), .A2(new_n252), .A3(KEYINPUT66), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT66), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(G20), .B2(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G150), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n287), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n286), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(KEYINPUT67), .A2(KEYINPUT9), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT67), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT9), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n299), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n298), .A2(new_n301), .A3(new_n302), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT10), .B1(new_n278), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n274), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT68), .B1(new_n308), .B2(G190), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT10), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n304), .A2(new_n305), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .A4(new_n275), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n299), .B1(new_n308), .B2(G169), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n274), .A2(G179), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n295), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(new_n202), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n289), .A2(new_n260), .B1(new_n214), .B2(G68), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n280), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT11), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n323), .ZN(new_n325));
  OR3_X1    g0125(.A1(new_n285), .A2(KEYINPUT12), .A3(G68), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT12), .B1(new_n285), .B2(G68), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n326), .A2(new_n327), .B1(G68), .B2(new_n281), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n324), .A2(new_n325), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n257), .A2(G232), .A3(G1698), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n257), .A2(G226), .A3(new_n258), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G97), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n264), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n269), .B1(new_n272), .B2(G238), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT13), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT13), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n334), .A2(new_n338), .A3(new_n335), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(G179), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G169), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n341), .B1(new_n337), .B2(new_n339), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT14), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n334), .A2(new_n338), .A3(new_n335), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n338), .B1(new_n334), .B2(new_n335), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n343), .B(G169), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n329), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n345), .A2(new_n346), .ZN(new_n350));
  INV_X1    g0150(.A(G200), .ZN(new_n351));
  OAI21_X1  g0151(.A(KEYINPUT69), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n329), .B1(new_n350), .B2(G190), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT69), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n354), .B(G200), .C1(new_n345), .C2(new_n346), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G107), .ZN(new_n358));
  OAI22_X1  g0158(.A1(new_n261), .A2(new_n227), .B1(new_n358), .B2(new_n257), .ZN(new_n359));
  NOR3_X1   g0159(.A1(new_n256), .A2(new_n225), .A3(G1698), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n264), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n269), .B1(new_n272), .B2(G244), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  XOR2_X1   g0163(.A(KEYINPUT15), .B(G87), .Z(new_n364));
  AOI22_X1  g0164(.A1(new_n364), .A2(new_n290), .B1(G20), .B2(G77), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n288), .A2(new_n295), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n287), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n281), .A2(G77), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(G77), .B2(new_n285), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n363), .A2(G169), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n361), .A2(new_n362), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n371), .A2(G179), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n363), .A2(new_n351), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n369), .A2(new_n367), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n371), .B2(new_n277), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n373), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n318), .A2(new_n357), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT17), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT16), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n256), .A2(new_n214), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT7), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n256), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n226), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n224), .A2(new_n226), .ZN(new_n386));
  OR2_X1    g0186(.A1(new_n386), .A2(new_n201), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n387), .A2(G20), .B1(G159), .B2(new_n295), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n380), .B1(new_n385), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT70), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n252), .B2(KEYINPUT3), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n253), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n252), .A3(KEYINPUT3), .ZN(new_n394));
  AOI21_X1  g0194(.A(G20), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(G68), .B1(new_n395), .B2(new_n382), .ZN(new_n396));
  NOR3_X1   g0196(.A1(new_n254), .A2(KEYINPUT70), .A3(G33), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(new_n253), .B2(new_n392), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n398), .A2(KEYINPUT7), .A3(G20), .ZN(new_n399));
  OAI211_X1 g0199(.A(KEYINPUT16), .B(new_n388), .C1(new_n396), .C2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n390), .A2(new_n400), .A3(new_n280), .ZN(new_n401));
  INV_X1    g0201(.A(new_n288), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n285), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(new_n281), .B2(new_n402), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n398), .A2(KEYINPUT71), .A3(G223), .A4(new_n258), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n220), .A2(new_n258), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT70), .B1(new_n254), .B2(G33), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n254), .A2(G33), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n394), .B(new_n406), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G87), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT71), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n258), .B(new_n394), .C1(new_n407), .C2(new_n408), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n412), .B1(new_n413), .B2(new_n262), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n405), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n264), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n271), .A2(new_n225), .B1(new_n268), .B2(new_n267), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(G200), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  AOI211_X1 g0219(.A(G190), .B(new_n417), .C1(new_n415), .C2(new_n264), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n401), .B(new_n404), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT73), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n379), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n401), .A2(new_n404), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n417), .B1(new_n415), .B2(new_n264), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n277), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(G200), .B2(new_n426), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n425), .A2(new_n428), .A3(KEYINPUT73), .A4(KEYINPUT17), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT74), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n423), .A2(new_n429), .A3(KEYINPUT74), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n426), .A2(G179), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n341), .B2(new_n426), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT18), .B1(new_n435), .B2(new_n424), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(KEYINPUT18), .A3(new_n424), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(KEYINPUT72), .A3(new_n438), .ZN(new_n439));
  AOI211_X1 g0239(.A(KEYINPUT72), .B(KEYINPUT18), .C1(new_n435), .C2(new_n424), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  AND4_X1   g0241(.A1(new_n432), .A2(new_n433), .A3(new_n439), .A4(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n378), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n444));
  NOR2_X1   g0244(.A1(G97), .A2(G107), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n214), .A2(new_n444), .B1(new_n445), .B2(new_n221), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT19), .ZN(new_n447));
  INV_X1    g0247(.A(G97), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n447), .B1(new_n289), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT77), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(KEYINPUT77), .B(new_n447), .C1(new_n289), .C2(new_n448), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n446), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n398), .A2(KEYINPUT76), .A3(new_n214), .A4(G68), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT76), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n214), .B(new_n394), .C1(new_n407), .C2(new_n408), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n456), .B2(new_n226), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n453), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n280), .ZN(new_n459));
  INV_X1    g0259(.A(new_n364), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n284), .ZN(new_n461));
  AOI211_X1 g0261(.A(new_n280), .B(new_n284), .C1(new_n266), .C2(G33), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n364), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n459), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n393), .A2(G244), .A3(G1698), .A4(new_n394), .ZN(new_n465));
  XNOR2_X1  g0265(.A(KEYINPUT75), .B(G116), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G33), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n413), .A2(new_n227), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n264), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G179), .ZN(new_n471));
  INV_X1    g0271(.A(G45), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(G1), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G274), .ZN(new_n474));
  OAI21_X1  g0274(.A(G250), .B1(new_n472), .B2(G1), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n474), .B1(new_n264), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n470), .A2(new_n471), .A3(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n465), .B(new_n467), .C1(new_n227), .C2(new_n413), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n476), .B1(new_n479), .B2(new_n264), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n478), .B1(G169), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n470), .A2(G190), .A3(new_n477), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n351), .B2(new_n480), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n462), .A2(G87), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n459), .A2(new_n461), .A3(new_n484), .ZN(new_n485));
  OAI22_X1  g0285(.A1(new_n464), .A2(new_n481), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT78), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n458), .A2(new_n280), .B1(new_n284), .B2(new_n460), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n463), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n489), .B(new_n478), .C1(G169), .C2(new_n480), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT78), .ZN(new_n491));
  INV_X1    g0291(.A(new_n480), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G200), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n493), .A2(new_n488), .A3(new_n484), .A4(new_n482), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n490), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n358), .B1(new_n383), .B2(new_n384), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT6), .ZN(new_n497));
  NOR3_X1   g0297(.A1(new_n497), .A2(new_n448), .A3(G107), .ZN(new_n498));
  XNOR2_X1  g0298(.A(G97), .B(G107), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n498), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OAI22_X1  g0300(.A1(new_n500), .A2(new_n214), .B1(new_n260), .B2(new_n319), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n280), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n284), .A2(new_n448), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n462), .A2(G97), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT4), .ZN(new_n506));
  OAI211_X1 g0306(.A(G244), .B(new_n394), .C1(new_n407), .C2(new_n408), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n506), .B1(new_n507), .B2(G1698), .ZN(new_n508));
  AND2_X1   g0308(.A1(KEYINPUT4), .A2(G244), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n253), .A2(new_n255), .A3(new_n509), .A4(new_n258), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n253), .A2(new_n255), .A3(G250), .A4(G1698), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G283), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n270), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g0314(.A1(KEYINPUT5), .A2(G41), .ZN(new_n515));
  NOR2_X1   g0315(.A1(KEYINPUT5), .A2(G41), .ZN(new_n516));
  OR2_X1    g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n264), .B1(new_n517), .B2(new_n473), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G257), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(G274), .A3(new_n473), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n514), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G190), .ZN(new_n523));
  OAI21_X1  g0323(.A(G200), .B1(new_n514), .B2(new_n521), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n505), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n520), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(new_n518), .B2(G257), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n508), .A2(new_n513), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n527), .B1(new_n528), .B2(new_n270), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n341), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n522), .A2(new_n471), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n525), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n487), .A2(new_n495), .A3(new_n534), .A4(KEYINPUT79), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n487), .A2(new_n495), .A3(new_n534), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT79), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n466), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n462), .A2(G116), .B1(new_n284), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n512), .B(new_n214), .C1(G33), .C2(new_n448), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n280), .B(new_n541), .C1(new_n466), .C2(new_n214), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT20), .ZN(new_n543));
  XNOR2_X1  g0343(.A(new_n542), .B(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n210), .A2(new_n258), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n211), .A2(G1698), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n393), .A2(new_n394), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  XNOR2_X1  g0348(.A(KEYINPUT80), .B(G303), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n256), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n264), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n473), .B1(new_n515), .B2(new_n516), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n270), .A2(new_n553), .A3(G270), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n554), .A2(new_n520), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n545), .A2(G169), .A3(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(KEYINPUT81), .A2(KEYINPUT21), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n558), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n545), .A2(G169), .A3(new_n560), .A4(new_n556), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n270), .B1(new_n548), .B2(new_n550), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n554), .A2(new_n520), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n562), .A2(new_n563), .A3(new_n471), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n545), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n556), .A2(G200), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n552), .A2(new_n555), .A3(G190), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n566), .A2(new_n544), .A3(new_n540), .A4(new_n567), .ZN(new_n568));
  AND4_X1   g0368(.A1(new_n559), .A2(new_n561), .A3(new_n565), .A4(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n394), .B1(new_n407), .B2(new_n408), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n210), .A2(G1698), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(G250), .B2(G1698), .ZN(new_n572));
  INV_X1    g0372(.A(G294), .ZN(new_n573));
  OAI22_X1  g0373(.A1(new_n570), .A2(new_n572), .B1(new_n252), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n264), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n518), .A2(G264), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(new_n520), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n351), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT83), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n577), .A2(KEYINPUT83), .A3(new_n351), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT82), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n575), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n574), .A2(KEYINPUT82), .A3(new_n264), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n583), .A2(new_n520), .A3(new_n584), .A4(new_n576), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n580), .B(new_n581), .C1(G190), .C2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n462), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n284), .A2(KEYINPUT25), .A3(new_n358), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT25), .B1(new_n284), .B2(new_n358), .ZN(new_n589));
  OAI22_X1  g0389(.A1(new_n587), .A2(new_n358), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n398), .A2(KEYINPUT22), .A3(new_n214), .A4(G87), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT22), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n214), .A2(G87), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(new_n256), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n214), .A2(G107), .ZN(new_n595));
  XNOR2_X1  g0395(.A(new_n595), .B(KEYINPUT23), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n466), .A2(new_n214), .A3(G33), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n591), .A2(new_n594), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT24), .ZN(new_n599));
  OR2_X1    g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n287), .B1(new_n598), .B2(new_n599), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n590), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n586), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n602), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n585), .A2(G169), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n575), .A2(new_n576), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(G179), .A3(new_n520), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n569), .A2(new_n603), .A3(new_n609), .ZN(new_n610));
  AND4_X1   g0410(.A1(new_n443), .A2(new_n535), .A3(new_n538), .A4(new_n610), .ZN(G372));
  NAND3_X1  g0411(.A1(new_n559), .A2(new_n561), .A3(new_n565), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n613), .A2(new_n609), .B1(new_n602), .B2(new_n586), .ZN(new_n614));
  INV_X1    g0414(.A(new_n486), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n614), .A2(KEYINPUT84), .A3(new_n615), .A4(new_n534), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT84), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n602), .B1(new_n605), .B2(new_n607), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n603), .B1(new_n618), .B2(new_n612), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n534), .A2(new_n615), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n533), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT26), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n616), .A2(new_n490), .A3(new_n621), .A4(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n487), .A2(new_n495), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n625), .B1(new_n628), .B2(new_n622), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n630), .A2(new_n443), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n435), .A2(KEYINPUT18), .A3(new_n424), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n632), .A2(new_n436), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n370), .A2(new_n372), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n356), .A2(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n635), .A2(KEYINPUT85), .A3(new_n349), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT85), .B1(new_n635), .B2(new_n349), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n423), .A2(KEYINPUT74), .A3(new_n429), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT74), .B1(new_n423), .B2(new_n429), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n633), .B1(new_n638), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n313), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n317), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n631), .A2(new_n644), .ZN(G369));
  AND2_X1   g0445(.A1(new_n603), .A2(new_n609), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n283), .A2(G20), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n266), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(G213), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(G343), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n604), .A2(new_n653), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n646), .A2(new_n654), .B1(new_n618), .B2(new_n653), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n613), .B2(new_n653), .ZN(new_n656));
  INV_X1    g0456(.A(new_n653), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n657), .B1(new_n544), .B2(new_n540), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n612), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n569), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n658), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n661), .A2(G330), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n646), .A2(new_n612), .A3(new_n657), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n618), .A2(new_n657), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n663), .A2(new_n666), .ZN(G399));
  NOR2_X1   g0467(.A1(new_n209), .A2(G41), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n445), .A2(new_n221), .A3(new_n242), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n669), .A2(G1), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n217), .B2(new_n669), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT28), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT29), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n675), .B(new_n657), .C1(new_n627), .C2(new_n629), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n522), .A2(new_n564), .A3(new_n606), .A4(new_n480), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT30), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n552), .A2(new_n555), .A3(G179), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n575), .A2(new_n576), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n682), .A2(KEYINPUT30), .A3(new_n480), .A4(new_n522), .ZN(new_n683));
  AOI21_X1  g0483(.A(G179), .B1(new_n552), .B2(new_n555), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n492), .A2(new_n529), .A3(new_n577), .A4(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n679), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n686), .A2(KEYINPUT31), .A3(new_n653), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT86), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT31), .B1(new_n686), .B2(new_n653), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n538), .A2(new_n610), .A3(new_n535), .A4(new_n657), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n623), .A2(KEYINPUT26), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n695), .B(new_n490), .C1(new_n620), .C2(new_n619), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n628), .A2(new_n625), .A3(new_n622), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n657), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(KEYINPUT29), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n676), .A2(new_n694), .A3(new_n699), .ZN(new_n700));
  XOR2_X1   g0500(.A(new_n700), .B(KEYINPUT87), .Z(new_n701));
  OAI21_X1  g0501(.A(new_n674), .B1(new_n701), .B2(G1), .ZN(G364));
  AOI21_X1  g0502(.A(new_n266), .B1(new_n647), .B2(G45), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n668), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n662), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(G330), .B2(new_n661), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n257), .A2(new_n208), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(KEYINPUT88), .B2(G355), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(KEYINPUT88), .B2(G355), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(G116), .B2(new_n208), .ZN(new_n711));
  MUX2_X1   g0511(.A(new_n217), .B(new_n250), .S(G45), .Z(new_n712));
  NAND2_X1  g0512(.A1(new_n570), .A2(new_n208), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n713), .B(KEYINPUT89), .Z(new_n714));
  AOI21_X1  g0514(.A(new_n711), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(G13), .A2(G33), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n214), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT90), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n213), .B1(G20), .B2(new_n341), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n705), .B1(new_n715), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n471), .A2(new_n351), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT91), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n214), .A2(G190), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G159), .ZN(new_n729));
  XOR2_X1   g0529(.A(new_n729), .B(KEYINPUT32), .Z(new_n730));
  OAI21_X1  g0530(.A(G20), .B1(new_n725), .B2(new_n277), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G97), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n471), .A2(new_n351), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n726), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n214), .A2(new_n277), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n351), .A2(G179), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI22_X1  g0539(.A1(G68), .A2(new_n735), .B1(new_n739), .B2(G87), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n736), .A2(new_n733), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n740), .B1(new_n202), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n471), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n726), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n257), .B1(new_n744), .B2(new_n260), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n736), .A2(new_n743), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n726), .A2(new_n737), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n746), .A2(new_n224), .B1(new_n747), .B2(new_n358), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n742), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n730), .A2(new_n732), .A3(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n741), .ZN(new_n751));
  INV_X1    g0551(.A(new_n744), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n751), .A2(G326), .B1(new_n752), .B2(G311), .ZN(new_n753));
  INV_X1    g0553(.A(new_n731), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n753), .B1(new_n754), .B2(new_n573), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT92), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n728), .A2(G329), .ZN(new_n757));
  XNOR2_X1  g0557(.A(KEYINPUT93), .B(KEYINPUT33), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n734), .B1(new_n758), .B2(G317), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(G317), .B2(new_n758), .ZN(new_n760));
  INV_X1    g0560(.A(new_n746), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n257), .B1(new_n761), .B2(G322), .ZN(new_n762));
  INV_X1    g0562(.A(new_n747), .ZN(new_n763));
  AOI22_X1  g0563(.A1(G303), .A2(new_n739), .B1(new_n763), .B2(G283), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n757), .A2(new_n760), .A3(new_n762), .A4(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n750), .B1(new_n756), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n723), .B1(new_n766), .B2(new_n720), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(new_n661), .B2(new_n718), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n707), .A2(new_n768), .ZN(G396));
  INV_X1    g0569(.A(new_n720), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n539), .A2(new_n744), .B1(new_n738), .B2(new_n358), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n257), .B(new_n771), .C1(G283), .C2(new_n735), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n728), .A2(G311), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n746), .A2(new_n573), .B1(new_n747), .B2(new_n221), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(G303), .B2(new_n751), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n772), .A2(new_n732), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G143), .A2(new_n761), .B1(new_n735), .B2(G150), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n751), .A2(G137), .B1(new_n752), .B2(G159), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(KEYINPUT34), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n738), .A2(new_n202), .B1(new_n747), .B2(new_n226), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n570), .B(new_n781), .C1(new_n728), .C2(G132), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n779), .A2(KEYINPUT34), .B1(new_n754), .B2(new_n224), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n776), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n770), .B1(new_n785), .B2(KEYINPUT95), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(KEYINPUT95), .B2(new_n785), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n720), .A2(new_n716), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT94), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n787), .B(new_n705), .C1(G77), .C2(new_n789), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n374), .A2(new_n376), .B1(new_n375), .B2(new_n657), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n373), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n634), .A2(new_n657), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT96), .ZN(new_n794));
  AND3_X1   g0594(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n794), .B1(new_n792), .B2(new_n793), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n790), .B1(new_n798), .B2(new_n716), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n630), .A2(new_n657), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n798), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n657), .B(new_n797), .C1(new_n627), .C2(new_n629), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n803), .A2(new_n694), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n705), .B1(new_n803), .B2(new_n694), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n799), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(G384));
  INV_X1    g0607(.A(KEYINPUT35), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n242), .B(new_n216), .C1(new_n500), .C2(new_n808), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n809), .A2(KEYINPUT97), .B1(new_n808), .B2(new_n500), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(KEYINPUT97), .B2(new_n809), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT36), .ZN(new_n812));
  OR3_X1    g0612(.A1(new_n386), .A2(new_n217), .A3(new_n260), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n266), .B(G13), .C1(new_n813), .C2(new_n246), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT38), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n388), .B1(new_n396), .B2(new_n399), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n817), .A2(new_n380), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n400), .A2(new_n280), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n404), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n651), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n440), .B1(new_n633), .B2(KEYINPUT72), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n822), .B1(new_n641), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n435), .A2(new_n424), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n651), .B(KEYINPUT98), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n424), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n825), .A2(new_n421), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(KEYINPUT37), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n820), .A2(new_n435), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n830), .A2(new_n822), .A3(new_n421), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n829), .B1(KEYINPUT37), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n816), .B1(new_n824), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n832), .ZN(new_n834));
  OAI211_X1 g0634(.A(KEYINPUT38), .B(new_n834), .C1(new_n442), .C2(new_n822), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n833), .A2(KEYINPUT99), .A3(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT99), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n837), .B(new_n816), .C1(new_n824), .C2(new_n832), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT40), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT102), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n687), .B1(new_n690), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n686), .A2(KEYINPUT102), .A3(KEYINPUT31), .A4(new_n653), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n692), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n349), .A2(new_n657), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n329), .A2(new_n653), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n349), .A2(new_n356), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  AND4_X1   g0648(.A1(new_n839), .A2(new_n844), .A3(new_n797), .A4(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n836), .A2(new_n838), .A3(new_n849), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n424), .B(new_n826), .C1(new_n633), .C2(new_n430), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n828), .B(KEYINPUT37), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT38), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n823), .A2(new_n432), .A3(new_n433), .ZN(new_n854));
  INV_X1    g0654(.A(new_n822), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n832), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n853), .B1(new_n856), .B2(KEYINPUT38), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n844), .A2(new_n848), .A3(new_n797), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT40), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n850), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n860), .A2(new_n443), .A3(new_n844), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(G330), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n443), .A2(G330), .A3(new_n844), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n378), .A2(new_n442), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n676), .B2(new_n699), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n867), .A2(new_n644), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n865), .B(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n349), .A2(new_n653), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n836), .A2(KEYINPUT39), .A3(new_n838), .ZN(new_n872));
  INV_X1    g0672(.A(new_n853), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n835), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT100), .B1(new_n874), .B2(KEYINPUT39), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n836), .A2(KEYINPUT100), .A3(KEYINPUT39), .A4(new_n838), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n871), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n802), .A2(new_n793), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n836), .A2(new_n879), .A3(new_n848), .A4(new_n838), .ZN(new_n880));
  OR3_X1    g0680(.A1(new_n632), .A2(new_n436), .A3(new_n826), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g0683(.A(KEYINPUT101), .B(KEYINPUT103), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n883), .B(new_n884), .ZN(new_n885));
  OAI22_X1  g0685(.A1(new_n869), .A2(new_n885), .B1(new_n266), .B2(new_n647), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n869), .A2(new_n885), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n815), .B1(new_n886), .B2(new_n887), .ZN(G367));
  NAND2_X1  g0688(.A1(new_n485), .A2(new_n653), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n889), .B(KEYINPUT104), .Z(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT105), .B1(new_n890), .B2(new_n615), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n490), .ZN(new_n892));
  MUX2_X1   g0692(.A(new_n891), .B(KEYINPUT105), .S(new_n892), .Z(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n719), .ZN(new_n894));
  INV_X1    g0694(.A(new_n714), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n895), .A2(new_n239), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n721), .B1(new_n208), .B2(new_n460), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n705), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n751), .A2(G311), .B1(new_n763), .B2(G97), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n739), .A2(KEYINPUT46), .A3(G116), .ZN(new_n900));
  INV_X1    g0700(.A(new_n549), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n899), .B(new_n900), .C1(new_n901), .C2(new_n746), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(G317), .B2(new_n728), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT46), .B1(new_n739), .B2(new_n466), .ZN(new_n904));
  INV_X1    g0704(.A(G283), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n734), .A2(new_n573), .B1(new_n744), .B2(new_n905), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n904), .A2(new_n906), .A3(new_n398), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n903), .B(new_n907), .C1(new_n358), .C2(new_n754), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n763), .A2(G77), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n202), .B2(new_n744), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n256), .B(new_n910), .C1(G143), .C2(new_n751), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n731), .A2(G68), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n728), .A2(G137), .ZN(new_n913));
  INV_X1    g0713(.A(G150), .ZN(new_n914));
  INV_X1    g0714(.A(G159), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n914), .A2(new_n746), .B1(new_n734), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(G58), .B2(new_n739), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n911), .A2(new_n912), .A3(new_n913), .A4(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT47), .B1(new_n908), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n919), .A2(new_n770), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n908), .A2(KEYINPUT47), .A3(new_n918), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n898), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n894), .A2(new_n922), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT108), .Z(new_n924));
  OR2_X1    g0724(.A1(new_n656), .A2(new_n662), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n925), .A2(new_n663), .A3(new_n664), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n701), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n533), .A2(new_n657), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n929), .A2(KEYINPUT106), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n534), .B1(new_n505), .B2(new_n657), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n929), .A2(KEYINPUT106), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n666), .A2(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT45), .Z(new_n935));
  NOR2_X1   g0735(.A1(new_n666), .A2(new_n933), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT44), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n935), .A2(new_n663), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n927), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n701), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n668), .B(KEYINPUT41), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n703), .ZN(new_n943));
  INV_X1    g0743(.A(new_n933), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n664), .ZN(new_n945));
  XNOR2_X1  g0745(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n622), .B1(new_n933), .B2(new_n618), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n947), .B1(new_n653), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT43), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n949), .B1(new_n950), .B2(new_n893), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n893), .A2(new_n950), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n951), .B(new_n952), .Z(new_n953));
  NOR2_X1   g0753(.A1(new_n663), .A2(new_n944), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n953), .B(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n924), .B1(new_n943), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(G387));
  NOR2_X1   g0757(.A1(new_n927), .A2(new_n669), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n701), .B2(new_n926), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n655), .A2(new_n719), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n714), .B1(new_n236), .B2(new_n472), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n671), .B2(new_n708), .ZN(new_n962));
  OR3_X1    g0762(.A1(new_n402), .A2(KEYINPUT50), .A3(G50), .ZN(new_n963));
  OAI21_X1  g0763(.A(KEYINPUT50), .B1(new_n402), .B2(G50), .ZN(new_n964));
  AOI211_X1 g0764(.A(G45), .B(new_n670), .C1(G68), .C2(G77), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n962), .A2(new_n966), .B1(new_n358), .B2(new_n209), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n705), .B1(new_n967), .B2(new_n722), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n402), .A2(new_n734), .B1(new_n260), .B2(new_n738), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n746), .A2(new_n202), .B1(new_n744), .B2(new_n226), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n741), .A2(new_n915), .B1(new_n747), .B2(new_n448), .ZN(new_n971));
  NOR4_X1   g0771(.A1(new_n969), .A2(new_n970), .A3(new_n971), .A4(new_n570), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n731), .A2(new_n364), .ZN(new_n973));
  INV_X1    g0773(.A(new_n728), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n972), .B(new_n973), .C1(new_n914), .C2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT109), .ZN(new_n976));
  AOI22_X1  g0776(.A1(G317), .A2(new_n761), .B1(new_n752), .B2(new_n549), .ZN(new_n977));
  INV_X1    g0777(.A(G322), .ZN(new_n978));
  INV_X1    g0778(.A(G311), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n741), .A2(new_n978), .B1(new_n734), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n980), .A2(KEYINPUT110), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(KEYINPUT110), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n977), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT48), .Z(new_n984));
  OAI22_X1  g0784(.A1(new_n754), .A2(new_n905), .B1(new_n573), .B2(new_n738), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n986), .A2(KEYINPUT49), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n570), .B1(new_n539), .B2(new_n747), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(new_n728), .B2(G326), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n986), .B2(KEYINPUT49), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n976), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n968), .B1(new_n991), .B2(new_n720), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n926), .A2(new_n704), .B1(new_n960), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n959), .A2(new_n993), .ZN(G393));
  AOI21_X1  g0794(.A(new_n663), .B1(new_n935), .B2(new_n937), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT111), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(new_n938), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n939), .B(new_n668), .C1(new_n998), .C2(new_n927), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n704), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n721), .B1(new_n448), .B2(new_n208), .C1(new_n895), .C2(new_n245), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n705), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n402), .A2(new_n744), .B1(new_n202), .B2(new_n734), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n738), .A2(new_n226), .B1(new_n747), .B2(new_n221), .ZN(new_n1004));
  NOR3_X1   g0804(.A1(new_n1003), .A2(new_n1004), .A3(new_n570), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT51), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n741), .A2(new_n914), .B1(new_n746), .B2(new_n915), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n728), .A2(G143), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1007), .A2(new_n1006), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n731), .A2(G77), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1005), .A2(new_n1008), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G317), .A2(new_n751), .B1(new_n761), .B2(G311), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT52), .Z(new_n1013));
  OAI22_X1  g0813(.A1(new_n901), .A2(new_n734), .B1(new_n744), .B2(new_n573), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n257), .B(new_n1014), .C1(G107), .C2(new_n763), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1013), .B(new_n1015), .C1(new_n539), .C2(new_n754), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n728), .A2(G322), .B1(G283), .B2(new_n739), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT112), .Z(new_n1018));
  OAI21_X1  g0818(.A(new_n1011), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1002), .B1(new_n1019), .B2(new_n720), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n933), .B2(new_n718), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n999), .A2(new_n1000), .A3(new_n1021), .ZN(G390));
  OAI211_X1 g0822(.A(new_n797), .B(new_n657), .C1(new_n697), .C2(new_n696), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1023), .A2(new_n793), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n848), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n874), .B(new_n871), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n876), .A2(new_n877), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n802), .A2(new_n793), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1028), .A2(new_n1025), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1029), .A2(new_n870), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1026), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(G330), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n858), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n876), .B(new_n877), .C1(new_n870), .C2(new_n1029), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n693), .A2(new_n848), .A3(G330), .A4(new_n797), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1036), .A2(new_n1037), .A3(new_n1026), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n867), .A2(new_n864), .A3(new_n644), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1025), .B1(new_n694), .B2(new_n798), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1028), .B1(new_n1033), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n844), .A2(G330), .A3(new_n797), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n1025), .ZN(new_n1044));
  AND3_X1   g0844(.A1(new_n1024), .A2(new_n1044), .A3(new_n1037), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1040), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(KEYINPUT113), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT113), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1040), .B(new_n1048), .C1(new_n1042), .C2(new_n1045), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n669), .B1(new_n1039), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1035), .A2(new_n1052), .A3(new_n1038), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n876), .A2(new_n716), .A3(new_n877), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n705), .B1(new_n789), .B2(new_n288), .ZN(new_n1056));
  INV_X1    g0856(.A(G132), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n738), .A2(new_n914), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT53), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n257), .B1(new_n1057), .B2(new_n746), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n1059), .B2(new_n1058), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n731), .A2(G159), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n728), .A2(G125), .ZN(new_n1063));
  XOR2_X1   g0863(.A(KEYINPUT54), .B(G143), .Z(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(G137), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n1065), .A2(new_n744), .B1(new_n1066), .B2(new_n734), .ZN(new_n1067));
  INV_X1    g0867(.A(G128), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n741), .A2(new_n1068), .B1(new_n747), .B2(new_n202), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .A4(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n751), .A2(G283), .B1(new_n752), .B2(G97), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n358), .B2(new_n734), .C1(new_n242), .C2(new_n746), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n257), .B(new_n1073), .C1(G87), .C2(new_n739), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n974), .A2(new_n573), .B1(new_n226), .B2(new_n747), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT114), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1074), .A2(new_n1010), .A3(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1071), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1056), .B1(new_n1080), .B2(new_n720), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1055), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n1039), .B2(new_n703), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1054), .A2(new_n1084), .ZN(G378));
  NOR2_X1   g0885(.A1(new_n298), .A2(new_n651), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n316), .B1(new_n307), .B2(new_n312), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(KEYINPUT55), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1087), .A2(KEYINPUT55), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1086), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT55), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n318), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1086), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1094), .A2(new_n1095), .A3(new_n1088), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n1091), .A2(new_n1092), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1092), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n716), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(G33), .A2(G41), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT115), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n202), .B(new_n1102), .C1(new_n398), .C2(G41), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n741), .A2(new_n242), .B1(new_n738), .B2(new_n260), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n460), .A2(new_n744), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n448), .A2(new_n734), .B1(new_n746), .B2(new_n358), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n747), .A2(new_n224), .ZN(new_n1107));
  NOR4_X1   g0907(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  AOI211_X1 g0908(.A(G41), .B(new_n398), .C1(new_n728), .C2(G283), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n1108), .A2(new_n1109), .A3(new_n912), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1103), .B1(new_n1110), .B2(KEYINPUT58), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT116), .ZN(new_n1112));
  OR2_X1    g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n739), .A2(new_n1064), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT117), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n731), .A2(G150), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G128), .A2(new_n761), .B1(new_n752), .B2(G137), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(G125), .A2(new_n751), .B1(new_n735), .B2(G132), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n1120), .A2(KEYINPUT59), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1102), .B1(G159), .B2(new_n763), .ZN(new_n1122));
  INV_X1    g0922(.A(G124), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1122), .B1(new_n974), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n1120), .B2(KEYINPUT59), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1121), .A2(new_n1125), .B1(KEYINPUT58), .B2(new_n1110), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1113), .A2(new_n1114), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n720), .ZN(new_n1128));
  OR2_X1    g0928(.A1(new_n789), .A2(G50), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1100), .A2(new_n705), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1027), .A2(new_n870), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n862), .A2(new_n1099), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n882), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1099), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n860), .A2(new_n1135), .A3(G330), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1032), .B(new_n1099), .C1(new_n850), .C2(new_n859), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1135), .B1(new_n860), .B2(G330), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1138), .A2(new_n1139), .B1(new_n878), .B2(new_n882), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1137), .A2(KEYINPUT119), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT119), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n883), .A2(new_n1142), .A3(new_n1133), .A4(new_n1136), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1131), .B1(new_n1144), .B2(new_n704), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1053), .A2(new_n1040), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT57), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1040), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n1036), .A2(new_n1037), .A3(new_n1026), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1033), .B1(new_n1036), .B2(new_n1026), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1148), .B1(new_n1151), .B2(new_n1052), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(KEYINPUT57), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n668), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1145), .B1(new_n1147), .B2(new_n1155), .ZN(G375));
  OAI21_X1  g0956(.A(new_n705), .B1(new_n789), .B2(G68), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n1065), .A2(new_n734), .B1(new_n1066), .B2(new_n746), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n741), .A2(new_n1057), .B1(new_n744), .B2(new_n914), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n738), .A2(new_n915), .B1(new_n747), .B2(new_n224), .ZN(new_n1160));
  NOR4_X1   g0960(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n570), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1161), .B1(new_n202), .B2(new_n754), .C1(new_n1068), .C2(new_n974), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n448), .A2(new_n738), .B1(new_n746), .B2(new_n905), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(G294), .B2(new_n751), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n973), .A2(new_n1164), .A3(new_n256), .A4(new_n909), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n466), .A2(new_n735), .B1(new_n752), .B2(G107), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1167), .A2(KEYINPUT120), .B1(G303), .B2(new_n728), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(KEYINPUT120), .B2(new_n1167), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1162), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1157), .B1(new_n1170), .B2(new_n720), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n716), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1171), .B1(new_n848), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1173), .B1(new_n1174), .B2(new_n703), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(new_n1148), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n941), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1176), .B1(new_n1052), .B2(new_n1178), .ZN(G381));
  INV_X1    g0979(.A(KEYINPUT121), .ZN(new_n1180));
  AOI21_X1  g0980(.A(G378), .B1(G375), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n1180), .B2(G375), .ZN(new_n1182));
  INV_X1    g0982(.A(G390), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(G393), .A2(G396), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n956), .A2(new_n806), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  OR3_X1    g0985(.A1(new_n1182), .A2(G381), .A3(new_n1185), .ZN(G407));
  NAND2_X1  g0986(.A1(new_n652), .A2(G213), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT122), .ZN(new_n1188));
  OAI211_X1 g0988(.A(G407), .B(G213), .C1(new_n1182), .C2(new_n1188), .ZN(G409));
  INV_X1    g0989(.A(new_n1188), .ZN(new_n1190));
  OAI211_X1 g0990(.A(G378), .B(new_n1145), .C1(new_n1147), .C2(new_n1155), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1146), .A2(new_n941), .A3(new_n1143), .A4(new_n1141), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT123), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n703), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1193), .B1(new_n1194), .B2(new_n1131), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1153), .A2(new_n704), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1196), .A2(KEYINPUT123), .A3(new_n1130), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1192), .A2(new_n1195), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1083), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1190), .B1(new_n1191), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1050), .A2(KEYINPUT60), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n1177), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1174), .A2(KEYINPUT60), .A3(new_n1148), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT125), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n669), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1203), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1208), .A2(G384), .A3(new_n1176), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n1177), .B2(new_n1202), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n806), .B1(new_n1211), .B2(new_n1175), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1209), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1201), .A2(KEYINPUT63), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(G387), .A2(new_n1183), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n956), .A2(G390), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  AND2_X1   g1017(.A1(G393), .A2(G396), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1217), .B1(new_n1184), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT61), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1218), .A2(new_n1184), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1215), .A2(new_n1221), .A3(new_n1216), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1214), .A2(new_n1219), .A3(new_n1220), .A4(new_n1222), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1191), .A2(new_n1200), .A3(KEYINPUT124), .ZN(new_n1224));
  AOI21_X1  g1024(.A(KEYINPUT124), .B1(new_n1191), .B2(new_n1200), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1187), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(G2897), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1209), .A2(new_n1212), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1190), .A2(G2897), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1229), .B1(new_n1213), .B2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(KEYINPUT63), .B1(new_n1227), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1227), .A2(new_n1213), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1223), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1220), .B1(new_n1231), .B2(new_n1201), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT62), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n1201), .B2(new_n1213), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1191), .A2(new_n1200), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT124), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1226), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1191), .A2(new_n1200), .A3(KEYINPUT124), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1241), .A2(new_n1236), .A3(new_n1213), .A4(new_n1242), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1238), .A2(new_n1243), .B1(new_n1222), .B2(new_n1219), .ZN(new_n1244));
  OAI21_X1  g1044(.A(KEYINPUT126), .B1(new_n1234), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1223), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT63), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1229), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1230), .B1(new_n1209), .B2(new_n1212), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1247), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1209), .A2(new_n1212), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1248), .A2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1246), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1219), .A2(new_n1222), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1243), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1239), .A2(new_n1188), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT61), .B1(new_n1251), .B2(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(KEYINPUT62), .B1(new_n1258), .B2(new_n1253), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1256), .B1(new_n1257), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT126), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1255), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1245), .A2(new_n1264), .ZN(G405));
  INV_X1    g1065(.A(KEYINPUT127), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1191), .B1(new_n1253), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(new_n1199), .B2(G375), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1213), .A2(KEYINPUT127), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1268), .B(new_n1269), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1270), .B(new_n1256), .ZN(G402));
endmodule


