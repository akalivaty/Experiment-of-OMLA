//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G210), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT70), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G101), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  OR2_X1    g007(.A1(KEYINPUT2), .A2(G113), .ZN(new_n194));
  AND3_X1   g008(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n195));
  AOI21_X1  g009(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n194), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  XOR2_X1   g011(.A(G116), .B(G119), .Z(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(G116), .B(G119), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n200), .B(new_n194), .C1(new_n196), .C2(new_n195), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G137), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G134), .ZN(new_n207));
  AND3_X1   g021(.A1(new_n205), .A2(new_n207), .A3(KEYINPUT65), .ZN(new_n208));
  OAI21_X1  g022(.A(G131), .B1(new_n207), .B2(KEYINPUT65), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n203), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G143), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G146), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n212), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(KEYINPUT1), .A3(G146), .ZN(new_n218));
  XNOR2_X1  g032(.A(G143), .B(G146), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n217), .B(new_n218), .C1(G128), .C2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT11), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n221), .B1(new_n204), .B2(G137), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n206), .A2(KEYINPUT11), .A3(G134), .ZN(new_n223));
  INV_X1    g037(.A(G131), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n205), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n205), .A2(new_n207), .A3(KEYINPUT65), .ZN(new_n226));
  OR3_X1    g040(.A1(new_n204), .A2(KEYINPUT65), .A3(G137), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT66), .A4(G131), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n210), .A2(new_n220), .A3(new_n225), .A4(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n222), .A2(new_n205), .A3(new_n223), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G131), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n225), .ZN(new_n232));
  AND2_X1   g046(.A1(KEYINPUT0), .A2(G128), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n214), .A2(new_n216), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT0), .B(G128), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n234), .B1(new_n219), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n232), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n229), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT30), .B1(new_n239), .B2(KEYINPUT64), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT64), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT30), .ZN(new_n242));
  AOI211_X1 g056(.A(new_n241), .B(new_n242), .C1(new_n229), .C2(new_n238), .ZN(new_n243));
  OAI211_X1 g057(.A(KEYINPUT68), .B(new_n202), .C1(new_n240), .C2(new_n243), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n199), .A2(new_n201), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n236), .B1(new_n231), .B2(new_n225), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n212), .A2(new_n214), .A3(new_n216), .ZN(new_n247));
  AOI21_X1  g061(.A(G128), .B1(new_n214), .B2(new_n216), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n226), .A2(new_n227), .A3(G131), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n249), .A2(new_n218), .B1(new_n203), .B2(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n228), .A2(new_n225), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n246), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n242), .B1(new_n253), .B2(new_n241), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n239), .A2(KEYINPUT64), .A3(KEYINPUT30), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n245), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n239), .A2(new_n202), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n193), .B(new_n244), .C1(new_n256), .C2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT31), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n240), .A2(new_n243), .ZN(new_n263));
  OAI22_X1  g077(.A1(new_n263), .A2(new_n245), .B1(new_n258), .B2(new_n257), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n264), .A2(KEYINPUT31), .A3(new_n193), .A4(new_n244), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT28), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n257), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n268), .A2(KEYINPUT71), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n253), .A2(new_n245), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n271), .B1(new_n239), .B2(new_n202), .ZN(new_n272));
  AOI211_X1 g086(.A(KEYINPUT72), .B(new_n245), .C1(new_n229), .C2(new_n238), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n270), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT71), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n269), .B1(new_n276), .B2(KEYINPUT28), .ZN(new_n277));
  INV_X1    g091(.A(new_n193), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n266), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(G472), .A2(G902), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(KEYINPUT32), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT32), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n262), .A2(new_n265), .B1(new_n277), .B2(new_n278), .ZN(new_n284));
  INV_X1    g098(.A(new_n281), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n269), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n239), .A2(new_n202), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT72), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n239), .A2(new_n271), .A3(new_n202), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT71), .B1(new_n291), .B2(new_n270), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n287), .B(new_n193), .C1(new_n292), .C2(new_n267), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n264), .A2(new_n278), .A3(new_n244), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT29), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n270), .A2(new_n288), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n268), .B1(new_n296), .B2(new_n267), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n297), .A2(KEYINPUT29), .A3(new_n193), .ZN(new_n298));
  INV_X1    g112(.A(G902), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G472), .B1(new_n295), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n282), .A2(new_n286), .A3(new_n301), .ZN(new_n302));
  OR2_X1    g116(.A1(KEYINPUT24), .A2(G110), .ZN(new_n303));
  NAND2_X1  g117(.A1(KEYINPUT24), .A2(G110), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(G119), .B(G128), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n303), .A2(KEYINPUT73), .A3(new_n304), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(KEYINPUT74), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT75), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n312), .A2(G125), .A3(G140), .ZN(new_n313));
  AOI21_X1  g127(.A(G140), .B1(new_n312), .B2(G125), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT16), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G125), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n316), .A2(KEYINPUT16), .A3(G140), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(G146), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(new_n316), .B2(KEYINPUT75), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n312), .A2(G125), .A3(G140), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n324), .A2(new_n213), .A3(new_n317), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n319), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT23), .ZN(new_n328));
  INV_X1    g142(.A(G119), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n328), .B1(new_n329), .B2(G128), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n211), .A2(KEYINPUT23), .A3(G119), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n330), .B(new_n331), .C1(G119), .C2(new_n211), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G110), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n311), .A2(new_n327), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n315), .A2(G146), .A3(new_n318), .ZN(new_n335));
  XNOR2_X1  g149(.A(G125), .B(G140), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n213), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n308), .B1(new_n307), .B2(new_n309), .ZN(new_n338));
  XOR2_X1   g152(.A(KEYINPUT76), .B(G110), .Z(new_n339));
  NOR2_X1   g153(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n335), .B(new_n337), .C1(new_n338), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n334), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(G221), .A2(G234), .ZN(new_n343));
  OR3_X1    g157(.A1(new_n343), .A2(KEYINPUT77), .A3(G953), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT22), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT77), .B1(new_n343), .B2(G953), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n345), .B1(new_n344), .B2(new_n346), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n206), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n349), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n347), .A3(G137), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n342), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n353), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n334), .A2(new_n341), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n299), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT25), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n354), .A2(KEYINPUT25), .A3(new_n299), .A4(new_n356), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G234), .ZN(new_n362));
  OAI21_X1  g176(.A(G217), .B1(new_n362), .B2(G902), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n356), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n355), .B1(new_n334), .B2(new_n341), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n364), .A2(G902), .ZN(new_n369));
  XOR2_X1   g183(.A(new_n369), .B(KEYINPUT78), .Z(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n365), .A2(KEYINPUT79), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT79), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n363), .B1(new_n359), .B2(new_n360), .ZN(new_n375));
  INV_X1    g189(.A(new_n372), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n379));
  AOI21_X1  g193(.A(G143), .B1(new_n187), .B2(G214), .ZN(new_n380));
  OAI21_X1  g194(.A(G131), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT17), .ZN(new_n382));
  INV_X1    g196(.A(G237), .ZN(new_n383));
  INV_X1    g197(.A(G953), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(G214), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n215), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n224), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n381), .A2(new_n382), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT91), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OAI211_X1 g205(.A(KEYINPUT17), .B(G131), .C1(new_n379), .C2(new_n380), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT90), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n386), .A2(new_n387), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n395), .A2(KEYINPUT90), .A3(KEYINPUT17), .A4(G131), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n381), .A2(new_n388), .A3(KEYINPUT91), .A4(new_n382), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n391), .A2(new_n397), .A3(new_n326), .A4(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(G113), .B(G122), .ZN(new_n400));
  INV_X1    g214(.A(G104), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n400), .B(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n322), .A2(G146), .A3(new_n323), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n337), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT88), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT88), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n337), .A2(new_n406), .A3(new_n403), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT89), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT18), .ZN(new_n410));
  OAI22_X1  g224(.A1(new_n395), .A2(new_n409), .B1(new_n410), .B2(new_n224), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n410), .A2(new_n224), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n386), .A2(KEYINPUT89), .A3(new_n412), .A4(new_n387), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n399), .A2(new_n402), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n402), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n407), .A2(new_n405), .B1(new_n411), .B2(new_n413), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n381), .A2(new_n388), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n336), .A2(KEYINPUT19), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT19), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n322), .B2(new_n323), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n213), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n419), .A2(new_n335), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n417), .B1(new_n418), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n416), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G475), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n299), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n399), .A2(new_n402), .A3(new_n415), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n402), .B1(new_n399), .B2(new_n415), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n299), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G475), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n426), .A2(KEYINPUT20), .A3(new_n427), .A4(new_n299), .ZN(new_n435));
  INV_X1    g249(.A(G478), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(KEYINPUT15), .ZN(new_n437));
  INV_X1    g251(.A(G116), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n438), .A2(G122), .ZN(new_n439));
  INV_X1    g253(.A(G122), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(G116), .ZN(new_n441));
  OAI21_X1  g255(.A(G107), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(G116), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n438), .A2(G122), .ZN(new_n444));
  INV_X1    g258(.A(G107), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT13), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(new_n211), .B2(G143), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n211), .A2(G143), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n215), .A2(KEYINPUT13), .A3(G128), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G134), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n215), .A2(G128), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(new_n450), .A3(new_n204), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n447), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT14), .B1(new_n438), .B2(G122), .ZN(new_n457));
  OAI211_X1 g271(.A(G107), .B(new_n457), .C1(new_n439), .C2(new_n441), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n443), .B(new_n444), .C1(KEYINPUT14), .C2(new_n445), .ZN(new_n459));
  INV_X1    g273(.A(new_n455), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n204), .B1(new_n454), .B2(new_n450), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n458), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(KEYINPUT9), .A2(G234), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(KEYINPUT9), .A2(G234), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n464), .A2(KEYINPUT80), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT80), .ZN(new_n467));
  INV_X1    g281(.A(new_n465), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n467), .B1(new_n468), .B2(new_n463), .ZN(new_n469));
  AND4_X1   g283(.A1(G217), .A2(new_n466), .A3(new_n469), .A4(new_n384), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n456), .A2(new_n462), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n470), .B1(new_n456), .B2(new_n462), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n299), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT92), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n437), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n474), .ZN(new_n476));
  OAI211_X1 g290(.A(KEYINPUT92), .B(new_n299), .C1(new_n471), .C2(new_n472), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n475), .B1(new_n478), .B2(new_n437), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n430), .A2(new_n434), .A3(new_n435), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(G234), .A2(G237), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(G952), .A3(new_n384), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  XOR2_X1   g297(.A(KEYINPUT21), .B(G898), .Z(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n481), .A2(G902), .A3(G953), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n483), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n480), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT83), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT3), .B1(new_n401), .B2(G107), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT3), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n445), .A3(G104), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n401), .A2(G107), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G101), .ZN(new_n496));
  INV_X1    g310(.A(G101), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n491), .A2(new_n493), .A3(new_n497), .A4(new_n494), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(KEYINPUT4), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n495), .A2(new_n500), .A3(G101), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n237), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT10), .ZN(new_n503));
  INV_X1    g317(.A(new_n218), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n247), .A2(new_n248), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n445), .A2(KEYINPUT82), .A3(G104), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT82), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(new_n401), .B2(G107), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n445), .A2(G104), .ZN(new_n509));
  OAI211_X1 g323(.A(G101), .B(new_n506), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n498), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n503), .B1(new_n505), .B2(new_n511), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n510), .A2(new_n498), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(KEYINPUT10), .A3(new_n220), .ZN(new_n514));
  INV_X1    g328(.A(new_n232), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n502), .A2(new_n512), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n511), .B(new_n220), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT12), .ZN(new_n518));
  NOR3_X1   g332(.A1(new_n517), .A2(new_n518), .A3(new_n515), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n513), .A2(new_n220), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n505), .A2(new_n511), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT12), .B1(new_n522), .B2(new_n232), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n516), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(G110), .B(G140), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n384), .A2(G227), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n516), .A2(new_n527), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n502), .A2(new_n512), .A3(new_n514), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n232), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n524), .A2(new_n528), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n490), .B(G469), .C1(new_n533), .C2(G902), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n466), .A2(new_n469), .A3(new_n299), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(G221), .ZN(new_n536));
  XOR2_X1   g350(.A(new_n536), .B(KEYINPUT81), .Z(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(G214), .B1(G237), .B2(G902), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(KEYINPUT84), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n499), .A2(new_n202), .A3(new_n501), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT5), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(new_n329), .A3(G116), .ZN(new_n545));
  OAI211_X1 g359(.A(G113), .B(new_n545), .C1(new_n198), .C2(new_n544), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n513), .A2(new_n201), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(G110), .B(G122), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n543), .A2(new_n547), .A3(new_n549), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(KEYINPUT6), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n248), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n554), .A2(new_n316), .A3(new_n218), .A4(new_n217), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n236), .A2(G125), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G224), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(G953), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n557), .B(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT6), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n548), .A2(new_n561), .A3(new_n550), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n553), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n549), .B(KEYINPUT8), .Z(new_n564));
  NAND2_X1  g378(.A1(new_n546), .A2(new_n201), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n511), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n564), .B1(new_n566), .B2(new_n547), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n557), .A2(new_n559), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n567), .B1(KEYINPUT7), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n559), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n555), .A2(new_n556), .B1(KEYINPUT7), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(KEYINPUT85), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n552), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n563), .A2(new_n573), .A3(new_n299), .ZN(new_n574));
  OAI21_X1  g388(.A(G210), .B1(G237), .B2(G902), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT86), .ZN(new_n576));
  XOR2_X1   g390(.A(new_n576), .B(KEYINPUT87), .Z(new_n577));
  NAND2_X1  g391(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n576), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n563), .A2(new_n573), .A3(new_n299), .A4(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n542), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(G469), .B1(new_n533), .B2(G902), .ZN(new_n582));
  INV_X1    g396(.A(G469), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n522), .A2(KEYINPUT12), .A3(new_n232), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n518), .B1(new_n517), .B2(new_n515), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n529), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n527), .B1(new_n532), .B2(new_n516), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n583), .B(new_n299), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n582), .A2(KEYINPUT83), .A3(new_n588), .ZN(new_n589));
  AND4_X1   g403(.A1(new_n489), .A2(new_n539), .A3(new_n581), .A4(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n302), .A2(new_n378), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G101), .ZN(G3));
  INV_X1    g406(.A(KEYINPUT93), .ZN(new_n593));
  INV_X1    g407(.A(G472), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n280), .A2(new_n299), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n595), .B1(new_n284), .B2(G902), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n589), .A2(new_n538), .A3(new_n534), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n599), .A2(KEYINPUT94), .A3(new_n378), .A4(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n378), .A2(new_n597), .A3(new_n600), .A4(new_n598), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT94), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n430), .A2(new_n434), .A3(new_n435), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n473), .A2(new_n436), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n456), .A2(new_n462), .ZN(new_n608));
  INV_X1    g422(.A(new_n470), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n456), .A2(new_n462), .A3(new_n470), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT33), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n299), .A2(G478), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n607), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n606), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(new_n488), .ZN(new_n618));
  INV_X1    g432(.A(new_n540), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n574), .A2(new_n576), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n619), .B1(new_n620), .B2(new_n580), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n605), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT34), .B(G104), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  AND3_X1   g438(.A1(new_n430), .A2(new_n434), .A3(new_n435), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT92), .B1(new_n612), .B2(new_n299), .ZN(new_n626));
  INV_X1    g440(.A(new_n477), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n437), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n475), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n488), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n625), .A2(KEYINPUT95), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT95), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n430), .A2(new_n630), .A3(new_n434), .A4(new_n435), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n633), .B1(new_n634), .B2(new_n488), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n605), .A2(new_n621), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n637), .B(KEYINPUT96), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT35), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(new_n445), .ZN(G9));
  INV_X1    g454(.A(KEYINPUT97), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n342), .B(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n353), .A2(KEYINPUT36), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n365), .B1(new_n645), .B2(new_n370), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n590), .A2(new_n597), .A3(new_n646), .A4(new_n598), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT37), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(G110), .Z(G12));
  AND3_X1   g463(.A1(new_n302), .A2(new_n621), .A3(new_n646), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n486), .A2(G900), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n482), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n634), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n650), .A2(KEYINPUT98), .A3(new_n600), .A4(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT98), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n302), .A2(new_n600), .A3(new_n621), .A4(new_n646), .ZN(new_n657));
  INV_X1    g471(.A(new_n654), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  NOR2_X1   g475(.A1(new_n625), .A2(new_n479), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n540), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n646), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n664), .B(KEYINPUT99), .Z(new_n665));
  NAND2_X1  g479(.A1(new_n264), .A2(new_n244), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n193), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n299), .B1(new_n193), .B2(new_n296), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n282), .A2(new_n286), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n578), .A2(new_n580), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT38), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n652), .B(KEYINPUT39), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n600), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT40), .ZN(new_n677));
  NOR4_X1   g491(.A1(new_n665), .A2(new_n672), .A3(new_n674), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(new_n215), .ZN(G45));
  NOR2_X1   g493(.A1(new_n617), .A2(new_n653), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n657), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(new_n213), .ZN(G48));
  OAI21_X1  g497(.A(new_n299), .B1(new_n586), .B2(new_n587), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(G469), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n538), .A3(new_n588), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT100), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n685), .A2(KEYINPUT100), .A3(new_n538), .A4(new_n588), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n688), .A2(new_n621), .A3(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n302), .A2(new_n378), .A3(new_n618), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT101), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT41), .B(G113), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  NAND4_X1  g508(.A1(new_n302), .A2(new_n378), .A3(new_n636), .A4(new_n690), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  AND3_X1   g510(.A1(new_n688), .A2(new_n489), .A3(new_n689), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n302), .A2(new_n621), .A3(new_n646), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G119), .ZN(G21));
  AND4_X1   g513(.A1(new_n621), .A2(new_n662), .A3(new_n688), .A4(new_n689), .ZN(new_n700));
  OR2_X1    g514(.A1(new_n297), .A2(new_n193), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n285), .B1(new_n266), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n280), .A2(new_n299), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n702), .B1(new_n703), .B2(G472), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n375), .A2(new_n376), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n700), .A2(new_n704), .A3(new_n705), .A4(new_n631), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G122), .ZN(G24));
  NAND4_X1  g521(.A1(new_n704), .A2(new_n646), .A3(new_n680), .A4(new_n690), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G125), .ZN(G27));
  NAND2_X1  g523(.A1(new_n302), .A2(new_n705), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT42), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n578), .A2(new_n580), .A3(new_n540), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n537), .B1(new_n582), .B2(new_n588), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR4_X1   g528(.A1(new_n710), .A2(new_n711), .A3(new_n681), .A4(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n714), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n302), .A2(new_n378), .A3(new_n680), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n711), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT102), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n717), .A2(new_n720), .A3(new_n711), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n715), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n224), .ZN(G33));
  NAND4_X1  g537(.A1(new_n302), .A2(new_n378), .A3(new_n654), .A4(new_n716), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G134), .ZN(G36));
  INV_X1    g539(.A(new_n588), .ZN(new_n726));
  XOR2_X1   g540(.A(new_n533), .B(KEYINPUT45), .Z(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(G469), .ZN(new_n728));
  NAND2_X1  g542(.A1(G469), .A2(G902), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT46), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n726), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n728), .A2(KEYINPUT46), .A3(new_n729), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n537), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n675), .ZN(new_n735));
  XOR2_X1   g549(.A(new_n735), .B(KEYINPUT103), .Z(new_n736));
  INV_X1    g550(.A(new_n712), .ZN(new_n737));
  INV_X1    g551(.A(new_n599), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n625), .A2(new_n616), .ZN(new_n739));
  XOR2_X1   g553(.A(new_n739), .B(KEYINPUT43), .Z(new_n740));
  NAND3_X1  g554(.A1(new_n738), .A2(new_n646), .A3(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n737), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n736), .B(new_n743), .C1(new_n742), .C2(new_n741), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT104), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n206), .ZN(G39));
  NOR4_X1   g560(.A1(new_n302), .A2(new_n378), .A3(new_n681), .A4(new_n737), .ZN(new_n747));
  XOR2_X1   g561(.A(new_n747), .B(KEYINPUT105), .Z(new_n748));
  XNOR2_X1  g562(.A(new_n734), .B(KEYINPUT47), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(KEYINPUT106), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n321), .ZN(G42));
  OAI21_X1  g566(.A(new_n708), .B1(new_n657), .B2(new_n681), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n753), .B1(new_n655), .B2(new_n659), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n663), .B1(new_n580), .B2(new_n620), .ZN(new_n755));
  XOR2_X1   g569(.A(new_n652), .B(KEYINPUT112), .Z(new_n756));
  NOR2_X1   g570(.A1(new_n646), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n755), .A2(new_n671), .A3(new_n757), .A4(new_n713), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n754), .A2(KEYINPUT52), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT52), .B1(new_n754), .B2(new_n758), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AND4_X1   g575(.A1(new_n691), .A2(new_n706), .A3(new_n695), .A4(new_n698), .ZN(new_n762));
  AOI211_X1 g576(.A(new_n488), .B(new_n542), .C1(new_n578), .C2(new_n580), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n634), .A2(KEYINPUT108), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n634), .A2(KEYINPUT108), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n617), .A2(KEYINPUT107), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT107), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n770), .B1(new_n606), .B2(new_n616), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n763), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  OAI211_X1 g586(.A(KEYINPUT109), .B(new_n763), .C1(new_n764), .C2(new_n765), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n768), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n601), .A2(new_n774), .A3(new_n604), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n591), .A2(new_n647), .ZN(new_n776));
  OAI21_X1  g590(.A(KEYINPUT110), .B1(new_n480), .B2(new_n653), .ZN(new_n777));
  AND4_X1   g591(.A1(new_n539), .A2(new_n777), .A3(new_n589), .A4(new_n712), .ZN(new_n778));
  OR3_X1    g592(.A1(new_n480), .A2(KEYINPUT110), .A3(new_n653), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n302), .A2(new_n778), .A3(new_n779), .A4(new_n646), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n704), .A2(new_n646), .A3(new_n680), .A4(new_n716), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n780), .A2(new_n724), .A3(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n762), .A2(new_n775), .A3(new_n776), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n722), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n761), .A2(KEYINPUT53), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT111), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n786), .B1(new_n783), .B2(new_n722), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n775), .A2(new_n776), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n691), .A2(new_n706), .A3(new_n695), .A4(new_n698), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n710), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n791), .A2(KEYINPUT42), .A3(new_n680), .A4(new_n716), .ZN(new_n792));
  INV_X1    g606(.A(new_n721), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n720), .B1(new_n717), .B2(new_n711), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n790), .A2(KEYINPUT111), .A3(new_n795), .A4(new_n782), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n787), .B(new_n796), .C1(new_n759), .C2(new_n760), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n797), .A2(KEYINPUT113), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT113), .B1(new_n797), .B2(new_n798), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n785), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n801), .A2(KEYINPUT54), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n797), .B(new_n798), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT54), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n384), .A2(G952), .ZN(new_n805));
  INV_X1    g619(.A(new_n378), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n688), .A2(new_n689), .A3(new_n712), .ZN(new_n807));
  NOR4_X1   g621(.A1(new_n671), .A2(new_n806), .A3(new_n482), .A4(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n617), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n805), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n740), .A2(new_n483), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n688), .A2(new_n689), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n704), .A2(new_n705), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n621), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n619), .A3(new_n674), .ZN(new_n816));
  XOR2_X1   g630(.A(new_n816), .B(KEYINPUT50), .Z(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT51), .ZN(new_n818));
  INV_X1    g632(.A(new_n808), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n819), .A2(new_n606), .A3(new_n616), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n704), .A2(new_n646), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n811), .A2(new_n807), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n811), .A2(new_n813), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n685), .A2(new_n588), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n538), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n712), .B(new_n824), .C1(new_n749), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n810), .B(new_n815), .C1(new_n818), .C2(new_n828), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n817), .A2(KEYINPUT114), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n817), .A2(KEYINPUT114), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n830), .A2(new_n831), .A3(new_n823), .A4(new_n827), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n829), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n822), .A2(new_n791), .ZN(new_n835));
  XOR2_X1   g649(.A(KEYINPUT115), .B(KEYINPUT48), .Z(new_n836));
  XNOR2_X1  g650(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n802), .A2(new_n804), .A3(new_n834), .A4(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n838), .B1(G952), .B2(G953), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n739), .A2(new_n542), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n674), .A2(new_n705), .A3(new_n538), .A4(new_n840), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n841), .A2(new_n671), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n825), .B(KEYINPUT49), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(G75));
  NAND2_X1  g658(.A1(new_n553), .A2(new_n562), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(new_n560), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT55), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT56), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n801), .A2(new_n850), .A3(G902), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n850), .B1(new_n801), .B2(G902), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n849), .B1(new_n853), .B2(new_n577), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n384), .A2(G952), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n801), .A2(G902), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT56), .B1(new_n857), .B2(new_n576), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n856), .B1(new_n858), .B2(new_n847), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n854), .A2(new_n859), .ZN(G51));
  NAND3_X1  g674(.A1(new_n853), .A2(G469), .A3(new_n727), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n801), .B(KEYINPUT54), .Z(new_n862));
  XNOR2_X1  g676(.A(new_n729), .B(KEYINPUT57), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n862), .A2(new_n863), .B1(new_n587), .B2(new_n586), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n855), .B1(new_n861), .B2(new_n864), .ZN(G54));
  OAI211_X1 g679(.A(KEYINPUT58), .B(G475), .C1(new_n851), .C2(new_n852), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n867));
  INV_X1    g681(.A(new_n426), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n856), .B1(new_n866), .B2(new_n868), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n867), .B1(new_n866), .B2(new_n868), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(G60));
  XNOR2_X1  g686(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n873));
  NAND2_X1  g687(.A1(G478), .A2(G902), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n873), .B(new_n874), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n862), .A2(new_n614), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n875), .B1(new_n802), .B2(new_n804), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n856), .B1(new_n877), .B2(new_n613), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n876), .A2(new_n878), .ZN(G63));
  NAND2_X1  g693(.A1(G217), .A2(G902), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT60), .Z(new_n881));
  XOR2_X1   g695(.A(new_n644), .B(KEYINPUT119), .Z(new_n882));
  NAND3_X1  g696(.A1(new_n801), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n856), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n368), .B1(new_n801), .B2(new_n881), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n886));
  OAI22_X1  g700(.A1(new_n884), .A2(new_n885), .B1(KEYINPUT120), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(KEYINPUT120), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT121), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n887), .B(new_n889), .ZN(G66));
  OAI21_X1  g704(.A(G953), .B1(new_n485), .B2(new_n558), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n891), .B1(new_n790), .B2(G953), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n845), .B1(G898), .B2(new_n384), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT122), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n892), .B(new_n894), .ZN(G69));
  NOR2_X1   g709(.A1(new_n420), .A2(new_n422), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n263), .B(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT123), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n897), .A2(KEYINPUT123), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n744), .A2(new_n750), .ZN(new_n900));
  INV_X1    g714(.A(new_n754), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(new_n678), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT62), .ZN(new_n903));
  OR4_X1    g717(.A1(new_n771), .A2(new_n769), .A3(new_n764), .A4(new_n765), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n905), .A2(KEYINPUT124), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n676), .B1(new_n905), .B2(KEYINPUT124), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n302), .A2(new_n378), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n906), .A2(new_n907), .A3(new_n909), .A4(new_n712), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n900), .A2(new_n903), .A3(new_n910), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT125), .Z(new_n912));
  OAI211_X1 g726(.A(new_n898), .B(new_n899), .C1(new_n912), .C2(G953), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n384), .B1(G227), .B2(G900), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n384), .A2(G900), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n754), .A2(new_n724), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n736), .A2(new_n791), .A3(new_n755), .ZN(new_n918));
  AND4_X1   g732(.A1(new_n795), .A2(new_n900), .A3(new_n917), .A4(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n916), .B1(new_n919), .B2(G953), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(KEYINPUT126), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n922), .B(new_n916), .C1(new_n919), .C2(G953), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n921), .A2(new_n897), .A3(new_n923), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n913), .A2(new_n914), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n914), .B1(new_n913), .B2(new_n924), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(G72));
  NAND2_X1  g741(.A1(new_n912), .A2(new_n790), .ZN(new_n928));
  NAND2_X1  g742(.A1(G472), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT63), .Z(new_n930));
  AOI21_X1  g744(.A(new_n667), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n919), .A2(new_n790), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n294), .B1(new_n932), .B2(new_n930), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n667), .A2(new_n294), .A3(new_n930), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT127), .Z(new_n935));
  AND2_X1   g749(.A1(new_n803), .A2(new_n935), .ZN(new_n936));
  NOR4_X1   g750(.A1(new_n931), .A2(new_n855), .A3(new_n933), .A4(new_n936), .ZN(G57));
endmodule


