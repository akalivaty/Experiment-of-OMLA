//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 1 0 1 0 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(KEYINPUT3), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT76), .A2(G107), .ZN(new_n191));
  NOR2_X1   g005(.A1(KEYINPUT76), .A2(G107), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n190), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT77), .ZN(new_n194));
  INV_X1    g008(.A(G107), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G104), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(G104), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(KEYINPUT3), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT77), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n190), .B(new_n199), .C1(new_n192), .C2(new_n191), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n194), .A2(new_n198), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G101), .ZN(new_n202));
  XOR2_X1   g016(.A(KEYINPUT78), .B(G101), .Z(new_n203));
  NAND4_X1  g017(.A1(new_n194), .A2(new_n203), .A3(new_n198), .A4(new_n200), .ZN(new_n204));
  AND2_X1   g018(.A1(new_n204), .A2(KEYINPUT79), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(KEYINPUT79), .ZN(new_n206));
  OAI211_X1 g020(.A(KEYINPUT4), .B(new_n202), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  OR2_X1    g021(.A1(new_n202), .A2(KEYINPUT4), .ZN(new_n208));
  XNOR2_X1  g022(.A(G116), .B(G119), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT2), .B(G113), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n211), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n209), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n207), .A2(new_n208), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT76), .B(G107), .ZN(new_n217));
  OR3_X1    g031(.A1(new_n217), .A2(KEYINPUT80), .A3(G104), .ZN(new_n218));
  OAI211_X1 g032(.A(KEYINPUT80), .B(new_n196), .C1(new_n217), .C2(G104), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(G101), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n194), .A2(new_n200), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT79), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n222), .A2(new_n223), .A3(new_n203), .A4(new_n198), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n204), .A2(KEYINPUT79), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n221), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT5), .ZN(new_n227));
  INV_X1    g041(.A(G119), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(G116), .ZN(new_n229));
  OAI211_X1 g043(.A(G113), .B(new_n229), .C1(new_n210), .C2(new_n227), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n226), .A2(new_n214), .A3(new_n230), .ZN(new_n231));
  XOR2_X1   g045(.A(G110), .B(G122), .Z(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n216), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT83), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n216), .A2(new_n231), .A3(KEYINPUT83), .A4(new_n233), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n233), .B1(new_n216), .B2(new_n231), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT6), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G143), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G146), .ZN(new_n244));
  INV_X1    g058(.A(G146), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G143), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n244), .A2(new_n246), .A3(G128), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT64), .B1(new_n243), .B2(G146), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT64), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(new_n245), .A3(G143), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(new_n250), .A3(new_n244), .ZN(new_n251));
  XOR2_X1   g065(.A(KEYINPUT0), .B(G128), .Z(new_n252));
  AOI22_X1  g066(.A1(KEYINPUT0), .A2(new_n247), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G125), .ZN(new_n254));
  OR2_X1    g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OR2_X1    g069(.A1(new_n255), .A2(KEYINPUT84), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT1), .B1(new_n243), .B2(G146), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G128), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n251), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT1), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n244), .A2(new_n246), .A3(new_n260), .A4(G128), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n254), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n255), .A2(KEYINPUT84), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n256), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G224), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(G953), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n266), .B(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n239), .A2(new_n240), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n242), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n230), .A2(new_n214), .ZN(new_n272));
  XOR2_X1   g086(.A(new_n226), .B(new_n272), .Z(new_n273));
  XOR2_X1   g087(.A(new_n232), .B(KEYINPUT8), .Z(new_n274));
  AOI22_X1  g088(.A1(new_n236), .A2(new_n237), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n268), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n255), .A2(new_n264), .B1(KEYINPUT7), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n266), .B1(KEYINPUT85), .B2(new_n268), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT7), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT85), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n279), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n277), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(G902), .B1(new_n275), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n271), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(G210), .B1(G237), .B2(G902), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n285), .B(KEYINPUT86), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n271), .A2(new_n283), .A3(new_n285), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n188), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(G128), .B(G143), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT13), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n243), .A2(G128), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n292), .B(G134), .C1(KEYINPUT13), .C2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G134), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G122), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G116), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n298), .B(KEYINPUT91), .ZN(new_n299));
  OR2_X1    g113(.A1(new_n297), .A2(G116), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n217), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n217), .B1(new_n299), .B2(new_n300), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n294), .B(new_n296), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n299), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n300), .B(KEYINPUT14), .ZN(new_n306));
  OAI21_X1  g120(.A(G107), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n291), .B(new_n295), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n301), .A3(new_n308), .ZN(new_n309));
  XOR2_X1   g123(.A(KEYINPUT9), .B(G234), .Z(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G217), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n311), .A2(new_n312), .A3(G953), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n304), .A2(new_n309), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n313), .B1(new_n304), .B2(new_n309), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G902), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G478), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(KEYINPUT15), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n316), .B(new_n317), .C1(KEYINPUT15), .C2(new_n319), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT92), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n323), .B(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(G125), .B(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n245), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT72), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G125), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G140), .ZN(new_n330));
  INV_X1    g144(.A(G140), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n331), .A3(G125), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n327), .B1(new_n333), .B2(new_n245), .ZN(new_n334));
  NOR2_X1   g148(.A1(G237), .A2(G953), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G214), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(KEYINPUT87), .A3(new_n243), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n243), .A2(KEYINPUT87), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(G214), .A3(new_n335), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT18), .ZN(new_n340));
  INV_X1    g154(.A(G131), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n337), .B(new_n339), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n337), .A2(new_n339), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G131), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n334), .B(new_n342), .C1(new_n344), .C2(new_n340), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n333), .A2(KEYINPUT19), .ZN(new_n346));
  OR2_X1    g160(.A1(new_n326), .A2(KEYINPUT19), .ZN(new_n347));
  AOI21_X1  g161(.A(G146), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n330), .A2(new_n332), .A3(KEYINPUT16), .ZN(new_n349));
  OR3_X1    g163(.A1(new_n254), .A2(KEYINPUT16), .A3(G140), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(G146), .A3(new_n350), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n337), .A2(new_n341), .A3(new_n339), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n341), .B1(new_n337), .B2(new_n339), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n345), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(G113), .B(G122), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(new_n189), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT17), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n337), .A2(new_n341), .A3(new_n339), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n344), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n349), .A2(new_n350), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n245), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n353), .A2(KEYINPUT17), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n362), .A2(new_n351), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n357), .B(KEYINPUT88), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n345), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n359), .A2(new_n368), .ZN(new_n369));
  NOR3_X1   g183(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(G475), .A2(G902), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n359), .A2(new_n368), .A3(KEYINPUT89), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT89), .B1(new_n359), .B2(new_n368), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n371), .B1(new_n375), .B2(KEYINPUT20), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n366), .A2(new_n345), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n368), .B1(new_n377), .B2(new_n357), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n317), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G475), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT90), .B1(new_n376), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT90), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT20), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT89), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n369), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n359), .A2(new_n368), .A3(KEYINPUT89), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n384), .B1(new_n388), .B2(new_n372), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n383), .B(new_n380), .C1(new_n389), .C2(new_n371), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n382), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(KEYINPUT93), .B(G952), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n392), .A2(G953), .ZN(new_n393));
  NAND2_X1  g207(.A1(G234), .A2(G237), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(KEYINPUT21), .B(G898), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(KEYINPUT94), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n394), .A2(G902), .A3(G953), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n396), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n325), .A2(new_n391), .A3(new_n400), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n290), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT11), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(new_n295), .B2(G137), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n295), .A2(G137), .ZN(new_n405));
  INV_X1    g219(.A(G137), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(KEYINPUT11), .A3(G134), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G131), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n404), .A2(new_n407), .A3(new_n341), .A4(new_n405), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n253), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n406), .A2(G134), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n295), .A2(G137), .ZN(new_n414));
  OAI21_X1  g228(.A(G131), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n262), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n215), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n412), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n418), .B1(new_n412), .B2(new_n417), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT28), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n412), .A2(new_n417), .A3(new_n418), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT28), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n335), .A2(G210), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(G101), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n421), .A2(KEYINPUT29), .A3(new_n424), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n317), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT67), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(KEYINPUT67), .A3(new_n317), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT66), .B1(new_n421), .B2(new_n424), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT66), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n412), .A2(new_n417), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n215), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n422), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n435), .B1(new_n438), .B2(KEYINPUT28), .ZN(new_n439));
  INV_X1    g253(.A(new_n428), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n434), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT29), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT30), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n412), .A2(new_n417), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n443), .B1(new_n412), .B2(new_n417), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n215), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n446), .A2(new_n422), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n442), .B1(new_n447), .B2(new_n428), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n432), .B(new_n433), .C1(new_n441), .C2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G472), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n446), .A2(new_n422), .A3(new_n428), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT31), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT65), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n440), .B1(new_n434), .B2(new_n439), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT31), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n447), .A2(new_n456), .A3(new_n428), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n451), .A2(KEYINPUT65), .A3(KEYINPUT31), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n454), .A2(new_n455), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT32), .ZN(new_n460));
  NOR2_X1   g274(.A1(G472), .A2(G902), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n460), .B1(new_n459), .B2(new_n461), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n450), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT68), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT68), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n466), .B(new_n450), .C1(new_n462), .C2(new_n463), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT22), .B(G137), .ZN(new_n468));
  INV_X1    g282(.A(G953), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(G221), .A3(G234), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n468), .B(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G128), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G119), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT23), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n473), .A2(KEYINPUT23), .A3(G119), .ZN(new_n477));
  INV_X1    g291(.A(G110), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n228), .A2(G128), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n476), .A2(new_n477), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT73), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n480), .B(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n474), .A2(new_n479), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT69), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT69), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n474), .A2(new_n479), .A3(new_n485), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT24), .B(G110), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT70), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n351), .B(new_n327), .C1(new_n482), .C2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT70), .ZN(new_n492));
  OR2_X1    g306(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n488), .A2(new_n492), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n493), .A2(new_n486), .A3(new_n484), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT71), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n364), .A2(new_n351), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n476), .A2(new_n479), .A3(new_n477), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G110), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT71), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n487), .A2(new_n489), .A3(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n496), .A2(new_n497), .A3(new_n499), .A4(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n491), .A2(new_n502), .A3(KEYINPUT74), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT74), .B1(new_n491), .B2(new_n502), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n472), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n491), .A2(new_n502), .A3(new_n471), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT25), .B1(new_n508), .B2(G902), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n312), .B1(G234), .B2(new_n317), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT25), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n506), .A2(new_n511), .A3(new_n317), .A4(new_n507), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n510), .A2(G902), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n506), .A2(new_n507), .A3(new_n514), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n465), .A2(new_n467), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(G221), .B1(new_n311), .B2(G902), .ZN(new_n518));
  XOR2_X1   g332(.A(new_n518), .B(KEYINPUT75), .Z(new_n519));
  NAND3_X1  g333(.A1(new_n207), .A2(new_n253), .A3(new_n208), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n244), .A2(new_n246), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n258), .A2(new_n521), .ZN(new_n522));
  OR2_X1    g336(.A1(new_n522), .A2(KEYINPUT81), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(KEYINPUT81), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n524), .A3(new_n261), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n220), .B(new_n525), .C1(new_n205), .C2(new_n206), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT10), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n411), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n263), .A2(new_n527), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n226), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n520), .A2(new_n528), .A3(new_n529), .A4(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n526), .B1(new_n226), .B2(new_n262), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n533), .A2(KEYINPUT12), .A3(new_n411), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT12), .B1(new_n533), .B2(new_n411), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g350(.A(G110), .B(G140), .ZN(new_n537));
  INV_X1    g351(.A(G227), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(G953), .ZN(new_n539));
  XOR2_X1   g353(.A(new_n537), .B(new_n539), .Z(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n532), .A2(new_n540), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n526), .A2(new_n527), .B1(new_n226), .B2(new_n530), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n529), .B1(new_n543), .B2(new_n520), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n536), .A2(new_n541), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(G469), .B1(new_n546), .B2(G902), .ZN(new_n547));
  INV_X1    g361(.A(new_n532), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n541), .B1(new_n548), .B2(new_n544), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n532), .B(new_n540), .C1(new_n534), .C2(new_n535), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G469), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n552), .A3(new_n317), .ZN(new_n553));
  AOI211_X1 g367(.A(KEYINPUT82), .B(new_n519), .C1(new_n547), .C2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT82), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n536), .A2(new_n541), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n542), .A2(new_n545), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(G469), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(G469), .A2(G902), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n553), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n519), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n555), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n554), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n402), .A2(new_n517), .A3(new_n563), .ZN(new_n564));
  XOR2_X1   g378(.A(new_n564), .B(new_n203), .Z(G3));
  INV_X1    g379(.A(G472), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(new_n459), .B2(new_n317), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n459), .A2(new_n461), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n554), .A2(new_n562), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n516), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(KEYINPUT95), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n271), .A2(new_n283), .A3(new_n285), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n285), .B1(new_n271), .B2(new_n283), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n187), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT33), .B1(new_n314), .B2(KEYINPUT96), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  OR2_X1    g392(.A1(new_n578), .A2(new_n316), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n316), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(G478), .A3(new_n317), .ZN(new_n582));
  INV_X1    g396(.A(new_n318), .ZN(new_n583));
  XNOR2_X1  g397(.A(KEYINPUT97), .B(G478), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n391), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n576), .A2(new_n400), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n573), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(new_n189), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(G6));
  OAI21_X1  g405(.A(new_n370), .B1(new_n373), .B2(new_n374), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT100), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n375), .A2(KEYINPUT99), .A3(KEYINPUT20), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT99), .B1(new_n375), .B2(KEYINPUT20), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT101), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n594), .B(KEYINPUT101), .C1(new_n595), .C2(new_n596), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n599), .A2(new_n380), .A3(new_n325), .A4(new_n600), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n601), .A2(new_n576), .A3(new_n400), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n573), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT35), .B(G107), .Z(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G9));
  NAND2_X1  g419(.A1(new_n560), .A2(new_n561), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(KEYINPUT82), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n519), .B1(new_n547), .B2(new_n553), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n555), .ZN(new_n609));
  INV_X1    g423(.A(new_n505), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n472), .A2(KEYINPUT36), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n610), .A2(new_n503), .A3(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n611), .B1(new_n504), .B2(new_n505), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n514), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT102), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n615), .A2(KEYINPUT102), .A3(new_n514), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n513), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(KEYINPUT103), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT103), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n513), .A2(new_n622), .A3(new_n618), .A4(new_n619), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n607), .A2(new_n609), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n570), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(new_n402), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT37), .B(G110), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G12));
  NAND3_X1  g443(.A1(new_n607), .A2(new_n609), .A3(new_n624), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n465), .A2(new_n467), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n630), .A2(new_n631), .A3(new_n576), .ZN(new_n632));
  INV_X1    g446(.A(G900), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n399), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n395), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n601), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G128), .ZN(G30));
  XNOR2_X1  g452(.A(new_n635), .B(KEYINPUT39), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n554), .A2(new_n562), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT40), .ZN(new_n641));
  INV_X1    g455(.A(new_n620), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n288), .A2(new_n289), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT38), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n569), .A2(KEYINPUT32), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n447), .A2(new_n440), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n317), .B1(new_n438), .B2(new_n428), .ZN(new_n649));
  OAI21_X1  g463(.A(G472), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n325), .A2(new_n391), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n652), .A2(new_n188), .A3(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n641), .A2(new_n642), .A3(new_n644), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G143), .ZN(G45));
  INV_X1    g470(.A(new_n635), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n585), .A2(new_n391), .A3(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n632), .A2(KEYINPUT104), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n466), .B1(new_n647), .B2(new_n450), .ZN(new_n662));
  INV_X1    g476(.A(new_n467), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n285), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n284), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n188), .B1(new_n666), .B2(new_n289), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n563), .A2(new_n664), .A3(new_n667), .A4(new_n624), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n661), .B1(new_n668), .B2(new_n658), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n660), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G146), .ZN(G48));
  AOI21_X1  g485(.A(new_n552), .B1(new_n551), .B2(new_n317), .ZN(new_n672));
  AOI211_X1 g486(.A(G469), .B(G902), .C1(new_n549), .C2(new_n550), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n672), .A2(new_n673), .A3(new_n519), .ZN(new_n674));
  AND4_X1   g488(.A1(new_n465), .A2(new_n467), .A3(new_n516), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n587), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT41), .B(G113), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G15));
  NAND2_X1  g492(.A1(new_n602), .A2(new_n675), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G116), .ZN(G18));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n667), .A2(new_n401), .A3(new_n674), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n624), .A2(new_n465), .A3(new_n467), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n624), .A2(new_n465), .A3(new_n467), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n682), .A2(new_n686), .A3(KEYINPUT105), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(new_n228), .ZN(G21));
  AND2_X1   g503(.A1(new_n421), .A2(new_n424), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n457), .B(new_n452), .C1(new_n690), .C2(new_n428), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n691), .A2(new_n461), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n567), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n516), .A2(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n576), .A2(new_n694), .A3(new_n400), .ZN(new_n695));
  INV_X1    g509(.A(new_n674), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n653), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G122), .ZN(G24));
  AND2_X1   g513(.A1(new_n693), .A2(new_n620), .ZN(new_n700));
  AND4_X1   g514(.A1(new_n667), .A2(new_n659), .A3(new_n700), .A4(new_n674), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n254), .ZN(G27));
  NAND3_X1  g516(.A1(new_n288), .A2(new_n187), .A3(new_n289), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n703), .A2(new_n586), .A3(new_n635), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n464), .A2(new_n516), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n704), .A2(KEYINPUT42), .A3(new_n608), .A4(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n465), .A2(new_n467), .A3(new_n516), .ZN(new_n707));
  NOR4_X1   g521(.A1(new_n707), .A2(new_n606), .A3(new_n658), .A4(new_n703), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n706), .B1(new_n708), .B2(KEYINPUT42), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G131), .ZN(G33));
  INV_X1    g524(.A(new_n703), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n517), .A2(new_n636), .A3(new_n608), .A4(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n707), .A2(new_n606), .A3(new_n703), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(KEYINPUT106), .A3(new_n636), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G134), .ZN(G36));
  INV_X1    g532(.A(new_n391), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT43), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n719), .A2(new_n585), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n391), .B(KEYINPUT109), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n585), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n721), .B1(new_n723), .B2(KEYINPUT43), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT110), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n570), .A2(new_n620), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT111), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n726), .A2(KEYINPUT112), .A3(KEYINPUT44), .A4(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n724), .A2(new_n725), .ZN(new_n730));
  AOI211_X1 g544(.A(KEYINPUT110), .B(new_n721), .C1(new_n723), .C2(KEYINPUT43), .ZN(new_n731));
  OAI211_X1 g545(.A(KEYINPUT44), .B(new_n728), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n729), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n726), .A2(new_n728), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n703), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n739));
  OAI21_X1  g553(.A(G469), .B1(new_n546), .B2(KEYINPUT45), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT107), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n546), .A2(KEYINPUT45), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n559), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT46), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n739), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n743), .A2(KEYINPUT108), .A3(KEYINPUT46), .A4(new_n559), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n746), .A2(new_n747), .A3(new_n553), .A4(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n639), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n561), .A3(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n735), .A2(new_n738), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G137), .ZN(G39));
  NAND2_X1  g568(.A1(new_n711), .A2(new_n657), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n755), .A2(new_n516), .A3(new_n586), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n749), .A2(KEYINPUT47), .A3(new_n561), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT47), .B1(new_n749), .B2(new_n561), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n631), .B(new_n756), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G140), .ZN(G42));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n762));
  AOI22_X1  g576(.A1(new_n587), .A2(new_n675), .B1(new_n695), .B2(new_n697), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n763), .B(new_n679), .C1(new_n685), .C2(new_n687), .ZN(new_n764));
  INV_X1    g578(.A(new_n400), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n286), .B1(new_n271), .B2(new_n283), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n187), .B(new_n765), .C1(new_n574), .C2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n586), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n571), .A2(new_n516), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n771));
  INV_X1    g585(.A(new_n323), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n391), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n771), .B1(new_n767), .B2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n290), .A2(KEYINPUT113), .A3(new_n765), .A4(new_n773), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n571), .A2(new_n775), .A3(new_n776), .A4(new_n516), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n627), .A2(new_n770), .A3(new_n777), .A4(new_n564), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n764), .A2(new_n778), .ZN(new_n779));
  AND4_X1   g593(.A1(new_n380), .A2(new_n599), .A3(new_n772), .A4(new_n600), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n625), .A2(new_n664), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n769), .A2(new_n608), .A3(new_n700), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n755), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n715), .A2(new_n659), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT42), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI22_X1  g601(.A1(new_n787), .A2(new_n706), .B1(new_n714), .B2(new_n716), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n779), .A2(new_n784), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT114), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n701), .B1(new_n632), .B2(new_n636), .ZN(new_n791));
  INV_X1    g605(.A(new_n653), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n667), .A2(new_n642), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n651), .A2(new_n608), .A3(new_n657), .ZN(new_n794));
  OR3_X1    g608(.A1(new_n793), .A2(KEYINPUT115), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(KEYINPUT115), .B1(new_n793), .B2(new_n794), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT104), .B1(new_n632), .B2(new_n659), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n668), .A2(new_n661), .A3(new_n658), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n791), .B(new_n797), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n670), .A2(KEYINPUT52), .A3(new_n791), .A4(new_n797), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n779), .A2(new_n788), .A3(new_n805), .A4(new_n784), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n790), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n762), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n717), .A2(new_n709), .ZN(new_n812));
  NOR4_X1   g626(.A1(new_n812), .A2(new_n764), .A3(new_n778), .A4(new_n783), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n804), .A2(KEYINPUT53), .A3(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n810), .A2(new_n762), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n724), .A2(new_n396), .ZN(new_n817));
  INV_X1    g631(.A(new_n694), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n188), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n644), .A2(new_n696), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  OR3_X1    g636(.A1(new_n820), .A2(KEYINPUT50), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n696), .A2(new_n703), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n817), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n700), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT50), .B1(new_n820), .B2(new_n822), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n823), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n824), .A2(new_n516), .A3(new_n396), .A4(new_n652), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n829), .A2(new_n391), .A3(new_n585), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n759), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n672), .A2(new_n673), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n519), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n832), .A2(new_n757), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(new_n711), .A3(new_n819), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT51), .B1(new_n831), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n825), .A2(new_n705), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n838), .A2(KEYINPUT48), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(KEYINPUT48), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n819), .A2(new_n667), .A3(new_n674), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n839), .A2(new_n393), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n837), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n819), .A2(new_n711), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n835), .B(KEYINPUT116), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n831), .B(KEYINPUT51), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n816), .A2(new_n843), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n829), .A2(new_n586), .ZN(new_n848));
  OAI22_X1  g662(.A1(new_n847), .A2(new_n848), .B1(G952), .B2(G953), .ZN(new_n849));
  XOR2_X1   g663(.A(new_n833), .B(KEYINPUT49), .Z(new_n850));
  NAND4_X1  g664(.A1(new_n652), .A2(new_n561), .A3(new_n516), .A4(new_n187), .ZN(new_n851));
  OR4_X1    g665(.A1(new_n644), .A2(new_n850), .A3(new_n851), .A4(new_n723), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n849), .A2(new_n852), .ZN(G75));
  NOR2_X1   g667(.A1(new_n469), .A2(G952), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT119), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n804), .A2(KEYINPUT53), .A3(new_n813), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n857), .B1(new_n808), .B2(new_n807), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n317), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT56), .B1(new_n859), .B2(G210), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n242), .A2(new_n270), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(new_n269), .ZN(new_n862));
  XOR2_X1   g676(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n863));
  XNOR2_X1  g677(.A(new_n862), .B(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n856), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT118), .B1(new_n858), .B2(new_n317), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n810), .A2(new_n814), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n867), .A2(new_n868), .A3(G902), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n287), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n864), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n865), .B1(new_n870), .B2(new_n872), .ZN(G51));
  XOR2_X1   g687(.A(new_n743), .B(KEYINPUT120), .Z(new_n874));
  NAND3_X1  g688(.A1(new_n866), .A2(new_n869), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT121), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n762), .B1(new_n810), .B2(new_n814), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n815), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n559), .B(KEYINPUT57), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n551), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n866), .A2(new_n869), .A3(new_n881), .A4(new_n874), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n876), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n854), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(G54));
  NAND4_X1  g699(.A1(new_n866), .A2(new_n869), .A3(KEYINPUT58), .A4(G475), .ZN(new_n886));
  INV_X1    g700(.A(new_n388), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n888), .A2(new_n889), .A3(new_n854), .ZN(G60));
  NAND2_X1  g704(.A1(G478), .A2(G902), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT59), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n581), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n856), .B1(new_n878), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n892), .B1(new_n811), .B2(new_n815), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(new_n579), .A3(new_n580), .ZN(new_n898));
  OAI211_X1 g712(.A(KEYINPUT122), .B(new_n856), .C1(new_n878), .C2(new_n893), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(G63));
  NAND2_X1  g714(.A1(G217), .A2(G902), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT60), .Z(new_n902));
  NAND2_X1  g716(.A1(new_n867), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n508), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n867), .A2(new_n615), .A3(new_n902), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n856), .A3(new_n905), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g721(.A(G953), .B1(new_n398), .B2(new_n267), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n908), .B1(new_n779), .B2(G953), .ZN(new_n909));
  INV_X1    g723(.A(G898), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n861), .B1(new_n910), .B2(G953), .ZN(new_n911));
  XNOR2_X1  g725(.A(KEYINPUT123), .B(KEYINPUT124), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n909), .B(new_n913), .ZN(G69));
  NOR2_X1   g728(.A1(new_n444), .A2(new_n445), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n346), .A2(new_n347), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n915), .B(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT125), .ZN(new_n918));
  AOI21_X1  g732(.A(G900), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n917), .B(KEYINPUT125), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(new_n538), .ZN(new_n921));
  AOI211_X1 g735(.A(new_n469), .B(new_n919), .C1(new_n921), .C2(G900), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n664), .B1(new_n832), .B2(new_n757), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n751), .B1(new_n729), .B2(new_n734), .ZN(new_n924));
  AOI22_X1  g738(.A1(new_n923), .A2(new_n756), .B1(new_n924), .B2(new_n738), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n752), .A2(new_n667), .A3(new_n792), .A4(new_n705), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n670), .A2(new_n791), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n928), .A2(new_n788), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n925), .A2(new_n926), .A3(new_n927), .A4(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n753), .A2(new_n760), .A3(new_n927), .A4(new_n929), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT126), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n920), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n928), .A2(new_n655), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n935), .B(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n774), .A2(new_n586), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n640), .A2(new_n517), .A3(new_n711), .A4(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n937), .A2(new_n925), .A3(new_n939), .ZN(new_n940));
  OAI22_X1  g754(.A1(new_n933), .A2(new_n917), .B1(new_n934), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n922), .B1(new_n941), .B2(new_n469), .ZN(G72));
  NAND3_X1  g756(.A1(new_n930), .A2(new_n932), .A3(new_n779), .ZN(new_n943));
  NAND2_X1  g757(.A1(G472), .A2(G902), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT63), .Z(new_n945));
  NAND2_X1  g759(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n447), .A2(new_n440), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n779), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n945), .B1(new_n940), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n854), .B1(new_n951), .B2(new_n648), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n809), .A2(new_n810), .ZN(new_n953));
  INV_X1    g767(.A(new_n648), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n953), .A2(new_n954), .A3(new_n945), .A4(new_n947), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n949), .A2(new_n952), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(KEYINPUT127), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n949), .A2(new_n958), .A3(new_n952), .A4(new_n955), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(G57));
endmodule


