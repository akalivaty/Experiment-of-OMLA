//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 0 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1267,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n209), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT65), .Z(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n211), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n214), .B(new_n219), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XOR2_X1   g0037(.A(G50), .B(G58), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  NAND3_X1  g0043(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(new_n217), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT8), .B(G58), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G20), .A2(G33), .ZN(new_n249));
  AOI22_X1  g0049(.A1(new_n248), .A2(new_n249), .B1(G20), .B2(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT15), .B(G87), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n209), .A2(G33), .ZN(new_n252));
  OR2_X1    g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n246), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n245), .B1(new_n208), .B2(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G77), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n256), .B1(G77), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n263), .A2(G232), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G107), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n269), .B1(new_n270), .B2(new_n268), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n272), .B1(new_n266), .B2(new_n267), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT69), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT69), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n271), .B1(new_n278), .B2(G238), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  OAI211_X1 g0080(.A(G1), .B(G13), .C1(new_n265), .C2(new_n280), .ZN(new_n281));
  OR2_X1    g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n208), .A2(G274), .ZN(new_n283));
  AND2_X1   g0083(.A1(KEYINPUT66), .A2(G41), .ZN(new_n284));
  NOR2_X1   g0084(.A1(KEYINPUT66), .A2(G41), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G45), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n283), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT67), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G41), .A2(G45), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n290), .B1(new_n291), .B2(G1), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n208), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n289), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n288), .B1(new_n294), .B2(G244), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n282), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G169), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n259), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G179), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n282), .A2(new_n299), .A3(new_n295), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g0101(.A(KEYINPUT74), .B(G200), .Z(new_n302));
  AOI21_X1  g0102(.A(new_n302), .B1(new_n282), .B2(new_n295), .ZN(new_n303));
  OAI211_X1 g0103(.A(G190), .B(new_n295), .C1(new_n279), .C2(new_n281), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n259), .ZN(new_n305));
  INV_X1    g0105(.A(G223), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(new_n275), .B2(new_n277), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT68), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n272), .ZN(new_n310));
  AND2_X1   g0110(.A1(KEYINPUT3), .A2(G33), .ZN(new_n311));
  NOR2_X1   g0111(.A1(KEYINPUT3), .A2(G33), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n310), .B(new_n260), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n311), .A2(new_n312), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n314), .A2(G222), .B1(G77), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n308), .A2(KEYINPUT70), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT70), .ZN(new_n318));
  INV_X1    g0118(.A(new_n316), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n318), .B1(new_n319), .B2(new_n307), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n317), .A2(new_n289), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n288), .B1(new_n294), .B2(G226), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT73), .B1(new_n323), .B2(G169), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n299), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n247), .A2(KEYINPUT71), .ZN(new_n327));
  INV_X1    g0127(.A(G58), .ZN(new_n328));
  OR3_X1    g0128(.A1(new_n328), .A2(KEYINPUT71), .A3(KEYINPUT8), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n327), .A2(new_n209), .A3(G33), .A4(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n249), .A2(G150), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT72), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT72), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n330), .A2(new_n335), .A3(new_n331), .ZN(new_n336));
  INV_X1    g0136(.A(new_n203), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n336), .B1(new_n209), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n245), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n257), .A2(G50), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n255), .B2(G50), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT73), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n342), .B1(new_n325), .B2(new_n343), .ZN(new_n344));
  OAI221_X1 g0144(.A(new_n301), .B1(new_n303), .B2(new_n305), .C1(new_n326), .C2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n341), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n333), .B(new_n336), .C1(new_n209), .C2(new_n337), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n346), .B1(new_n347), .B2(new_n245), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT75), .B1(new_n348), .B2(KEYINPUT9), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT75), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT9), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n342), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n348), .A2(KEYINPUT9), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n321), .A2(G190), .A3(new_n322), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n354), .B(new_n355), .C1(new_n323), .C2(new_n302), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n353), .A2(new_n356), .A3(KEYINPUT10), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT10), .ZN(new_n358));
  INV_X1    g0158(.A(new_n355), .ZN(new_n359));
  AOI211_X1 g0159(.A(new_n351), .B(new_n346), .C1(new_n347), .C2(new_n245), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n302), .B1(new_n321), .B2(new_n322), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n349), .A2(new_n352), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n358), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n357), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G68), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT7), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n268), .B2(G20), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n315), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n328), .A2(new_n366), .ZN(new_n371));
  OAI21_X1  g0171(.A(G20), .B1(new_n371), .B2(new_n202), .ZN(new_n372));
  INV_X1    g0172(.A(G159), .ZN(new_n373));
  INV_X1    g0173(.A(new_n249), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT77), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n376), .A2(KEYINPUT16), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n246), .B1(new_n376), .B2(KEYINPUT16), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n327), .A2(new_n329), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n257), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n379), .B2(new_n255), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT78), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT78), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n380), .B(new_n383), .C1(new_n379), .C2(new_n255), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n377), .A2(new_n378), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G200), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G87), .ZN(new_n387));
  INV_X1    g0187(.A(G226), .ZN(new_n388));
  OAI221_X1 g0188(.A(new_n387), .B1(new_n313), .B2(new_n306), .C1(new_n274), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n289), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n288), .B1(new_n294), .B2(G232), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n386), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n390), .A2(new_n391), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n392), .B1(G190), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n385), .A2(new_n394), .ZN(new_n395));
  XOR2_X1   g0195(.A(KEYINPUT80), .B(KEYINPUT17), .Z(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT81), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(KEYINPUT17), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT81), .ZN(new_n399));
  INV_X1    g0199(.A(new_n396), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n385), .A2(new_n394), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n397), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT79), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n390), .A2(new_n299), .A3(new_n391), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n393), .B2(G169), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n385), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT18), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n385), .B2(new_n405), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n403), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n409), .A2(new_n403), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n402), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI211_X1 g0212(.A(G232), .B(G1698), .C1(new_n311), .C2(new_n312), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G33), .A2(G97), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n413), .B(new_n414), .C1(new_n313), .C2(new_n388), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n289), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n288), .B1(new_n294), .B2(G238), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT13), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT76), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT13), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n416), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n419), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n416), .A2(new_n417), .A3(KEYINPUT76), .A4(new_n421), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(G169), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT14), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT14), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n423), .A2(new_n427), .A3(G169), .A4(new_n424), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n419), .A2(G179), .A3(new_n422), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n426), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n255), .A2(G68), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT12), .ZN(new_n432));
  INV_X1    g0232(.A(new_n257), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n432), .B1(new_n433), .B2(new_n366), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n257), .A2(KEYINPUT12), .A3(G68), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n431), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT11), .ZN(new_n437));
  INV_X1    g0237(.A(G50), .ZN(new_n438));
  OAI22_X1  g0238(.A1(new_n374), .A2(new_n438), .B1(new_n209), .B2(G68), .ZN(new_n439));
  INV_X1    g0239(.A(G77), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n252), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n245), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n436), .B1(new_n437), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n437), .B2(new_n442), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n430), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(G190), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n446), .B1(new_n418), .B2(KEYINPUT13), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n444), .B1(new_n422), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n423), .A2(G200), .A3(new_n424), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n445), .A2(new_n451), .ZN(new_n452));
  NOR4_X1   g0252(.A1(new_n345), .A2(new_n365), .A3(new_n412), .A4(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  XOR2_X1   g0254(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n455));
  INV_X1    g0255(.A(G244), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n313), .B2(new_n456), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n273), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n263), .A2(new_n268), .A3(KEYINPUT4), .A4(G244), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n289), .ZN(new_n461));
  OR2_X1    g0261(.A1(KEYINPUT66), .A2(G41), .ZN(new_n462));
  NAND2_X1  g0262(.A1(KEYINPUT66), .A2(G41), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT5), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT5), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n208), .B(G45), .C1(new_n465), .C2(G41), .ZN(new_n466));
  OAI211_X1 g0266(.A(G257), .B(new_n281), .C1(new_n464), .C2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n466), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n465), .B1(new_n284), .B2(new_n285), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n468), .A2(new_n469), .A3(G274), .A4(new_n281), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n461), .A2(G190), .A3(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n257), .A2(G97), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n208), .A2(G33), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n257), .A2(new_n475), .A3(new_n217), .A4(new_n244), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n474), .B1(new_n477), .B2(G97), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT7), .B1(new_n315), .B2(new_n209), .ZN(new_n480));
  NOR4_X1   g0280(.A1(new_n311), .A2(new_n312), .A3(new_n367), .A4(G20), .ZN(new_n481));
  OAI21_X1  g0281(.A(G107), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT6), .ZN(new_n483));
  AND2_X1   g0283(.A1(G97), .A2(G107), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(new_n205), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n270), .A2(KEYINPUT6), .A3(G97), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n487), .A2(G20), .B1(G77), .B2(new_n249), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n482), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n479), .B1(new_n489), .B2(new_n245), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n473), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n471), .B1(new_n460), .B2(new_n289), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(new_n386), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT83), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n461), .A2(new_n472), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G200), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT83), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n496), .A2(new_n497), .A3(new_n490), .A4(new_n473), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n492), .A2(G179), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n297), .B2(new_n492), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n489), .A2(new_n245), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n502), .A2(KEYINPUT84), .A3(new_n478), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT84), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n246), .B1(new_n482), .B2(new_n488), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n504), .B1(new_n505), .B2(new_n479), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n499), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT85), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n494), .A2(new_n498), .B1(new_n501), .B2(new_n507), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT85), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n268), .A2(new_n209), .A3(G68), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT19), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n209), .B1(new_n414), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(G87), .B2(new_n206), .ZN(new_n517));
  INV_X1    g0317(.A(G97), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n515), .B1(new_n252), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n514), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n520), .A2(new_n245), .B1(new_n433), .B2(new_n251), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n477), .A2(G87), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(G116), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n265), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n456), .A2(new_n272), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(new_n312), .B2(new_n311), .ZN(new_n528));
  INV_X1    g0328(.A(G238), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n526), .B(new_n528), .C1(new_n313), .C2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n289), .ZN(new_n531));
  OR3_X1    g0331(.A1(new_n287), .A2(G1), .A3(G274), .ZN(new_n532));
  INV_X1    g0332(.A(G250), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n287), .B2(G1), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n281), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n302), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n523), .B(new_n538), .C1(new_n446), .C2(new_n536), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n521), .B1(new_n251), .B2(new_n476), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n536), .A2(new_n297), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n540), .B(new_n541), .C1(G179), .C2(new_n536), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n510), .A2(new_n513), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n268), .A2(new_n209), .A3(G87), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT22), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT22), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n268), .A2(new_n547), .A3(new_n209), .A4(G87), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT24), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT23), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n209), .B2(G107), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n270), .A2(KEYINPUT23), .A3(G20), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n552), .A2(new_n553), .B1(new_n525), .B2(new_n209), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n549), .A2(new_n550), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n550), .B1(new_n549), .B2(new_n554), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n245), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n433), .A2(KEYINPUT25), .A3(new_n270), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT25), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n257), .B2(G107), .ZN(new_n560));
  AOI22_X1  g0360(.A1(G107), .A2(new_n477), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(G257), .B(G1698), .C1(new_n311), .C2(new_n312), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G33), .A2(G294), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n563), .B(new_n564), .C1(new_n313), .C2(new_n533), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n289), .ZN(new_n566));
  OAI211_X1 g0366(.A(G264), .B(new_n281), .C1(new_n464), .C2(new_n466), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n566), .A2(new_n446), .A3(new_n470), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT88), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n566), .A2(KEYINPUT88), .A3(new_n567), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n470), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n386), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n562), .B1(new_n568), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n571), .A2(G179), .A3(new_n470), .A4(new_n572), .ZN(new_n576));
  INV_X1    g0376(.A(new_n470), .ZN(new_n577));
  OAI21_X1  g0377(.A(G169), .B1(new_n569), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n576), .A2(new_n578), .B1(new_n557), .B2(new_n561), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT21), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n257), .A2(new_n475), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT86), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(new_n246), .A4(G116), .ZN(new_n584));
  OAI21_X1  g0384(.A(KEYINPUT86), .B1(new_n476), .B2(new_n524), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n433), .A2(new_n524), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(G20), .B1(G33), .B2(G283), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(G33), .B2(new_n518), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT87), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n524), .A2(G20), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n245), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n591), .B1(new_n245), .B2(new_n592), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n590), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT20), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(KEYINPUT20), .B(new_n590), .C1(new_n594), .C2(new_n595), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n588), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(G257), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(new_n266), .B2(new_n267), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n602), .A2(new_n263), .B1(new_n315), .B2(G303), .ZN(new_n603));
  OAI211_X1 g0403(.A(G264), .B(G1698), .C1(new_n311), .C2(new_n312), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n281), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(G270), .B(new_n281), .C1(new_n464), .C2(new_n466), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n470), .ZN(new_n607));
  OAI21_X1  g0407(.A(G169), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n581), .B1(new_n600), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n584), .A2(new_n585), .B1(new_n524), .B2(new_n433), .ZN(new_n610));
  INV_X1    g0410(.A(new_n595), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n593), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT20), .B1(new_n612), .B2(new_n590), .ZN(new_n613));
  INV_X1    g0413(.A(new_n599), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n610), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n605), .A2(new_n607), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(G179), .A3(new_n616), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n606), .A2(new_n470), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n266), .A2(G303), .A3(new_n267), .ZN(new_n619));
  OAI21_X1  g0419(.A(G257), .B1(new_n311), .B2(new_n312), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n310), .A2(new_n260), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n604), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n289), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n297), .B1(new_n618), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n615), .A2(KEYINPUT21), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(G200), .B1(new_n605), .B2(new_n607), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n618), .A2(G190), .A3(new_n623), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n598), .A2(new_n599), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .A4(new_n610), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n609), .A2(new_n617), .A3(new_n625), .A4(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n580), .A2(new_n631), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n454), .A2(new_n544), .A3(new_n632), .ZN(G372));
  NOR2_X1   g0433(.A1(new_n326), .A2(new_n344), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n407), .A2(new_n409), .ZN(new_n635));
  INV_X1    g0435(.A(new_n301), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n451), .A2(new_n636), .B1(new_n444), .B2(new_n430), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n637), .A2(KEYINPUT90), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n402), .B1(new_n637), .B2(KEYINPUT90), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n635), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT91), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n357), .B2(new_n364), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT10), .B1(new_n353), .B2(new_n356), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n362), .A2(new_n358), .A3(new_n363), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n644), .A3(KEYINPUT91), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n634), .B1(new_n640), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n490), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n543), .A2(new_n501), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n542), .B1(new_n649), .B2(KEYINPUT26), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n539), .A2(new_n542), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n508), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT26), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n609), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n617), .A2(new_n625), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT89), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT89), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n579), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n566), .A2(KEYINPUT88), .A3(new_n567), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT88), .B1(new_n566), .B2(new_n567), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n662), .A2(new_n663), .A3(new_n577), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n568), .B1(new_n664), .B2(G200), .ZN(new_n665));
  INV_X1    g0465(.A(new_n562), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n511), .A2(new_n543), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n655), .B1(new_n661), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n647), .B1(new_n454), .B2(new_n670), .ZN(G369));
  NAND3_X1  g0471(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n580), .B1(new_n666), .B2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n579), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(new_n678), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT93), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n658), .A2(new_n677), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n579), .A2(new_n678), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n659), .A2(new_n660), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n600), .A2(new_n678), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n631), .A2(KEYINPUT92), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT92), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n689), .B1(new_n630), .B2(new_n691), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n688), .A2(new_n689), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n683), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n687), .A2(new_n697), .ZN(G399));
  INV_X1    g0498(.A(new_n212), .ZN(new_n699));
  INV_X1    g0499(.A(new_n286), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n215), .B2(new_n702), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n669), .A2(new_n678), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT29), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n652), .A2(new_n653), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n542), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(KEYINPUT26), .B2(new_n649), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n579), .A2(new_n656), .A3(new_n657), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n668), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n677), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT29), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n651), .B1(new_n509), .B2(KEYINPUT85), .ZN(new_n717));
  NOR4_X1   g0517(.A1(new_n575), .A2(new_n630), .A3(new_n579), .A4(new_n677), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(new_n718), .A3(new_n513), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT94), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT31), .ZN(new_n721));
  INV_X1    g0521(.A(new_n535), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n722), .B1(new_n530), .B2(new_n289), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(new_n618), .A3(G179), .A4(new_n623), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n724), .A2(new_n662), .A3(new_n663), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n492), .A2(KEYINPUT30), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n263), .A2(G238), .A3(new_n268), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n525), .B1(new_n268), .B2(new_n527), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n281), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n299), .B1(new_n730), .B2(new_n722), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n492), .A2(new_n616), .A3(new_n731), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n725), .A2(new_n727), .B1(new_n732), .B2(new_n573), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n623), .A2(G179), .A3(new_n470), .A4(new_n606), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(new_n536), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(new_n492), .A3(new_n571), .A4(new_n572), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI211_X1 g0538(.A(new_n721), .B(new_n678), .C1(new_n733), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n725), .A2(new_n727), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n732), .A2(new_n573), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n738), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(KEYINPUT31), .B1(new_n742), .B2(new_n677), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n720), .B1(new_n739), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n735), .A2(new_n571), .A3(new_n572), .ZN(new_n745));
  INV_X1    g0545(.A(new_n731), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n618), .A2(new_n623), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n495), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n745), .A2(new_n726), .B1(new_n664), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(KEYINPUT30), .B1(new_n725), .B2(new_n492), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n677), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n721), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n742), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n752), .A2(KEYINPUT94), .A3(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n719), .A2(new_n744), .A3(new_n754), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n709), .A2(new_n716), .B1(G330), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n706), .B1(new_n756), .B2(G1), .ZN(G364));
  AND2_X1   g0557(.A1(new_n209), .A2(G13), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n208), .B1(new_n758), .B2(G45), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n701), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n695), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n693), .A2(G330), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n693), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n212), .A2(new_n268), .ZN(new_n770));
  INV_X1    g0570(.A(G355), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n770), .A2(new_n771), .B1(G116), .B2(new_n212), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n699), .A2(new_n268), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(new_n287), .B2(new_n216), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n239), .A2(G45), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n217), .B1(G20), .B2(new_n297), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n767), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n761), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n209), .A2(G179), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n537), .A2(new_n446), .A3(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G107), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n209), .A2(new_n299), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT95), .Z(new_n787));
  NOR2_X1   g0587(.A1(G190), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n446), .A2(G200), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n785), .B1(new_n789), .B2(new_n440), .C1(new_n328), .C2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n786), .A2(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(G190), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n793), .A2(new_n446), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n795), .A2(new_n366), .B1(new_n797), .B2(new_n438), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n790), .A2(new_n299), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G20), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n782), .A2(new_n788), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n373), .ZN(new_n803));
  XOR2_X1   g0603(.A(KEYINPUT96), .B(KEYINPUT32), .Z(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n801), .A2(new_n518), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n537), .A2(G190), .A3(new_n782), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(G87), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n315), .B1(new_n803), .B2(new_n805), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR4_X1   g0611(.A1(new_n792), .A2(new_n798), .A3(new_n806), .A4(new_n811), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n812), .A2(KEYINPUT97), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(KEYINPUT97), .ZN(new_n814));
  INV_X1    g0614(.A(G329), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n315), .B1(new_n802), .B2(new_n815), .ZN(new_n816));
  XOR2_X1   g0616(.A(KEYINPUT33), .B(G317), .Z(new_n817));
  INV_X1    g0617(.A(G294), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n795), .A2(new_n817), .B1(new_n801), .B2(new_n818), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n816), .B(new_n819), .C1(G326), .C2(new_n796), .ZN(new_n820));
  INV_X1    g0620(.A(new_n789), .ZN(new_n821));
  INV_X1    g0621(.A(new_n791), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G311), .A2(new_n821), .B1(new_n822), .B2(G322), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G283), .A2(new_n784), .B1(new_n808), .B2(G303), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n820), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n813), .A2(new_n814), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n781), .B1(new_n826), .B2(new_n778), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n762), .A2(new_n764), .B1(new_n769), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G396));
  OAI22_X1  g0629(.A1(new_n303), .A2(new_n305), .B1(new_n259), .B2(new_n678), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n301), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n298), .A2(new_n300), .A3(new_n678), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n707), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n833), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n669), .A2(new_n678), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n755), .A2(G330), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n761), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n838), .B2(new_n837), .ZN(new_n840));
  INV_X1    g0640(.A(new_n761), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n778), .A2(new_n765), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n841), .B1(new_n440), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n778), .ZN(new_n844));
  INV_X1    g0644(.A(G303), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n315), .B1(new_n801), .B2(new_n518), .C1(new_n797), .C2(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n822), .A2(G294), .B1(G107), .B2(new_n808), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n524), .B2(new_n789), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n794), .A2(KEYINPUT98), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n794), .A2(KEYINPUT98), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n846), .B(new_n848), .C1(G283), .C2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n784), .A2(G87), .ZN(new_n854));
  INV_X1    g0654(.A(G311), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n854), .B1(new_n855), .B2(new_n802), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT99), .ZN(new_n857));
  AOI22_X1  g0657(.A1(G137), .A2(new_n796), .B1(new_n794), .B2(G150), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n789), .B2(new_n373), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(G143), .B2(new_n822), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT34), .Z(new_n861));
  NAND2_X1  g0661(.A1(new_n784), .A2(G68), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n438), .B2(new_n807), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n863), .A2(KEYINPUT100), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n863), .A2(KEYINPUT100), .ZN(new_n865));
  INV_X1    g0665(.A(G132), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n268), .B1(new_n802), .B2(new_n866), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n867), .A2(KEYINPUT101), .B1(new_n800), .B2(G58), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(KEYINPUT101), .B2(new_n867), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n864), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n853), .A2(new_n857), .B1(new_n861), .B2(new_n870), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n843), .B1(new_n844), .B2(new_n871), .C1(new_n835), .C2(new_n766), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n840), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(G384));
  INV_X1    g0674(.A(new_n385), .ZN(new_n875));
  INV_X1    g0675(.A(new_n675), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n412), .A2(new_n878), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n385), .A2(new_n405), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n877), .A2(new_n880), .A3(new_n395), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT103), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT37), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n877), .A2(new_n880), .A3(new_n884), .A4(new_n395), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n882), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n883), .B1(new_n882), .B2(new_n885), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n879), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT38), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n879), .B(KEYINPUT38), .C1(new_n886), .C2(new_n887), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n739), .A2(new_n743), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n631), .A2(new_n667), .A3(new_n680), .A4(new_n678), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n893), .B1(new_n544), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n444), .A2(new_n677), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n445), .A2(new_n451), .A3(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n444), .B(new_n677), .C1(new_n430), .C2(new_n450), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n833), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n892), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT40), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n882), .ZN(new_n905));
  INV_X1    g0705(.A(new_n885), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n877), .B1(new_n402), .B2(new_n635), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n889), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n891), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(new_n901), .A3(KEYINPUT40), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n904), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n453), .A2(new_n895), .ZN(new_n913));
  OAI21_X1  g0713(.A(G330), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n913), .B2(new_n912), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n910), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n890), .A2(KEYINPUT39), .A3(new_n891), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n445), .A2(new_n677), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n635), .A2(new_n876), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n897), .A2(new_n898), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n836), .B2(new_n832), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n921), .B1(new_n892), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n920), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n709), .A2(new_n453), .A3(new_n716), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n647), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n926), .B(new_n928), .Z(new_n929));
  OAI22_X1  g0729(.A1(new_n915), .A2(new_n929), .B1(new_n208), .B2(new_n758), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n929), .B2(new_n915), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n487), .A2(KEYINPUT35), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n487), .A2(KEYINPUT35), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n932), .A2(G116), .A3(new_n218), .A4(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT36), .Z(new_n935));
  NOR3_X1   g0735(.A1(new_n371), .A2(new_n215), .A3(new_n440), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT102), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n936), .A2(new_n937), .B1(new_n201), .B2(G68), .ZN(new_n939));
  AOI211_X1 g0739(.A(new_n208), .B(G13), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  OR3_X1    g0740(.A1(new_n931), .A2(new_n935), .A3(new_n940), .ZN(G367));
  OAI21_X1  g0741(.A(new_n511), .B1(new_n490), .B2(new_n678), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n501), .A2(new_n648), .A3(new_n677), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n696), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT104), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n945), .A2(new_n579), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n677), .B1(new_n949), .B2(new_n508), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n683), .A2(new_n684), .A3(new_n945), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n950), .B1(new_n951), .B2(KEYINPUT42), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(KEYINPUT42), .B2(new_n951), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n523), .A2(new_n678), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n543), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n542), .B2(new_n954), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n953), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n957), .B1(new_n953), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n948), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n946), .B(KEYINPUT104), .ZN(new_n962));
  OR3_X1    g0762(.A1(new_n959), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n701), .B(KEYINPUT41), .Z(new_n964));
  XOR2_X1   g0764(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n687), .B2(new_n945), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n685), .A2(new_n686), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n968), .A2(new_n944), .A3(new_n965), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n685), .A2(new_n686), .A3(new_n945), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT45), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n696), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n683), .A2(new_n684), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n685), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n694), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n974), .A2(new_n695), .A3(new_n685), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n976), .A2(new_n756), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT45), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n971), .B(new_n980), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n981), .A2(new_n697), .A3(new_n969), .A4(new_n967), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n973), .A2(new_n979), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n964), .B1(new_n983), .B2(new_n756), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n961), .B(new_n963), .C1(new_n984), .C2(new_n760), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n773), .A2(new_n235), .ZN(new_n986));
  INV_X1    g0786(.A(new_n251), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n780), .B1(new_n699), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n841), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n821), .A2(G283), .B1(G97), .B2(new_n784), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n845), .B2(new_n791), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT106), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n808), .A2(KEYINPUT46), .A3(G116), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(KEYINPUT46), .B1(new_n808), .B2(G116), .ZN(new_n995));
  XOR2_X1   g0795(.A(KEYINPUT107), .B(G317), .Z(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n802), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n268), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n801), .B2(new_n270), .C1(new_n855), .C2(new_n797), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n995), .B(new_n1000), .C1(G294), .C2(new_n852), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n994), .B(new_n1001), .C1(new_n992), .C2(new_n993), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n852), .A2(G159), .ZN(new_n1003));
  INV_X1    g0803(.A(G137), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n268), .B1(new_n802), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n801), .A2(new_n366), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(G143), .C2(new_n796), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n201), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n821), .A2(new_n1008), .B1(G58), .B2(new_n808), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n822), .A2(G150), .B1(G77), .B2(new_n784), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1003), .A2(new_n1007), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1002), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT47), .Z(new_n1013));
  OAI221_X1 g0813(.A(new_n989), .B1(new_n768), .B2(new_n956), .C1(new_n1013), .C2(new_n844), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n985), .A2(new_n1014), .ZN(G387));
  NAND3_X1  g0815(.A1(new_n976), .A2(new_n760), .A3(new_n977), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n770), .A2(new_n703), .B1(G107), .B2(new_n212), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n232), .A2(new_n287), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n703), .ZN(new_n1019));
  AOI211_X1 g0819(.A(G45), .B(new_n1019), .C1(G68), .C2(G77), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n247), .A2(G50), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT50), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n774), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1017), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n761), .B1(new_n1024), .B2(new_n780), .ZN(new_n1025));
  INV_X1    g0825(.A(G150), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n268), .B1(new_n802), .B2(new_n1026), .C1(new_n797), .C2(new_n373), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n987), .B2(new_n800), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n821), .A2(G68), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n795), .A2(new_n379), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n822), .B2(G50), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G77), .A2(new_n808), .B1(new_n784), .B2(G97), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n268), .B1(new_n998), .B2(G326), .ZN(new_n1034));
  INV_X1    g0834(.A(G283), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n807), .A2(new_n818), .B1(new_n801), .B2(new_n1035), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n821), .A2(G303), .B1(G322), .B2(new_n796), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n855), .B2(new_n851), .C1(new_n791), .C2(new_n996), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT48), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1036), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n1039), .B2(new_n1038), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT49), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1034), .B1(new_n524), .B2(new_n783), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1033), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1025), .B1(new_n1045), .B2(new_n778), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n683), .B2(new_n768), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n978), .A2(new_n701), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n756), .B1(new_n976), .B2(new_n977), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1016), .B(new_n1047), .C1(new_n1048), .C2(new_n1049), .ZN(G393));
  NAND2_X1  g0850(.A1(new_n983), .A2(new_n701), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n979), .B1(new_n973), .B2(new_n982), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n973), .A2(new_n760), .A3(new_n982), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n779), .B1(new_n518), .B2(new_n212), .C1(new_n774), .C2(new_n242), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n761), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n822), .A2(G311), .B1(G317), .B2(new_n796), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT52), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n852), .A2(G303), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n801), .A2(new_n524), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n268), .B(new_n1061), .C1(G322), .C2(new_n998), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n821), .A2(G294), .B1(G283), .B2(new_n808), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1060), .A2(new_n1062), .A3(new_n785), .A4(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n791), .A2(new_n373), .B1(new_n1026), .B2(new_n797), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT51), .Z(new_n1066));
  NAND2_X1  g0866(.A1(new_n852), .A2(new_n1008), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n801), .A2(new_n440), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n315), .B(new_n1068), .C1(G143), .C2(new_n998), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n821), .A2(new_n248), .B1(G68), .B2(new_n808), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1067), .A2(new_n1069), .A3(new_n854), .A4(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n1059), .A2(new_n1064), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1057), .B1(new_n1072), .B2(new_n778), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n945), .B2(new_n768), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1055), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1054), .A2(new_n1076), .ZN(G390));
  AOI21_X1  g0877(.A(new_n841), .B1(new_n379), .B2(new_n842), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n315), .B1(new_n998), .B2(G125), .ZN(new_n1079));
  INV_X1    g0879(.A(G128), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1079), .B1(new_n801), .B2(new_n373), .C1(new_n797), .C2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n808), .A2(G150), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT53), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1081), .B(new_n1083), .C1(G137), .C2(new_n852), .ZN(new_n1084));
  XOR2_X1   g0884(.A(KEYINPUT54), .B(G143), .Z(new_n1085));
  NAND2_X1  g0885(.A1(new_n821), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n866), .B2(new_n791), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n1008), .B2(new_n784), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n315), .B1(new_n801), .B2(new_n440), .C1(new_n797), .C2(new_n1035), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n809), .B1(new_n789), .B2(new_n518), .C1(new_n524), .C2(new_n791), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1089), .B(new_n1090), .C1(G107), .C2(new_n852), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n862), .B1(new_n818), .B2(new_n802), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT114), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1084), .A2(new_n1088), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1078), .B1(new_n1094), .B2(new_n844), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n917), .A2(new_n918), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1095), .B1(new_n1096), .B2(new_n765), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n836), .A2(new_n832), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n922), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n919), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1096), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n755), .A2(G330), .A3(new_n835), .A4(new_n922), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n832), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n715), .B2(new_n831), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n923), .A2(KEYINPUT108), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n922), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n919), .B1(new_n891), .B2(new_n909), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1103), .A2(new_n1104), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(KEYINPUT110), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n543), .B1(new_n511), .B2(new_n512), .ZN(new_n1117));
  AOI221_X4 g0917(.A(KEYINPUT85), .B1(new_n501), .B2(new_n507), .C1(new_n494), .C2(new_n498), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n1117), .A2(new_n894), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n752), .A2(new_n753), .ZN(new_n1120));
  OAI21_X1  g0920(.A(G330), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n922), .A2(new_n835), .ZN(new_n1122));
  OAI21_X1  g0922(.A(KEYINPUT109), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(G330), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n719), .B2(new_n893), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT109), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1125), .A2(new_n1126), .A3(new_n899), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n917), .A2(new_n918), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1128), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT110), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1103), .A2(new_n1132), .A3(new_n1104), .A4(new_n1114), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1116), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1098), .B1(new_n1134), .B2(new_n759), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(KEYINPUT115), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT115), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1137), .B(new_n1098), .C1(new_n1134), .C2(new_n759), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1125), .A2(new_n835), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1139), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1140), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n755), .A2(G330), .A3(new_n835), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n923), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(KEYINPUT111), .ZN(new_n1144));
  AND4_X1   g0944(.A1(new_n1126), .A2(new_n895), .A3(new_n899), .A4(G330), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1126), .B1(new_n1125), .B2(new_n899), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT111), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1142), .A2(new_n1148), .A3(new_n923), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1144), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1141), .B1(new_n1150), .B2(new_n1099), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n453), .A2(new_n1125), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n927), .A2(new_n647), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(KEYINPUT112), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT112), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1153), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1099), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1148), .B1(new_n1142), .B2(new_n923), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1128), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1157), .B1(new_n1159), .B2(new_n1149), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1155), .B(new_n1156), .C1(new_n1160), .C2(new_n1141), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1154), .A2(new_n1161), .A3(KEYINPUT113), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1096), .A2(new_n1102), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1132), .B1(new_n1164), .B2(new_n1104), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(KEYINPUT113), .B1(new_n1154), .B2(new_n1161), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n1162), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1154), .A2(new_n1161), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n701), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1136), .B(new_n1138), .C1(new_n1168), .C2(new_n1171), .ZN(G378));
  NAND2_X1  g0972(.A1(new_n1170), .A2(new_n1156), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT119), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n900), .B1(new_n890), .B2(new_n891), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n911), .B(G330), .C1(new_n1175), .C2(KEYINPUT40), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n342), .A2(new_n876), .ZN(new_n1177));
  XOR2_X1   g0977(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1178));
  XOR2_X1   g0978(.A(new_n1177), .B(new_n1178), .Z(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT117), .ZN(new_n1181));
  OR2_X1    g0981(.A1(new_n326), .A2(new_n344), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1181), .B1(new_n646), .B2(new_n1182), .ZN(new_n1183));
  AOI211_X1 g0983(.A(KEYINPUT117), .B(new_n634), .C1(new_n642), .C2(new_n645), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1180), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n643), .A2(new_n644), .A3(KEYINPUT91), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT91), .B1(new_n643), .B2(new_n644), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1182), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT117), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n646), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(new_n1190), .A3(new_n1179), .ZN(new_n1191));
  AND2_X1   g0991(.A1(new_n1185), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1176), .A2(new_n1192), .A3(KEYINPUT118), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1185), .A2(KEYINPUT118), .A3(new_n1191), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n904), .A2(new_n1194), .A3(G330), .A4(new_n911), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n926), .ZN(new_n1196));
  AND3_X1   g0996(.A1(new_n1193), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1196), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1174), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1200));
  OAI21_X1  g1000(.A(KEYINPUT119), .B1(new_n1200), .B2(new_n926), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1173), .A2(KEYINPUT57), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT57), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1153), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1203), .A2(new_n1207), .A3(new_n701), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n795), .A2(new_n866), .B1(new_n801), .B2(new_n1026), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n822), .A2(G128), .B1(new_n808), .B2(new_n1085), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n1004), .B2(new_n789), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1209), .B(new_n1211), .C1(G125), .C2(new_n796), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1213), .A2(KEYINPUT59), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1213), .A2(KEYINPUT59), .ZN(new_n1215));
  AOI211_X1 g1015(.A(G33), .B(G41), .C1(new_n998), .C2(G124), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n373), .B2(new_n783), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1217), .B(KEYINPUT116), .Z(new_n1218));
  NOR3_X1   g1018(.A1(new_n1214), .A2(new_n1215), .A3(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n783), .A2(new_n328), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G77), .B2(new_n808), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1221), .B1(new_n270), .B2(new_n791), .C1(new_n251), .C2(new_n789), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n315), .B(new_n286), .C1(new_n802), .C2(new_n1035), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n795), .A2(new_n518), .B1(new_n797), .B2(new_n524), .ZN(new_n1224));
  NOR4_X1   g1024(.A1(new_n1222), .A2(new_n1006), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1225), .A2(KEYINPUT58), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(KEYINPUT58), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n438), .B1(G33), .B2(G41), .C1(new_n700), .C2(new_n268), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n778), .B1(new_n1219), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n842), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1230), .B(new_n761), .C1(new_n1008), .C2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1192), .B2(new_n765), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1206), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1233), .B1(new_n1234), .B2(new_n760), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1208), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(G375));
  NAND2_X1  g1037(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NOR4_X1   g1039(.A1(new_n1162), .A2(new_n1167), .A3(new_n964), .A4(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n841), .B1(new_n366), .B2(new_n842), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n268), .B1(new_n998), .B2(G303), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1242), .B1(new_n801), .B2(new_n251), .C1(new_n797), .C2(new_n818), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n822), .A2(G283), .B1(G97), .B2(new_n808), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1244), .B1(new_n440), .B2(new_n783), .C1(new_n270), .C2(new_n789), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1243), .B(new_n1245), .C1(G116), .C2(new_n852), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1246), .A2(KEYINPUT120), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(KEYINPUT120), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n268), .B1(new_n802), .B2(new_n1080), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n1249), .B(new_n1220), .C1(G50), .C2(new_n800), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n797), .A2(new_n866), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1251), .A2(KEYINPUT121), .B1(new_n808), .B2(G159), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n852), .B2(new_n1085), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(G137), .A2(new_n822), .B1(new_n821), .B2(G150), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1254), .B(new_n1255), .C1(KEYINPUT121), .C2(new_n1251), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1247), .A2(new_n1248), .A3(new_n1256), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n1241), .B1(new_n844), .B2(new_n1257), .C1(new_n1111), .C2(new_n766), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n1151), .B2(new_n759), .ZN(new_n1259));
  OR2_X1    g1059(.A1(new_n1240), .A2(new_n1259), .ZN(G381));
  OR3_X1    g1060(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1261));
  NOR4_X1   g1061(.A1(G381), .A2(G387), .A3(G390), .A4(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1168), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1171), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1135), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1262), .A2(new_n1236), .A3(new_n1265), .ZN(G407));
  NAND4_X1  g1066(.A1(new_n1236), .A2(G213), .A3(new_n676), .A4(new_n1265), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(G407), .A2(G213), .A3(new_n1267), .ZN(G409));
  NAND2_X1  g1068(.A1(G387), .A2(KEYINPUT125), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT125), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n985), .A2(new_n1270), .A3(new_n1014), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(G393), .B(new_n828), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(G390), .A2(new_n1272), .ZN(new_n1273));
  OR3_X1    g1073(.A1(new_n1272), .A2(new_n1053), .A3(new_n1075), .ZN(new_n1274));
  AND4_X1   g1074(.A1(new_n1269), .A2(new_n1271), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1269), .A2(new_n1271), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1208), .A2(G378), .A3(new_n1235), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1233), .B1(new_n1202), .B2(new_n760), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1173), .A2(new_n1234), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1279), .B1(new_n1280), .B2(new_n964), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1265), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n1278), .A2(new_n1282), .B1(G213), .B2(new_n676), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT123), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT60), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n701), .B1(new_n1238), .B2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1154), .A2(new_n1161), .A3(KEYINPUT60), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1238), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT122), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1286), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1287), .A2(KEYINPUT122), .A3(new_n1238), .ZN(new_n1291));
  AOI211_X1 g1091(.A(new_n873), .B(new_n1259), .C1(new_n1290), .C2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1286), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(new_n1291), .A3(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1259), .ZN(new_n1296));
  AOI21_X1  g1096(.A(G384), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1284), .B1(new_n1292), .B2(new_n1297), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1287), .A2(KEYINPUT122), .A3(new_n1238), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT122), .B1(new_n1287), .B2(new_n1238), .ZN(new_n1300));
  NOR3_X1   g1100(.A1(new_n1299), .A2(new_n1300), .A3(new_n1286), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n873), .B1(new_n1301), .B2(new_n1259), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1295), .A2(G384), .A3(new_n1296), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1302), .A2(KEYINPUT123), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n676), .A2(G213), .ZN(new_n1305));
  INV_X1    g1105(.A(G2897), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1298), .A2(new_n1304), .A3(new_n1307), .ZN(new_n1308));
  OAI221_X1 g1108(.A(new_n1284), .B1(new_n1306), .B2(new_n1305), .C1(new_n1292), .C2(new_n1297), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT124), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1308), .A2(KEYINPUT124), .A3(new_n1309), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1283), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1292), .A2(new_n1297), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1315), .A2(new_n1305), .A3(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(KEYINPUT62), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT61), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT62), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1283), .A2(new_n1320), .A3(new_n1316), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1318), .A2(new_n1319), .A3(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1277), .B1(new_n1314), .B2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1283), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1313), .ZN(new_n1325));
  AOI21_X1  g1125(.A(KEYINPUT124), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1324), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1283), .A2(KEYINPUT63), .A3(new_n1316), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT63), .B1(new_n1283), .B2(new_n1316), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1319), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1327), .A2(new_n1328), .A3(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1323), .A2(new_n1332), .ZN(G405));
  INV_X1    g1133(.A(KEYINPUT127), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1277), .A2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT126), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1316), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1338));
  NOR3_X1   g1138(.A1(new_n1236), .A2(new_n1338), .A3(new_n1135), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1278), .ZN(new_n1340));
  OAI211_X1 g1140(.A(new_n1336), .B(new_n1337), .C1(new_n1339), .C2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(G375), .A2(new_n1265), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1337), .A2(new_n1336), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1316), .A2(KEYINPUT126), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1342), .A2(new_n1278), .A3(new_n1343), .A4(new_n1344), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1335), .A2(new_n1341), .A3(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(KEYINPUT127), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1346), .A2(new_n1348), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1335), .A2(new_n1341), .A3(new_n1345), .A4(new_n1347), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1349), .A2(new_n1350), .ZN(G402));
endmodule


