//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n631,
    new_n632, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n815, new_n816, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941;
  INV_X1    g000(.A(KEYINPUT40), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT4), .ZN(new_n203));
  INV_X1    g002(.A(G148gat), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT72), .B1(new_n204), .B2(G141gat), .ZN(new_n205));
  OR3_X1    g004(.A1(new_n204), .A2(KEYINPUT72), .A3(G141gat), .ZN(new_n206));
  XOR2_X1   g005(.A(KEYINPUT73), .B(G148gat), .Z(new_n207));
  INV_X1    g006(.A(G141gat), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n205), .B(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(G155gat), .B(G162gat), .Z(new_n210));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n211), .B1(KEYINPUT74), .B2(G155gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT75), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n209), .A2(KEYINPUT75), .A3(new_n213), .ZN(new_n217));
  XOR2_X1   g016(.A(G141gat), .B(G148gat), .Z(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(new_n211), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n216), .A2(new_n217), .B1(new_n210), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G113gat), .B(G120gat), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT1), .B1(new_n221), .B2(KEYINPUT67), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(KEYINPUT67), .B2(new_n221), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224));
  INV_X1    g023(.A(G134gat), .ZN(new_n225));
  NOR3_X1   g024(.A1(new_n224), .A2(new_n225), .A3(G127gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(G127gat), .B(G134gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n226), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G113gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G120gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT68), .B(G120gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n230), .B1(new_n231), .B2(new_n229), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT1), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n227), .A2(new_n233), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n223), .A2(new_n228), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n203), .B1(new_n220), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n203), .A3(new_n235), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT79), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT80), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n240), .B1(new_n238), .B2(new_n239), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n237), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n243), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n245), .A2(new_n236), .A3(new_n241), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n220), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n248), .A2(new_n235), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n220), .A2(new_n247), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n244), .A2(new_n246), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT39), .ZN(new_n253));
  NAND2_X1  g052(.A1(G225gat), .A2(G233gat), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n252), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(G57gat), .B(G85gat), .Z(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT78), .ZN(new_n258));
  XOR2_X1   g057(.A(G1gat), .B(G29gat), .Z(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n260), .B(new_n261), .Z(new_n262));
  NAND2_X1  g061(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n220), .B(new_n235), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n264), .A2(new_n255), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT39), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n266), .B1(new_n252), .B2(new_n255), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n202), .B1(new_n263), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n267), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n269), .A2(KEYINPUT40), .A3(new_n262), .A4(new_n256), .ZN(new_n270));
  AOI211_X1 g069(.A(KEYINPUT5), .B(new_n255), .C1(new_n249), .C2(new_n250), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n244), .A2(new_n271), .A3(new_n246), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n273), .B1(new_n264), .B2(new_n255), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n236), .A2(KEYINPUT76), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n251), .A2(new_n254), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT76), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n237), .A2(new_n277), .A3(new_n238), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n274), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n272), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n262), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n283));
  INV_X1    g082(.A(G169gat), .ZN(new_n284));
  INV_X1    g083(.A(G176gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287));
  OR3_X1    g086(.A1(new_n286), .A2(KEYINPUT26), .A3(new_n287), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n287), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n289));
  XOR2_X1   g088(.A(KEYINPUT27), .B(G183gat), .Z(new_n290));
  INV_X1    g089(.A(KEYINPUT28), .ZN(new_n291));
  NOR3_X1   g090(.A1(new_n290), .A2(new_n291), .A3(G190gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n293));
  AOI21_X1  g092(.A(G190gat), .B1(new_n293), .B2(KEYINPUT27), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT27), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n295), .A2(KEYINPUT65), .A3(G183gat), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT28), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n288), .B(new_n289), .C1(new_n292), .C2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n287), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT23), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n299), .B1(new_n286), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n301), .B1(new_n300), .B2(new_n299), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT24), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n303), .A2(G183gat), .A3(G190gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(G183gat), .B(G190gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n304), .B1(new_n305), .B2(new_n303), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT25), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT64), .B(G176gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(KEYINPUT23), .A3(new_n284), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT25), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(new_n310), .A3(new_n301), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n298), .B(new_n307), .C1(new_n306), .C2(new_n311), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n312), .A2(G226gat), .A3(G233gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT29), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n312), .A2(new_n314), .B1(G226gat), .B2(G233gat), .ZN(new_n315));
  XOR2_X1   g114(.A(G197gat), .B(G204gat), .Z(new_n316));
  AOI21_X1  g115(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G211gat), .B(G218gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  OR3_X1    g120(.A1(new_n313), .A2(new_n315), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n321), .B1(new_n313), .B2(new_n315), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XOR2_X1   g123(.A(G8gat), .B(G36gat), .Z(new_n325));
  XNOR2_X1  g124(.A(new_n325), .B(KEYINPUT71), .ZN(new_n326));
  XNOR2_X1  g125(.A(G64gat), .B(G92gat), .ZN(new_n327));
  XOR2_X1   g126(.A(new_n326), .B(new_n327), .Z(new_n328));
  OAI21_X1  g127(.A(new_n283), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n328), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n322), .A2(KEYINPUT30), .A3(new_n323), .A4(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n324), .A2(new_n328), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n329), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n268), .A2(new_n270), .A3(new_n282), .A4(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G228gat), .ZN(new_n335));
  INV_X1    g134(.A(G233gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT3), .B1(new_n320), .B2(new_n314), .ZN(new_n338));
  OR2_X1    g137(.A1(new_n220), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT82), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n337), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n220), .A2(new_n338), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n320), .B1(new_n250), .B2(new_n314), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT29), .B1(new_n220), .B2(new_n247), .ZN(new_n345));
  OAI221_X1 g144(.A(new_n339), .B1(new_n340), .B2(new_n337), .C1(new_n345), .C2(new_n320), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G22gat), .ZN(new_n348));
  INV_X1    g147(.A(G22gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n344), .A2(new_n349), .A3(new_n346), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT31), .B(G50gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT81), .ZN(new_n353));
  XOR2_X1   g152(.A(G78gat), .B(G106gat), .Z(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n349), .B1(new_n344), .B2(new_n346), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n355), .B1(new_n356), .B2(KEYINPUT83), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n351), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n348), .A2(KEYINPUT83), .A3(new_n350), .A4(new_n355), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n334), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n262), .B1(new_n272), .B2(new_n279), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT84), .B1(new_n363), .B2(KEYINPUT6), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n324), .A2(new_n328), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(KEYINPUT38), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n330), .B1(new_n324), .B2(KEYINPUT37), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n368), .B1(KEYINPUT37), .B2(new_n324), .ZN(new_n369));
  MUX2_X1   g168(.A(KEYINPUT38), .B(new_n367), .S(new_n369), .Z(new_n370));
  INV_X1    g169(.A(KEYINPUT6), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n272), .A2(new_n279), .A3(new_n262), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n282), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n363), .A2(KEYINPUT6), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT84), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n365), .B(new_n370), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n377), .ZN(new_n378));
  XOR2_X1   g177(.A(KEYINPUT69), .B(KEYINPUT34), .Z(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  OR2_X1    g179(.A1(new_n312), .A2(new_n235), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n312), .A2(new_n235), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n381), .A2(G227gat), .A3(G233gat), .A4(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT33), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  XOR2_X1   g184(.A(G15gat), .B(G43gat), .Z(new_n386));
  XNOR2_X1  g185(.A(G71gat), .B(G99gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n386), .B(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n380), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n381), .A2(new_n382), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT32), .ZN(new_n392));
  INV_X1    g191(.A(G227gat), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n391), .B(new_n392), .C1(new_n393), .C2(new_n336), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n391), .B1(new_n393), .B2(new_n336), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(KEYINPUT32), .A3(new_n383), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n385), .A2(new_n380), .A3(new_n388), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n390), .A2(new_n394), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n394), .ZN(new_n399));
  INV_X1    g198(.A(new_n397), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n399), .B1(new_n400), .B2(new_n389), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT70), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT36), .ZN(new_n404));
  OR2_X1    g203(.A1(new_n403), .A2(KEYINPUT36), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n398), .A2(new_n401), .A3(new_n403), .A4(KEYINPUT36), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n333), .B1(new_n373), .B2(new_n374), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n408), .B1(new_n409), .B2(new_n361), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n378), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n402), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n360), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT35), .ZN(new_n416));
  INV_X1    g215(.A(new_n333), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n358), .A2(new_n402), .A3(new_n417), .A4(new_n359), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT85), .B(KEYINPUT35), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n376), .B1(new_n373), .B2(new_n374), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n419), .B(new_n421), .C1(new_n422), .C2(new_n364), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n416), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n412), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G15gat), .B(G22gat), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT16), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n426), .B1(new_n427), .B2(G1gat), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n428), .B1(G1gat), .B2(new_n426), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(G8gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(G71gat), .ZN(new_n432));
  INV_X1    g231(.A(G78gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(G71gat), .A2(G78gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g235(.A1(G57gat), .A2(G64gat), .ZN(new_n437));
  NOR2_X1   g236(.A1(G57gat), .A2(G64gat), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n436), .B1(new_n439), .B2(KEYINPUT9), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n432), .A2(new_n433), .A3(KEYINPUT9), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT90), .B1(new_n437), .B2(new_n438), .ZN(new_n443));
  INV_X1    g242(.A(G57gat), .ZN(new_n444));
  INV_X1    g243(.A(G64gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT90), .ZN(new_n447));
  NAND2_X1  g246(.A1(G57gat), .A2(G64gat), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI221_X4 g248(.A(KEYINPUT91), .B1(new_n435), .B2(new_n442), .C1(new_n443), .C2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT91), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n443), .A2(new_n449), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n442), .A2(new_n435), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n441), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT92), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(KEYINPUT92), .B(new_n441), .C1(new_n450), .C2(new_n454), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT21), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n459), .A2(KEYINPUT21), .ZN(new_n461));
  NAND2_X1  g260(.A1(G231gat), .A2(G233gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(G127gat), .ZN(new_n464));
  OAI211_X1 g263(.A(G231gat), .B(G233gat), .C1(new_n459), .C2(KEYINPUT21), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n464), .B1(new_n463), .B2(new_n465), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n431), .B(new_n460), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n468), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n460), .A2(new_n431), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n471), .A3(new_n466), .ZN(new_n472));
  XOR2_X1   g271(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(G155gat), .ZN(new_n474));
  XOR2_X1   g273(.A(G183gat), .B(G211gat), .Z(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n469), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n476), .B1(new_n469), .B2(new_n472), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(G190gat), .B(G218gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(G99gat), .A2(G106gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT8), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT95), .ZN(new_n483));
  OR2_X1    g282(.A1(G85gat), .A2(G92gat), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n483), .B1(new_n482), .B2(new_n484), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G85gat), .A2(G92gat), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n488), .A2(KEYINPUT94), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT93), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT7), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT7), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n492), .B1(new_n488), .B2(KEYINPUT93), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n491), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  XOR2_X1   g293(.A(G99gat), .B(G106gat), .Z(new_n495));
  NOR3_X1   g294(.A1(new_n487), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n495), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n484), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT95), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n484), .A3(new_n483), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n493), .A2(new_n489), .ZN(new_n502));
  NOR4_X1   g301(.A1(new_n488), .A2(new_n492), .A3(KEYINPUT93), .A4(KEYINPUT94), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n497), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n496), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT14), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n507), .B1(G29gat), .B2(G36gat), .ZN(new_n508));
  OR3_X1    g307(.A1(new_n507), .A2(G29gat), .A3(G36gat), .ZN(new_n509));
  XOR2_X1   g308(.A(KEYINPUT87), .B(G36gat), .Z(new_n510));
  INV_X1    g309(.A(G29gat), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n508), .B(new_n509), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G43gat), .ZN(new_n513));
  INV_X1    g312(.A(G50gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(G43gat), .A2(G50gat), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT15), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT88), .B(G43gat), .ZN(new_n519));
  AOI211_X1 g318(.A(KEYINPUT15), .B(new_n515), .C1(new_n519), .C2(new_n514), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n517), .B1(new_n520), .B2(new_n512), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT17), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n518), .A2(new_n521), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n506), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n495), .B1(new_n487), .B2(new_n494), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n501), .A2(new_n504), .A3(new_n497), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n528), .B1(new_n524), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT96), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n527), .A2(new_n532), .A3(KEYINPUT96), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n480), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n535), .ZN(new_n537));
  INV_X1    g336(.A(new_n480), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n537), .A2(new_n538), .A3(new_n533), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G134gat), .B(G162gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT41), .ZN(new_n542));
  INV_X1    g341(.A(G232gat), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n542), .B1(new_n543), .B2(new_n336), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n541), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT97), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n545), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n536), .A2(KEYINPUT97), .A3(new_n548), .A4(new_n539), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT98), .B1(new_n479), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT98), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n550), .B(new_n553), .C1(new_n477), .C2(new_n478), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n523), .A2(new_n526), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(new_n431), .ZN(new_n557));
  NAND2_X1  g356(.A1(G229gat), .A2(G233gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT89), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n522), .A2(new_n430), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT18), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n557), .A2(KEYINPUT18), .A3(new_n559), .A4(new_n560), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n431), .A2(new_n524), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n560), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n559), .B(KEYINPUT13), .Z(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n563), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G113gat), .B(G141gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT86), .B(G197gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(KEYINPUT11), .B(G169gat), .Z(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT12), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n563), .A2(new_n564), .A3(new_n568), .A4(new_n575), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NOR3_X1   g378(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT90), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n447), .B1(new_n446), .B2(new_n448), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n453), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT91), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n452), .A2(new_n451), .A3(new_n453), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT92), .B1(new_n585), .B2(new_n441), .ZN(new_n586));
  INV_X1    g385(.A(new_n458), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n531), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT100), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n440), .B1(new_n583), .B2(new_n584), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n531), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n588), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT101), .ZN(new_n595));
  INV_X1    g394(.A(new_n590), .ZN(new_n596));
  XOR2_X1   g395(.A(KEYINPUT99), .B(KEYINPUT10), .Z(new_n597));
  AOI21_X1  g396(.A(new_n597), .B1(new_n588), .B2(new_n593), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n459), .A2(KEYINPUT10), .A3(new_n506), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n596), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G120gat), .B(G148gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(G176gat), .B(G204gat), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n603), .B(new_n604), .Z(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  OR3_X1    g405(.A1(new_n595), .A2(new_n602), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n606), .B1(new_n595), .B2(new_n602), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n555), .A2(new_n579), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n425), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n375), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(G1gat), .ZN(G1324gat));
  INV_X1    g414(.A(G8gat), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n616), .B1(new_n613), .B2(new_n333), .ZN(new_n617));
  XNOR2_X1  g416(.A(KEYINPUT102), .B(KEYINPUT16), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(new_n616), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n612), .A2(new_n417), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(KEYINPUT42), .B1(new_n617), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n621), .B1(KEYINPUT42), .B2(new_n620), .ZN(G1325gat));
  NAND2_X1  g421(.A1(new_n406), .A2(new_n407), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT104), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n613), .A2(G15gat), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(G15gat), .B1(new_n613), .B2(new_n402), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n627), .A2(KEYINPUT103), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(KEYINPUT103), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(G1326gat));
  NOR2_X1   g429(.A1(new_n612), .A2(new_n361), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT43), .B(G22gat), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(G1327gat));
  AOI21_X1  g432(.A(new_n550), .B1(new_n412), .B2(new_n424), .ZN(new_n634));
  INV_X1    g433(.A(new_n479), .ZN(new_n635));
  INV_X1    g434(.A(new_n579), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n635), .A2(new_n636), .A3(new_n609), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n373), .A2(new_n374), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n638), .A2(G29gat), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n640), .B(KEYINPUT45), .Z(new_n641));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n410), .B1(new_n362), .B2(new_n377), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT106), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n364), .B1(new_n639), .B2(KEYINPUT84), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n361), .A2(new_n417), .A3(new_n402), .A4(new_n421), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT35), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n648), .B1(new_n409), .B2(new_n414), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n644), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n416), .A2(new_n423), .A3(KEYINPUT106), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n643), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n642), .B1(new_n652), .B2(new_n550), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n634), .A2(KEYINPUT44), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n637), .B(KEYINPUT105), .Z(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(G29gat), .B1(new_n657), .B2(new_n639), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n641), .A2(new_n658), .ZN(G1328gat));
  INV_X1    g458(.A(KEYINPUT46), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n333), .B(new_n510), .C1(KEYINPUT107), .C2(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n638), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(KEYINPUT107), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n653), .A2(new_n333), .A3(new_n654), .A4(new_n656), .ZN(new_n665));
  INV_X1    g464(.A(new_n510), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT108), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT108), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n664), .A2(new_n670), .A3(new_n667), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(G1329gat));
  INV_X1    g471(.A(new_n519), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n673), .B1(new_n657), .B2(new_n408), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n638), .A2(new_n413), .A3(new_n673), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT47), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n655), .A2(new_n625), .A3(new_n656), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n675), .B1(new_n679), .B2(new_n673), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n678), .B1(new_n680), .B2(KEYINPUT47), .ZN(G1330gat));
  AOI211_X1 g480(.A(G50gat), .B(new_n361), .C1(new_n638), .C2(KEYINPUT109), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(KEYINPUT109), .B2(new_n638), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n653), .A2(new_n360), .A3(new_n654), .A4(new_n656), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(G50gat), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT48), .B1(new_n685), .B2(KEYINPUT110), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n683), .B(new_n685), .C1(KEYINPUT110), .C2(KEYINPUT48), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(G1331gat));
  NOR3_X1   g489(.A1(new_n647), .A2(new_n644), .A3(new_n649), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT106), .B1(new_n416), .B2(new_n423), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n412), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n555), .A2(new_n636), .A3(new_n609), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n639), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(new_n444), .ZN(G1332gat));
  NAND2_X1  g496(.A1(new_n695), .A2(KEYINPUT111), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT111), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n693), .A2(new_n699), .A3(new_n694), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n417), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n698), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(KEYINPUT112), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT112), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n698), .A2(new_n704), .A3(new_n700), .A4(new_n701), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1333gat));
  AND2_X1   g507(.A1(new_n698), .A2(new_n700), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n709), .A2(G71gat), .A3(new_n625), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n432), .B1(new_n695), .B2(new_n413), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n710), .A2(KEYINPUT50), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT50), .B1(new_n710), .B2(new_n711), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(G1334gat));
  NAND2_X1  g513(.A1(new_n709), .A2(new_n360), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g515(.A1(new_n635), .A2(new_n579), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(new_n610), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n653), .A2(new_n654), .A3(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(G85gat), .B1(new_n721), .B2(new_n639), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n693), .A2(new_n551), .A3(new_n717), .ZN(new_n723));
  NAND2_X1  g522(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n650), .A2(new_n651), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n550), .B1(new_n726), .B2(new_n412), .ZN(new_n727));
  INV_X1    g526(.A(new_n724), .ZN(new_n728));
  NOR2_X1   g527(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n727), .A2(new_n717), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n725), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n639), .A2(G85gat), .A3(new_n610), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT114), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n722), .B1(new_n734), .B2(new_n736), .ZN(G1336gat));
  INV_X1    g536(.A(G92gat), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n738), .B1(new_n720), .B2(new_n333), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n609), .A2(new_n738), .A3(new_n333), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT115), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n733), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n740), .A2(new_n741), .A3(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n744), .ZN(new_n746));
  OAI21_X1  g545(.A(KEYINPUT52), .B1(new_n746), .B2(new_n739), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1337gat));
  OAI21_X1  g547(.A(G99gat), .B1(new_n721), .B2(new_n624), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n610), .A2(new_n413), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  OR2_X1    g550(.A1(new_n751), .A2(G99gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n749), .B1(new_n734), .B2(new_n752), .ZN(G1338gat));
  INV_X1    g552(.A(KEYINPUT117), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n361), .A2(new_n610), .A3(G106gat), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n728), .B1(new_n727), .B2(new_n717), .ZN(new_n756));
  NOR4_X1   g555(.A1(new_n652), .A2(new_n550), .A3(new_n718), .A4(new_n730), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n653), .A2(new_n360), .A3(new_n654), .A4(new_n719), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G106gat), .ZN(new_n760));
  XOR2_X1   g559(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n761));
  AND4_X1   g560(.A1(new_n754), .A2(new_n758), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  AOI22_X1  g561(.A1(new_n733), .A2(new_n755), .B1(new_n759), .B2(G106gat), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n754), .B1(new_n763), .B2(new_n761), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n758), .A2(new_n760), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT53), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n762), .B1(new_n764), .B2(new_n766), .ZN(G1339gat));
  NAND4_X1  g566(.A1(new_n552), .A2(new_n636), .A3(new_n554), .A4(new_n610), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT54), .ZN(new_n770));
  INV_X1    g569(.A(new_n597), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n506), .B1(new_n457), .B2(new_n458), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n772), .B2(new_n592), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n599), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n770), .B1(new_n774), .B2(new_n596), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n773), .A2(new_n590), .A3(new_n599), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n769), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n770), .B(new_n596), .C1(new_n598), .C2(new_n600), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n778), .A2(new_n779), .A3(new_n606), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n779), .B1(new_n778), .B2(new_n606), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n777), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n601), .A2(KEYINPUT54), .A3(new_n776), .ZN(new_n783));
  AOI211_X1 g582(.A(KEYINPUT54), .B(new_n590), .C1(new_n773), .C2(new_n599), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT118), .B1(new_n784), .B2(new_n605), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n778), .A2(new_n779), .A3(new_n606), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n783), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n607), .B(new_n782), .C1(new_n787), .C2(KEYINPUT55), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n559), .B1(new_n557), .B2(new_n560), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n566), .A2(new_n567), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n574), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n791), .A2(KEYINPUT119), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(KEYINPUT119), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(new_n578), .A3(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n788), .A2(new_n550), .A3(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n609), .A2(new_n578), .A3(new_n792), .A4(new_n793), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(new_n636), .B2(new_n788), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n795), .B1(new_n797), .B2(new_n550), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n768), .B1(new_n798), .B2(new_n635), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n361), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT120), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n800), .B(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n802), .A2(new_n402), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n639), .A2(new_n333), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n805), .A2(new_n229), .A3(new_n636), .ZN(new_n806));
  INV_X1    g605(.A(new_n799), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n807), .A2(new_n639), .A3(new_n418), .ZN(new_n808));
  AOI21_X1  g607(.A(G113gat), .B1(new_n808), .B2(new_n579), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n806), .A2(new_n809), .ZN(G1340gat));
  OAI21_X1  g609(.A(G120gat), .B1(new_n805), .B2(new_n610), .ZN(new_n811));
  INV_X1    g610(.A(new_n231), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n808), .A2(new_n812), .A3(new_n609), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(G1341gat));
  OAI21_X1  g613(.A(G127gat), .B1(new_n805), .B2(new_n479), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n808), .A2(new_n464), .A3(new_n635), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(G1342gat));
  OAI21_X1  g616(.A(G134gat), .B1(new_n805), .B2(new_n550), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n808), .A2(new_n225), .A3(new_n551), .ZN(new_n819));
  XOR2_X1   g618(.A(new_n819), .B(KEYINPUT56), .Z(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(G1343gat));
  NAND2_X1  g620(.A1(new_n799), .A2(new_n360), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(KEYINPUT57), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n804), .A2(new_n408), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n795), .ZN(new_n826));
  INV_X1    g625(.A(new_n796), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT121), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n636), .B1(new_n788), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n780), .A2(new_n781), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n769), .B1(new_n830), .B2(new_n783), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n831), .A2(KEYINPUT121), .A3(new_n607), .A4(new_n782), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n827), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n550), .B1(new_n833), .B2(KEYINPUT122), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT122), .ZN(new_n835));
  AOI211_X1 g634(.A(new_n835), .B(new_n827), .C1(new_n829), .C2(new_n832), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n826), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n479), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n361), .B1(new_n838), .B2(new_n768), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n579), .B(new_n825), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(G141gat), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT123), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n624), .A2(new_n360), .ZN(new_n844));
  NOR4_X1   g643(.A1(new_n807), .A2(new_n639), .A3(new_n333), .A4(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n845), .A2(new_n208), .A3(new_n579), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n843), .A2(new_n847), .A3(KEYINPUT58), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n842), .B(new_n846), .C1(KEYINPUT123), .C2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(G1344gat));
  INV_X1    g650(.A(new_n207), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n845), .A2(new_n852), .A3(new_n609), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n823), .A2(new_n824), .ZN(new_n854));
  INV_X1    g653(.A(new_n839), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n854), .B1(new_n855), .B2(KEYINPUT57), .ZN(new_n856));
  AOI211_X1 g655(.A(KEYINPUT59), .B(new_n852), .C1(new_n856), .C2(new_n609), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n361), .A2(KEYINPUT57), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n829), .A2(new_n832), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n835), .B1(new_n860), .B2(new_n827), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n833), .A2(KEYINPUT122), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n550), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n635), .B1(new_n863), .B2(new_n826), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT124), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n768), .B(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n859), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n822), .A2(KEYINPUT57), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n824), .A2(new_n610), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n858), .B1(new_n870), .B2(G148gat), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n853), .B1(new_n857), .B2(new_n871), .ZN(G1345gat));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n635), .ZN(new_n873));
  XNOR2_X1  g672(.A(KEYINPUT74), .B(G155gat), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n479), .A2(new_n874), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n845), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(G1346gat));
  AOI21_X1  g677(.A(G162gat), .B1(new_n845), .B2(new_n551), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n551), .A2(G162gat), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n856), .B2(new_n880), .ZN(G1347gat));
  NOR2_X1   g680(.A1(new_n375), .A2(new_n417), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n882), .B(KEYINPUT125), .Z(new_n883));
  NAND3_X1  g682(.A1(new_n802), .A2(new_n402), .A3(new_n883), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n884), .A2(new_n284), .A3(new_n636), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n807), .A2(new_n375), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n886), .A2(new_n333), .A3(new_n414), .ZN(new_n887));
  AOI21_X1  g686(.A(G169gat), .B1(new_n887), .B2(new_n579), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n885), .A2(new_n888), .ZN(G1348gat));
  AOI21_X1  g688(.A(G176gat), .B1(new_n887), .B2(new_n609), .ZN(new_n890));
  INV_X1    g689(.A(new_n883), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n891), .A2(new_n308), .A3(new_n751), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n890), .B1(new_n802), .B2(new_n892), .ZN(G1349gat));
  OAI21_X1  g692(.A(G183gat), .B1(new_n884), .B2(new_n479), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n479), .A2(new_n290), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n887), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT60), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT60), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n894), .A2(new_n899), .A3(new_n896), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(G1350gat));
  INV_X1    g700(.A(G190gat), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n887), .A2(new_n902), .A3(new_n551), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n803), .A2(new_n551), .A3(new_n883), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(G190gat), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n904), .B(G190gat), .C1(new_n884), .C2(new_n550), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n903), .B1(new_n906), .B2(new_n908), .ZN(G1351gat));
  NOR2_X1   g708(.A1(new_n844), .A2(new_n417), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n886), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(G197gat), .B1(new_n911), .B2(new_n579), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n891), .A2(new_n625), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n866), .B1(new_n837), .B2(new_n479), .ZN(new_n914));
  INV_X1    g713(.A(new_n859), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n913), .B(new_n868), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n579), .A2(G197gat), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n912), .B1(new_n917), .B2(new_n918), .ZN(G1352gat));
  INV_X1    g718(.A(G204gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n911), .A2(new_n920), .A3(new_n609), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n921), .B(KEYINPUT62), .Z(new_n922));
  OAI21_X1  g721(.A(G204gat), .B1(new_n916), .B2(new_n610), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1353gat));
  INV_X1    g723(.A(KEYINPUT63), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n925), .B(G211gat), .C1(new_n916), .C2(new_n479), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n479), .A2(G211gat), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n886), .A2(new_n910), .A3(new_n927), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT126), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n867), .A2(new_n635), .A3(new_n868), .A4(new_n913), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n925), .B1(new_n931), .B2(G211gat), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT127), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(G211gat), .B1(new_n916), .B2(new_n479), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(KEYINPUT63), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT127), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n935), .A2(new_n936), .A3(new_n926), .A4(new_n929), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n933), .A2(new_n937), .ZN(G1354gat));
  OAI21_X1  g737(.A(G218gat), .B1(new_n916), .B2(new_n550), .ZN(new_n939));
  INV_X1    g738(.A(G218gat), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n911), .A2(new_n940), .A3(new_n551), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1355gat));
endmodule


