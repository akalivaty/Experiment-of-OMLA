//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 1 1 1 1 0 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1232, new_n1233, new_n1234, new_n1235, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  AOI22_X1  g0008(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n211), .B1(KEYINPUT64), .B2(new_n214), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n214), .A2(KEYINPUT64), .ZN(new_n216));
  AOI22_X1  g0016(.A1(new_n215), .A2(new_n216), .B1(G1), .B2(G20), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT65), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT0), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(new_n201), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n224), .B1(new_n228), .B2(new_n230), .C1(new_n217), .C2(new_n218), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n220), .A2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT66), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n236), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n226), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G150), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n226), .A2(new_n253), .ZN(new_n254));
  OAI22_X1  g0054(.A1(new_n250), .A2(new_n251), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n255), .B1(G20), .B2(new_n203), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n225), .B1(new_n221), .B2(new_n253), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n261), .B(new_n225), .C1(new_n253), .C2(new_n221), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n260), .A2(G20), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G50), .A3(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(G50), .B2(new_n261), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT9), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n267), .B(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G41), .A2(G45), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(G1), .ZN(new_n271));
  AND2_X1   g0071(.A1(G1), .A2(G13), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n271), .A2(new_n274), .A3(G274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(KEYINPUT67), .B1(new_n270), .B2(G1), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT67), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n278), .B(new_n260), .C1(G41), .C2(G45), .ZN(new_n279));
  AND3_X1   g0079(.A1(new_n277), .A2(new_n274), .A3(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n280), .A2(G226), .ZN(new_n281));
  AND2_X1   g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(new_n225), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT3), .B(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(G222), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G77), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(G1698), .ZN(new_n288));
  INV_X1    g0088(.A(G223), .ZN(new_n289));
  OAI221_X1 g0089(.A(new_n286), .B1(new_n287), .B2(new_n284), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  AOI211_X1 g0090(.A(new_n276), .B(new_n281), .C1(new_n283), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G190), .ZN(new_n292));
  INV_X1    g0092(.A(G200), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n269), .B(new_n292), .C1(new_n293), .C2(new_n291), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT10), .ZN(new_n295));
  INV_X1    g0095(.A(G179), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  OAI221_X1 g0097(.A(new_n297), .B1(G169), .B2(new_n291), .C1(new_n259), .C2(new_n266), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(KEYINPUT73), .B(KEYINPUT14), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT3), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G33), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n301), .A2(new_n303), .A3(G232), .A4(G1698), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n301), .A2(new_n303), .A3(G226), .A4(new_n285), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n304), .B(new_n305), .C1(new_n253), .C2(new_n205), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n283), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n277), .A2(G238), .A3(new_n274), .A4(new_n279), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n308), .A2(new_n275), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT13), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n307), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n310), .B1(new_n307), .B2(new_n309), .ZN(new_n312));
  OAI211_X1 g0112(.A(G169), .B(new_n300), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n307), .A2(new_n309), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT13), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n307), .A2(new_n309), .A3(new_n310), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(G179), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT14), .ZN(new_n319));
  OAI21_X1  g0119(.A(G169), .B1(new_n311), .B2(new_n312), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT72), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G169), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(new_n315), .B2(new_n316), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT72), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n318), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n226), .A2(G33), .A3(G77), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n327), .B1(new_n226), .B2(G68), .C1(new_n254), .C2(new_n202), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT70), .ZN(new_n329));
  AND3_X1   g0129(.A1(new_n328), .A2(new_n329), .A3(new_n257), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n329), .B1(new_n328), .B2(new_n257), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT11), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n328), .A2(new_n257), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT70), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT11), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n328), .A2(new_n329), .A3(new_n257), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G13), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n338), .A2(G1), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n226), .A2(G68), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT12), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n339), .B(new_n340), .C1(KEYINPUT71), .C2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT71), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n342), .B1(new_n343), .B2(KEYINPUT12), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n339), .A2(new_n340), .A3(KEYINPUT71), .A4(new_n341), .ZN(new_n345));
  INV_X1    g0145(.A(G68), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(new_n260), .B2(G20), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n344), .A2(new_n345), .B1(new_n263), .B2(new_n347), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n332), .A2(new_n337), .A3(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n326), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT69), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n315), .A2(new_n316), .ZN(new_n353));
  INV_X1    g0153(.A(G190), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n311), .A2(new_n312), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n356), .A2(KEYINPUT69), .A3(G190), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n349), .B1(new_n356), .B2(new_n293), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n351), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G238), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n288), .A2(new_n363), .B1(new_n206), .B2(new_n284), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n301), .A2(new_n303), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n365), .A2(new_n238), .A3(G1698), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n283), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n276), .B1(new_n280), .B2(G244), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n323), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n264), .A2(G77), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n262), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n261), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n372), .B1(new_n287), .B2(new_n373), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n250), .A2(new_n254), .B1(new_n226), .B2(new_n287), .ZN(new_n375));
  XNOR2_X1  g0175(.A(KEYINPUT15), .B(G87), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n376), .A2(new_n251), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n257), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n370), .A2(new_n379), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n367), .A2(new_n368), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n380), .B1(new_n296), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT68), .B1(new_n381), .B2(new_n293), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n369), .A2(new_n354), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n379), .B1(new_n384), .B2(KEYINPUT68), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR4_X1   g0188(.A1(new_n299), .A2(new_n362), .A3(new_n382), .A4(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n238), .B1(new_n272), .B2(new_n273), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n390), .A2(new_n277), .A3(new_n279), .ZN(new_n391));
  AND3_X1   g0191(.A1(new_n391), .A2(KEYINPUT74), .A3(new_n275), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT74), .B1(new_n391), .B2(new_n275), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT75), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n391), .A2(new_n275), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT74), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT75), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n391), .A2(KEYINPUT74), .A3(new_n275), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AND2_X1   g0200(.A1(KEYINPUT76), .A2(G190), .ZN(new_n401));
  NOR2_X1   g0201(.A1(KEYINPUT76), .A2(G190), .ZN(new_n402));
  OR2_X1    g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n284), .A2(G223), .A3(new_n285), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G87), .ZN(new_n405));
  INV_X1    g0205(.A(G226), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n404), .B(new_n405), .C1(new_n288), .C2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n403), .B1(new_n407), .B2(new_n283), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n394), .A2(new_n400), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n283), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n410), .A2(new_n397), .A3(new_n399), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n293), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n250), .B1(new_n260), .B2(G20), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(new_n263), .B1(new_n373), .B2(new_n250), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT7), .B1(new_n365), .B2(new_n226), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT7), .ZN(new_n418));
  AOI211_X1 g0218(.A(new_n418), .B(G20), .C1(new_n301), .C2(new_n303), .ZN(new_n419));
  OAI21_X1  g0219(.A(G68), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(G58), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n421), .A2(new_n346), .ZN(new_n422));
  OAI21_X1  g0222(.A(G20), .B1(new_n422), .B2(new_n201), .ZN(new_n423));
  INV_X1    g0223(.A(new_n254), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G159), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n420), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT16), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n258), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n420), .A2(KEYINPUT16), .A3(new_n427), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n416), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT77), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n413), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n433), .B1(new_n413), .B2(new_n432), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT17), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT17), .B1(new_n413), .B2(new_n432), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n418), .B1(new_n284), .B2(G20), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n365), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n346), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n429), .B1(new_n442), .B2(new_n426), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n431), .A2(new_n443), .A3(new_n257), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n415), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n394), .A2(new_n400), .A3(new_n296), .A4(new_n410), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n411), .A2(new_n323), .ZN(new_n447));
  AND4_X1   g0247(.A1(new_n439), .A2(new_n445), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n444), .A2(new_n415), .B1(new_n323), .B2(new_n411), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n439), .B1(new_n449), .B2(new_n446), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n436), .A2(new_n438), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n389), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g0254(.A(G97), .B(G107), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT6), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n456), .A2(new_n205), .A3(G107), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n460), .A2(G20), .B1(G77), .B2(new_n424), .ZN(new_n461));
  OAI21_X1  g0261(.A(G107), .B1(new_n417), .B2(new_n419), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n258), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(KEYINPUT79), .B1(new_n253), .B2(G1), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT79), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(new_n260), .A3(G33), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n262), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G97), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n261), .A2(G97), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n470), .B(KEYINPUT78), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT80), .B1(new_n463), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n472), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n458), .B1(new_n456), .B2(new_n455), .ZN(new_n475));
  OAI22_X1  g0275(.A1(new_n475), .A2(new_n226), .B1(new_n287), .B2(new_n254), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n206), .B1(new_n440), .B2(new_n441), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n257), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT80), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n474), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n301), .A2(new_n303), .A3(G244), .A4(new_n285), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT4), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n284), .A2(KEYINPUT4), .A3(G244), .A4(new_n285), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n284), .A2(G250), .A3(G1698), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G283), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n483), .A2(new_n484), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT5), .B(G41), .ZN(new_n488));
  INV_X1    g0288(.A(G45), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(G1), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n488), .A2(new_n490), .B1(new_n272), .B2(new_n273), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n487), .A2(new_n283), .B1(G257), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  NOR2_X1   g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(G274), .B1(new_n282), .B2(new_n225), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n492), .A2(new_n354), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(G200), .B1(new_n492), .B2(new_n498), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n473), .B(new_n480), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n474), .A2(new_n478), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n492), .A2(G179), .A3(new_n498), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n323), .B1(new_n492), .B2(new_n498), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n260), .A2(G45), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G250), .ZN(new_n507));
  OAI22_X1  g0307(.A1(new_n496), .A2(new_n506), .B1(new_n283), .B2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n301), .A2(new_n303), .A3(G238), .A4(new_n285), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n301), .A2(new_n303), .A3(G244), .A4(G1698), .ZN(new_n510));
  INV_X1    g0310(.A(G116), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n509), .B(new_n510), .C1(new_n253), .C2(new_n511), .ZN(new_n512));
  AOI211_X1 g0312(.A(new_n354), .B(new_n508), .C1(new_n283), .C2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n284), .A2(new_n226), .A3(G68), .ZN(new_n514));
  NAND3_X1  g0314(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n226), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(G87), .B2(new_n207), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT19), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n251), .B2(new_n205), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n514), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n257), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n376), .A2(new_n373), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n468), .A2(G87), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n513), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n508), .B1(new_n512), .B2(new_n283), .ZN(new_n526));
  OR2_X1    g0326(.A1(new_n526), .A2(new_n293), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n512), .A2(new_n283), .ZN(new_n528));
  INV_X1    g0328(.A(new_n508), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(G179), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n323), .B2(new_n526), .ZN(new_n531));
  INV_X1    g0331(.A(new_n468), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n521), .B(new_n522), .C1(new_n532), .C2(new_n376), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n525), .A2(new_n527), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n501), .A2(new_n505), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT87), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT86), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n261), .A2(G107), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(KEYINPUT25), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT25), .ZN(new_n540));
  NOR4_X1   g0340(.A1(new_n261), .A2(KEYINPUT86), .A3(new_n540), .A4(G107), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n536), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n339), .A2(G20), .A3(new_n206), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT86), .B1(new_n543), .B2(new_n540), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n538), .A2(new_n537), .A3(KEYINPUT25), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(KEYINPUT87), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n543), .A2(new_n540), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n542), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n468), .A2(G107), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n301), .A2(new_n303), .A3(G257), .A4(G1698), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n301), .A2(new_n303), .A3(G250), .A4(new_n285), .ZN(new_n552));
  INV_X1    g0352(.A(G294), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n551), .B(new_n552), .C1(new_n253), .C2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n497), .B1(new_n554), .B2(new_n283), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n495), .A2(G264), .A3(new_n274), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT88), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n495), .A2(KEYINPUT88), .A3(G264), .A4(new_n274), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n293), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n555), .A2(new_n560), .A3(new_n354), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n301), .A2(new_n303), .A3(new_n226), .A4(G87), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT83), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n284), .A2(KEYINPUT83), .A3(new_n226), .A4(G87), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT22), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT84), .ZN(new_n569));
  INV_X1    g0369(.A(new_n564), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT22), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n566), .A2(new_n567), .A3(new_n569), .A4(KEYINPUT22), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n253), .A2(new_n511), .A3(G20), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT23), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n226), .B2(G107), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n573), .A2(new_n574), .A3(new_n579), .ZN(new_n580));
  XOR2_X1   g0380(.A(KEYINPUT85), .B(KEYINPUT24), .Z(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n258), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n573), .A2(new_n581), .A3(new_n574), .A4(new_n579), .ZN(new_n584));
  AOI221_X4 g0384(.A(new_n550), .B1(new_n562), .B2(new_n563), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n535), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n365), .A2(G303), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n301), .A2(new_n303), .A3(G264), .A4(G1698), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n301), .A2(new_n303), .A3(G257), .A4(new_n285), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT82), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n587), .A2(KEYINPUT82), .A3(new_n588), .A4(new_n589), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n283), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n491), .A2(KEYINPUT81), .A3(G270), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n495), .A2(G270), .A3(new_n274), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT81), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n497), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n595), .A2(new_n600), .A3(new_n403), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n274), .B1(new_n592), .B2(new_n593), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT81), .B1(new_n491), .B2(G270), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n597), .A2(new_n598), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n498), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(G200), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n261), .A2(G116), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n468), .B2(G116), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n486), .B(new_n226), .C1(G33), .C2(new_n205), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n511), .A2(G20), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(new_n257), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT20), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n609), .A2(new_n257), .A3(KEYINPUT20), .A4(new_n610), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n601), .A2(new_n606), .A3(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n616), .A2(new_n296), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n602), .A2(new_n605), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT21), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n595), .A2(new_n600), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n323), .B1(new_n608), .B2(new_n615), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n623), .B(new_n621), .C1(new_n602), .C2(new_n605), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n617), .B(new_n620), .C1(new_n624), .C2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n583), .A2(new_n584), .ZN(new_n628));
  INV_X1    g0428(.A(new_n550), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT89), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n323), .B1(new_n555), .B2(new_n560), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n555), .A2(new_n560), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n630), .A2(new_n631), .B1(new_n632), .B2(G179), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT89), .B1(new_n632), .B2(new_n323), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n628), .A2(new_n629), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n627), .A2(new_n635), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n454), .A2(new_n586), .A3(new_n636), .ZN(G372));
  INV_X1    g0437(.A(new_n534), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n638), .A2(new_n505), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n531), .A2(new_n533), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n503), .A2(new_n504), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n473), .A2(new_n480), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n647), .A2(KEYINPUT90), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n638), .B1(new_n647), .B2(KEYINPUT90), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(new_n640), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n620), .B1(new_n624), .B2(new_n626), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n586), .B1(new_n635), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n644), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n454), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n350), .B1(new_n361), .B2(new_n382), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n409), .A2(new_n412), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT77), .B1(new_n656), .B2(new_n445), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n413), .A2(new_n432), .A3(new_n433), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n437), .B1(new_n659), .B2(KEYINPUT17), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n451), .B1(new_n655), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n295), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n654), .A2(new_n298), .A3(new_n663), .ZN(G369));
  NAND2_X1  g0464(.A1(new_n339), .A2(new_n226), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n339), .A2(new_n667), .A3(new_n226), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(G213), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT91), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(new_n616), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n651), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n627), .B2(new_n672), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n628), .A2(new_n629), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n633), .A2(new_n634), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n671), .B1(new_n628), .B2(new_n629), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n678), .B1(new_n585), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n635), .A2(new_n671), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n675), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n651), .A2(new_n671), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n681), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n684), .A2(new_n688), .ZN(G399));
  INV_X1    g0489(.A(new_n222), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G1), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n230), .B2(new_n692), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n643), .B1(new_n639), .B2(new_n640), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n652), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n640), .B1(new_n648), .B2(new_n649), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n671), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT29), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n653), .A2(new_n671), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n702), .B1(KEYINPUT29), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  AOI211_X1 g0505(.A(new_n296), .B(new_n508), .C1(new_n283), .C2(new_n512), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n706), .A2(new_n492), .A3(new_n560), .A4(new_n555), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n705), .B1(new_n707), .B2(new_n622), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n487), .A2(new_n283), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n491), .A2(G257), .ZN(new_n710));
  AND4_X1   g0510(.A1(G179), .A2(new_n709), .A3(new_n710), .A4(new_n526), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n711), .A2(new_n619), .A3(KEYINPUT30), .A4(new_n632), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n492), .A2(new_n498), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n526), .A2(G179), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n622), .A2(new_n561), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n708), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT31), .B1(new_n716), .B2(new_n701), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n636), .A2(new_n586), .A3(new_n671), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G330), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT92), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n704), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n696), .B1(new_n724), .B2(G1), .ZN(G364));
  NOR2_X1   g0525(.A1(new_n674), .A2(G330), .ZN(new_n726));
  XOR2_X1   g0526(.A(new_n726), .B(KEYINPUT93), .Z(new_n727));
  NOR2_X1   g0527(.A1(new_n338), .A2(G20), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n260), .B1(new_n728), .B2(G45), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n691), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n727), .A2(new_n675), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(G20), .B1(KEYINPUT95), .B2(G169), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(KEYINPUT95), .A2(G169), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n225), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n226), .A2(new_n296), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G200), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n354), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G179), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G190), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  AOI22_X1  g0546(.A1(new_n743), .A2(G311), .B1(G294), .B2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(G326), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n740), .A2(new_n293), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n403), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n747), .B1(new_n748), .B2(new_n753), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT98), .Z(new_n755));
  NAND2_X1  g0555(.A1(new_n741), .A2(new_n403), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G322), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n744), .A2(G20), .A3(new_n354), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n284), .B1(new_n760), .B2(G329), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n750), .A2(G190), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  XOR2_X1   g0563(.A(KEYINPUT33), .B(G317), .Z(new_n764));
  OAI211_X1 g0564(.A(new_n758), .B(new_n761), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n296), .A2(G200), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n226), .B1(new_n766), .B2(KEYINPUT96), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(KEYINPUT96), .B2(new_n766), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(G190), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n765), .B1(G283), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G303), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n768), .A2(new_n354), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n772), .A2(KEYINPUT97), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(KEYINPUT97), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n755), .B(new_n770), .C1(new_n771), .C2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n775), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G87), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n760), .A2(G159), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT32), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n365), .B(new_n780), .C1(G68), .C2(new_n762), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n769), .A2(G107), .ZN(new_n782));
  INV_X1    g0582(.A(new_n746), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n753), .A2(new_n202), .B1(new_n205), .B2(new_n783), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n421), .A2(new_n756), .B1(new_n742), .B2(new_n287), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n778), .A2(new_n781), .A3(new_n782), .A4(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n738), .B1(new_n776), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G13), .A2(G33), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n737), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n690), .A2(new_n365), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT94), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n794), .A2(G355), .B1(new_n511), .B2(new_n690), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n248), .A2(G45), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n690), .A2(new_n284), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(G45), .B2(new_n230), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n795), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n732), .B(new_n788), .C1(new_n792), .C2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n791), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n674), .B2(new_n801), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n733), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(G396));
  NAND2_X1  g0604(.A1(new_n382), .A2(new_n671), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n386), .A2(new_n387), .B1(new_n379), .B2(new_n701), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n805), .B1(new_n806), .B2(new_n382), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n703), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n807), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n653), .A2(new_n671), .A3(new_n809), .ZN(new_n810));
  AND3_X1   g0610(.A1(new_n723), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n723), .B1(new_n808), .B2(new_n810), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n811), .A2(new_n812), .A3(new_n731), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n738), .A2(new_n790), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n731), .B1(new_n814), .B2(G77), .ZN(new_n815));
  INV_X1    g0615(.A(new_n769), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n346), .ZN(new_n817));
  INV_X1    g0617(.A(G132), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n284), .B1(new_n818), .B2(new_n759), .C1(new_n783), .C2(new_n421), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G137), .A2(new_n752), .B1(new_n743), .B2(G159), .ZN(new_n820));
  INV_X1    g0620(.A(G143), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n820), .B1(new_n821), .B2(new_n756), .C1(new_n252), .C2(new_n763), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT34), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n817), .B(new_n819), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n824), .B1(new_n823), .B2(new_n822), .C1(new_n202), .C2(new_n775), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G116), .A2(new_n743), .B1(new_n757), .B2(G294), .ZN(new_n826));
  XNOR2_X1  g0626(.A(KEYINPUT99), .B(G283), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n826), .B1(new_n771), .B2(new_n753), .C1(new_n763), .C2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n775), .A2(new_n206), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n769), .A2(G87), .ZN(new_n830));
  INV_X1    g0630(.A(G311), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n365), .B1(new_n831), .B2(new_n759), .C1(new_n783), .C2(new_n205), .ZN(new_n832));
  NOR4_X1   g0632(.A1(new_n828), .A2(new_n829), .A3(new_n830), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(KEYINPUT100), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n833), .A2(KEYINPUT100), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n825), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n815), .B1(new_n836), .B2(new_n737), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n809), .B2(new_n790), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT101), .Z(new_n839));
  NOR2_X1   g0639(.A1(new_n813), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G384));
  NOR2_X1   g0641(.A1(new_n728), .A2(new_n260), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT38), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n445), .A2(new_n670), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n660), .B2(new_n451), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n449), .A2(new_n446), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n657), .A2(new_n658), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT102), .B1(new_n445), .B2(new_n670), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT102), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT91), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n669), .B(new_n850), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n849), .B(new_n851), .C1(new_n444), .C2(new_n415), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n848), .A2(new_n852), .A3(KEYINPUT37), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n657), .A2(new_n658), .A3(new_n846), .A4(new_n844), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n847), .A2(new_n853), .B1(new_n854), .B2(KEYINPUT37), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n843), .B1(new_n845), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n844), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n452), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n854), .A2(KEYINPUT37), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n434), .A2(new_n435), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n860), .A2(new_n853), .A3(new_n846), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n858), .A2(new_n862), .A3(KEYINPUT38), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n856), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT39), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n848), .A2(new_n852), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n446), .A2(new_n449), .B1(new_n413), .B2(new_n432), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n867), .B1(new_n868), .B2(KEYINPUT103), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n413), .A2(new_n432), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n846), .A2(new_n870), .A3(KEYINPUT103), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT37), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n867), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n872), .A2(new_n861), .B1(new_n452), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n863), .B1(new_n874), .B2(KEYINPUT38), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n866), .B1(new_n865), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n351), .A2(new_n701), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n451), .A2(new_n670), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n810), .A2(new_n805), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n332), .A2(new_n337), .A3(new_n348), .ZN(new_n882));
  INV_X1    g0682(.A(new_n318), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT14), .B1(new_n324), .B2(KEYINPUT72), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n320), .A2(new_n321), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n359), .B1(new_n355), .B2(new_n357), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n882), .B(new_n701), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n701), .A2(new_n882), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n361), .B(new_n889), .C1(new_n326), .C2(new_n349), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n881), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n879), .B1(new_n893), .B2(new_n864), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n878), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n663), .A2(new_n298), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n454), .B2(new_n704), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n895), .B(new_n897), .Z(new_n898));
  INV_X1    g0698(.A(G330), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n454), .A2(new_n721), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n807), .B1(new_n888), .B2(new_n890), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n721), .A2(new_n901), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n858), .A2(new_n862), .A3(KEYINPUT38), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT38), .B1(new_n858), .B2(new_n862), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT40), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n721), .A2(new_n901), .A3(KEYINPUT40), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n872), .A2(new_n861), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n452), .A2(new_n873), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT38), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n908), .B1(new_n911), .B2(new_n903), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n899), .B1(new_n900), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n913), .B2(new_n900), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n842), .B1(new_n898), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n898), .B2(new_n915), .ZN(new_n917));
  AOI211_X1 g0717(.A(new_n511), .B(new_n228), .C1(new_n460), .C2(KEYINPUT35), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(KEYINPUT35), .B2(new_n460), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT36), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n230), .A2(new_n287), .A3(new_n422), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n346), .A2(G50), .ZN(new_n922));
  OAI211_X1 g0722(.A(G1), .B(new_n338), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n917), .A2(new_n920), .A3(new_n923), .ZN(G367));
  INV_X1    g0724(.A(KEYINPUT45), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n646), .A2(new_n701), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(new_n505), .A3(new_n501), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n645), .A2(new_n646), .A3(new_n701), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n688), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n930), .A2(KEYINPUT106), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(KEYINPUT106), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n925), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n930), .A2(KEYINPUT106), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n930), .A2(KEYINPUT106), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(KEYINPUT45), .A3(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT44), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n688), .B2(new_n929), .ZN(new_n938));
  INV_X1    g0738(.A(new_n929), .ZN(new_n939));
  OAI211_X1 g0739(.A(KEYINPUT44), .B(new_n939), .C1(new_n686), .C2(new_n687), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n933), .A2(new_n936), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(KEYINPUT107), .A3(new_n683), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n682), .B(new_n685), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(new_n675), .Z(new_n945));
  NAND2_X1  g0745(.A1(new_n724), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n933), .A2(new_n936), .A3(new_n684), .A4(new_n941), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n943), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT107), .B1(new_n942), .B2(new_n683), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n724), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n691), .B(KEYINPUT41), .Z(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n730), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n683), .A2(new_n929), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT105), .Z(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT104), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n686), .A2(new_n929), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(KEYINPUT42), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n505), .B1(new_n939), .B2(new_n678), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n671), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n958), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n960), .A2(new_n958), .A3(new_n962), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n964), .B(new_n965), .C1(KEYINPUT42), .C2(new_n959), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n701), .A2(new_n524), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n534), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n642), .B2(new_n967), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n957), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n966), .A2(new_n970), .A3(new_n957), .ZN(new_n974));
  AND3_X1   g0774(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n973), .B1(new_n972), .B2(new_n974), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(KEYINPUT108), .B1(new_n954), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT108), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n942), .A2(new_n683), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT107), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n983), .A2(new_n943), .A3(new_n947), .A4(new_n948), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n952), .B1(new_n984), .B2(new_n724), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n977), .B(new_n980), .C1(new_n985), .C2(new_n730), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n979), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n235), .A2(new_n797), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n376), .A2(new_n222), .ZN(new_n989));
  NOR3_X1   g0789(.A1(new_n989), .A2(new_n737), .A3(new_n791), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n732), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n783), .A2(new_n346), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n365), .B(new_n992), .C1(G137), .C2(new_n760), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n769), .A2(G77), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G143), .A2(new_n752), .B1(new_n743), .B2(G50), .ZN(new_n995));
  AOI22_X1  g0795(.A1(G159), .A2(new_n762), .B1(new_n757), .B2(G150), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n993), .A2(new_n994), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G58), .B2(new_n777), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n284), .B1(new_n760), .B2(G317), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n756), .B2(new_n771), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G311), .A2(new_n752), .B1(new_n762), .B2(G294), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n206), .B2(new_n783), .C1(new_n742), .C2(new_n827), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n1000), .B(new_n1002), .C1(G97), .C2(new_n769), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n777), .A2(G116), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT46), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n998), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT47), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n991), .B1(new_n801), .B2(new_n969), .C1(new_n1007), .C2(new_n738), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n987), .A2(new_n1008), .ZN(G387));
  NOR2_X1   g0809(.A1(new_n947), .A2(new_n692), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n724), .B2(new_n945), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(KEYINPUT109), .B(G322), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n752), .A2(new_n1012), .B1(new_n757), .B2(G317), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n771), .B2(new_n742), .C1(new_n831), .C2(new_n763), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT48), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1015), .B1(new_n553), .B2(new_n775), .C1(new_n783), .C2(new_n827), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT49), .Z(new_n1017));
  OAI221_X1 g0817(.A(new_n365), .B1(new_n748), .B2(new_n759), .C1(new_n816), .C2(new_n511), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT110), .Z(new_n1019));
  NOR2_X1   g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n783), .A2(new_n376), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n365), .B(new_n1021), .C1(G150), .C2(new_n760), .ZN(new_n1022));
  XOR2_X1   g0822(.A(KEYINPUT8), .B(G58), .Z(new_n1023));
  AOI22_X1  g0823(.A1(G159), .A2(new_n752), .B1(new_n762), .B2(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G50), .A2(new_n757), .B1(new_n743), .B2(G68), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1022), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n775), .A2(new_n287), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(G97), .C2(new_n769), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n737), .B1(new_n1020), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n241), .A2(G45), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n693), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n1030), .A2(new_n797), .B1(new_n1031), .B2(new_n794), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n693), .B(new_n489), .C1(new_n346), .C2(new_n287), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT50), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n1023), .B2(new_n202), .ZN(new_n1035));
  NOR3_X1   g0835(.A1(new_n250), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n1032), .A2(new_n1037), .B1(G107), .B2(new_n222), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n732), .B1(new_n1038), .B2(new_n792), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1029), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n682), .B2(new_n791), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n945), .B2(new_n730), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1011), .A2(new_n1042), .ZN(G393));
  INV_X1    g0843(.A(KEYINPUT113), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n981), .A2(KEYINPUT111), .A3(new_n948), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT111), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n942), .A2(new_n1046), .A3(new_n683), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1045), .A2(new_n946), .A3(new_n1047), .ZN(new_n1048));
  AND3_X1   g0848(.A1(new_n1048), .A2(new_n984), .A3(new_n691), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n730), .ZN(new_n1051));
  INV_X1    g0851(.A(G159), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n753), .A2(new_n252), .B1(new_n1052), .B2(new_n756), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT51), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n763), .A2(new_n202), .B1(new_n250), .B2(new_n742), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n783), .A2(new_n287), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n284), .B1(new_n759), .B2(new_n821), .ZN(new_n1057));
  NOR4_X1   g0857(.A1(new_n1055), .A2(new_n830), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1054), .B(new_n1058), .C1(new_n346), .C2(new_n775), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G317), .A2(new_n752), .B1(new_n757), .B2(G311), .ZN(new_n1060));
  XOR2_X1   g0860(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n1061));
  XNOR2_X1  g0861(.A(new_n1060), .B(new_n1061), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G303), .A2(new_n762), .B1(new_n743), .B2(G294), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n746), .A2(G116), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n284), .B1(new_n760), .B2(new_n1012), .ZN(new_n1065));
  AND4_X1   g0865(.A1(new_n782), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1062), .B(new_n1066), .C1(new_n775), .C2(new_n827), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n738), .B1(new_n1059), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n245), .A2(new_n797), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n791), .B(new_n737), .C1(G97), .C2(new_n690), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n732), .B(new_n1068), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n929), .B2(new_n801), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1051), .A2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1044), .B1(new_n1049), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1048), .A2(new_n984), .A3(new_n691), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1075), .A2(KEYINPUT113), .A3(new_n1051), .A4(new_n1072), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1074), .A2(new_n1076), .ZN(G390));
  OAI221_X1 g0877(.A(new_n671), .B1(new_n382), .B2(new_n806), .C1(new_n698), .C2(new_n699), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n805), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n891), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n877), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1080), .A2(new_n1081), .A3(new_n875), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n877), .B1(new_n880), .B2(new_n891), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1082), .B1(new_n876), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n899), .B1(new_n719), .B2(new_n720), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n901), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT114), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n723), .A2(new_n809), .A3(new_n891), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1082), .B(new_n1089), .C1(new_n876), .C2(new_n1083), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n892), .B1(new_n722), .B2(new_n807), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1089), .A2(new_n805), .A3(new_n1078), .A4(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n723), .A2(new_n809), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1087), .B1(new_n1095), .B2(new_n892), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1094), .B1(new_n1096), .B2(new_n881), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n454), .A2(new_n1085), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n897), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(KEYINPUT115), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n692), .B1(new_n1092), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n1092), .B2(new_n1101), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1092), .A2(new_n730), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n731), .B1(new_n814), .B2(new_n1023), .ZN(new_n1105));
  INV_X1    g0905(.A(G283), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n206), .A2(new_n763), .B1(new_n753), .B2(new_n1106), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n205), .A2(new_n742), .B1(new_n756), .B2(new_n511), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n769), .A2(G68), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n284), .B(new_n1056), .C1(G294), .C2(new_n760), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n778), .A2(new_n1109), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  XOR2_X1   g0912(.A(KEYINPUT54), .B(G143), .Z(new_n1113));
  AOI22_X1  g0913(.A1(new_n762), .A2(G137), .B1(new_n743), .B2(new_n1113), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1114), .B1(new_n818), .B2(new_n756), .C1(new_n1052), .C2(new_n783), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n365), .B1(new_n760), .B2(G125), .ZN(new_n1116));
  INV_X1    g0916(.A(G128), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1116), .B1(new_n753), .B2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(KEYINPUT53), .B1(new_n775), .B2(new_n252), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1119), .B(new_n1120), .C1(new_n202), .C2(new_n816), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n775), .A2(KEYINPUT53), .A3(new_n252), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1112), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1105), .B1(new_n1123), .B2(new_n737), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n876), .B2(new_n790), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1103), .A2(new_n1104), .A3(new_n1125), .ZN(G378));
  INV_X1    g0926(.A(KEYINPUT120), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n267), .A2(new_n851), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n295), .A2(new_n298), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1131), .B1(new_n295), .B2(new_n298), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1129), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n299), .A2(new_n1130), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1136), .A2(new_n1132), .A3(new_n1128), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n899), .B1(new_n875), .B2(new_n908), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n907), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(KEYINPUT119), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n907), .A2(new_n1139), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT118), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1138), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n907), .A2(new_n1139), .A3(KEYINPUT118), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1141), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT119), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n912), .A2(G330), .ZN(new_n1148));
  AOI21_X1  g0948(.A(KEYINPUT40), .B1(new_n864), .B2(new_n902), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1143), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1138), .ZN(new_n1151));
  AND4_X1   g0951(.A1(new_n1147), .A2(new_n1150), .A3(new_n1145), .A4(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1127), .B1(new_n1146), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1150), .A2(new_n1145), .A3(new_n1151), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1140), .A2(KEYINPUT119), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1144), .A2(new_n1147), .A3(new_n1145), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1156), .A2(KEYINPUT120), .A3(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1153), .A2(new_n895), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT121), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n895), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1159), .A2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1153), .A2(new_n1160), .A3(new_n895), .A4(new_n1158), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1099), .A2(KEYINPUT122), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1088), .A2(new_n1097), .A3(new_n1090), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1099), .A2(KEYINPUT122), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1166), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1164), .A2(new_n1165), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT57), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1169), .A2(KEYINPUT57), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT123), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1161), .A2(KEYINPUT123), .A3(new_n1162), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1156), .A2(new_n895), .A3(new_n1157), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n692), .B1(new_n1173), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1172), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1164), .A2(new_n1165), .A3(new_n730), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n731), .B1(new_n814), .B2(G50), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G125), .A2(new_n752), .B1(new_n762), .B2(G132), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G128), .A2(new_n757), .B1(new_n743), .B2(G137), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(new_n252), .C2(new_n783), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n777), .B2(new_n1113), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(G33), .A2(G41), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT116), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n816), .A2(new_n1052), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(G124), .C2(new_n760), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1189), .A2(new_n1190), .A3(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n816), .A2(new_n421), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT117), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(G116), .A2(new_n752), .B1(new_n757), .B2(G107), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n205), .B2(new_n763), .C1(new_n376), .C2(new_n742), .ZN(new_n1200));
  AOI211_X1 g1000(.A(G41), .B(new_n284), .C1(new_n760), .C2(G283), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n346), .B2(new_n783), .ZN(new_n1202));
  NOR4_X1   g1002(.A1(new_n1198), .A2(new_n1200), .A3(new_n1027), .A4(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(KEYINPUT58), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1203), .A2(KEYINPUT58), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1192), .B(new_n202), .C1(G41), .C2(new_n284), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1195), .A2(new_n1204), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1183), .B1(new_n1207), .B2(new_n737), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n1138), .B2(new_n790), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1182), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1181), .A2(new_n1210), .ZN(G375));
  OR2_X1    g1011(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1212), .A2(new_n953), .A3(new_n1100), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n892), .A2(new_n789), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n731), .B1(new_n814), .B2(G68), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n284), .B1(new_n759), .B2(new_n1117), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(G132), .A2(new_n752), .B1(new_n762), .B2(new_n1113), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n202), .B2(new_n783), .C1(new_n252), .C2(new_n742), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1216), .B(new_n1218), .C1(G137), .C2(new_n757), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1219), .B(new_n1197), .C1(new_n1052), .C2(new_n775), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n763), .A2(new_n511), .B1(new_n1106), .B2(new_n756), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n753), .A2(new_n553), .B1(new_n206), .B2(new_n742), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n759), .A2(new_n771), .ZN(new_n1223));
  NOR4_X1   g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1021), .A4(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n205), .B2(new_n775), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n994), .A2(new_n365), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT124), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1220), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1215), .B1(new_n1228), .B2(new_n737), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1097), .A2(new_n730), .B1(new_n1214), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1213), .A2(new_n1230), .ZN(G381));
  INV_X1    g1031(.A(G390), .ZN(new_n1232));
  INV_X1    g1032(.A(G378), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  OR3_X1    g1035(.A1(new_n1235), .A2(G375), .A3(G387), .ZN(G407));
  INV_X1    g1036(.A(G343), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(G213), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(KEYINPUT125), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1233), .A2(new_n1239), .ZN(new_n1240));
  OAI211_X1 g1040(.A(G407), .B(G213), .C1(G375), .C2(new_n1240), .ZN(G409));
  INV_X1    g1041(.A(KEYINPUT61), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1181), .A2(G378), .A3(new_n1210), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1179), .A2(new_n730), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1244), .B(new_n1209), .C1(new_n1170), .C2(new_n952), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1233), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1239), .B1(new_n1243), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1100), .A2(KEYINPUT60), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1248), .A2(new_n1212), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n691), .B1(new_n1248), .B2(new_n1212), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1230), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n840), .ZN(new_n1252));
  OAI211_X1 g1052(.A(G384), .B(new_n1230), .C1(new_n1249), .C2(new_n1250), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1252), .A2(new_n1253), .B1(G2897), .B2(new_n1239), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1238), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1257), .A2(G2897), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1254), .B1(new_n1256), .B2(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1242), .B1(new_n1247), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT126), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1256), .A2(KEYINPUT62), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1247), .A2(new_n1262), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n1257), .B(new_n1255), .C1(new_n1243), .C2(new_n1246), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1263), .B1(new_n1264), .B2(KEYINPUT62), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT126), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1266), .B(new_n1242), .C1(new_n1247), .C2(new_n1259), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1261), .A2(new_n1265), .A3(new_n1267), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(G393), .B(new_n803), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n987), .A2(G390), .A3(new_n1008), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(G390), .B1(new_n987), .B2(new_n1008), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1270), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(G387), .A2(new_n1232), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(new_n1269), .A3(new_n1271), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1268), .A2(new_n1277), .ZN(new_n1278));
  OR2_X1    g1078(.A1(new_n1264), .A2(KEYINPUT63), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1277), .A2(KEYINPUT61), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1247), .A2(KEYINPUT63), .A3(new_n1256), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1243), .A2(new_n1246), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1256), .A2(new_n1258), .ZN(new_n1283));
  OAI22_X1  g1083(.A1(new_n1282), .A2(new_n1257), .B1(new_n1254), .B2(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .A4(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1278), .A2(new_n1285), .ZN(G405));
  NOR2_X1   g1086(.A1(new_n1256), .A2(KEYINPUT127), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1272), .A2(new_n1273), .A3(new_n1270), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1269), .B1(new_n1275), .B2(new_n1271), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1287), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1274), .B(new_n1276), .C1(KEYINPUT127), .C2(new_n1256), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT127), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1243), .B1(new_n1293), .B2(new_n1255), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1294), .B1(new_n1233), .B2(G375), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1292), .B(new_n1295), .ZN(G402));
endmodule


