//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1241, new_n1242, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(KEYINPUT67), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n217), .A2(KEYINPUT67), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n211), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  INV_X1    g0024(.A(new_n206), .ZN(new_n225));
  OR2_X1    g0025(.A1(new_n225), .A2(KEYINPUT66), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(KEYINPUT66), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n226), .A2(G50), .A3(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(KEYINPUT65), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n234), .B1(new_n211), .B2(G13), .ZN(new_n235));
  INV_X1    g0035(.A(G13), .ZN(new_n236));
  NAND4_X1  g0036(.A1(new_n236), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g0038(.A(new_n238), .B(G250), .C1(G257), .C2(G264), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT0), .ZN(new_n240));
  NAND3_X1  g0040(.A1(new_n224), .A2(new_n233), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g0041(.A(new_n241), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G232), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT2), .B(G226), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G250), .B(G257), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G264), .B(G270), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G358));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT68), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G50), .B(G68), .ZN(new_n255));
  XNOR2_X1  g0055(.A(G58), .B(G77), .ZN(new_n256));
  XOR2_X1   g0056(.A(new_n255), .B(new_n256), .Z(new_n257));
  XNOR2_X1  g0057(.A(new_n254), .B(new_n257), .ZN(G351));
  INV_X1    g0058(.A(KEYINPUT9), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n208), .A2(KEYINPUT73), .A3(G20), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT73), .ZN(new_n261));
  AOI21_X1  g0061(.A(G50), .B1(new_n204), .B2(new_n205), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n261), .B1(new_n262), .B2(new_n231), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G20), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G150), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT8), .ZN(new_n266));
  NOR3_X1   g0066(.A1(new_n266), .A2(KEYINPUT72), .A3(G58), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(G58), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(new_n270), .A3(KEYINPUT72), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n268), .A2(new_n271), .A3(new_n231), .A4(G33), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n260), .A2(new_n263), .A3(new_n265), .A4(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT71), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g0076(.A1(KEYINPUT71), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(new_n230), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  NOR3_X1   g0079(.A1(new_n236), .A2(new_n231), .A3(G1), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n207), .ZN(new_n281));
  INV_X1    g0081(.A(G1), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G20), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n276), .A2(new_n230), .A3(new_n277), .A4(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n281), .B1(new_n284), .B2(new_n207), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n259), .B1(new_n279), .B2(new_n286), .ZN(new_n287));
  AOI211_X1 g0087(.A(KEYINPUT9), .B(new_n285), .C1(new_n273), .C2(new_n278), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT74), .ZN(new_n289));
  OR3_X1    g0089(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT3), .ZN(new_n291));
  INV_X1    g0091(.A(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(KEYINPUT3), .A2(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(G222), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(G223), .A3(G1698), .ZN(new_n298));
  AND2_X1   g0098(.A1(KEYINPUT3), .A2(G33), .ZN(new_n299));
  NOR2_X1   g0099(.A1(KEYINPUT3), .A2(G33), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G77), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n297), .A2(new_n298), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G41), .ZN(new_n306));
  OAI211_X1 g0106(.A(G1), .B(G13), .C1(new_n292), .C2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n282), .B1(G41), .B2(G45), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G45), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT69), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT69), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G45), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n311), .A2(new_n313), .A3(new_n306), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n282), .A2(G274), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n309), .A2(G226), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n305), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT70), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n305), .A2(new_n316), .A3(KEYINPUT70), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n319), .A2(KEYINPUT75), .A3(G200), .A4(new_n320), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n305), .A2(new_n316), .A3(KEYINPUT70), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT70), .B1(new_n305), .B2(new_n316), .ZN(new_n323));
  OAI21_X1  g0123(.A(G190), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT10), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n321), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n319), .A2(G200), .A3(new_n320), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT75), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n289), .B1(new_n287), .B2(new_n288), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n290), .A2(new_n326), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n324), .B(new_n327), .C1(new_n287), .C2(new_n288), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT76), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n332), .A2(new_n333), .A3(KEYINPUT10), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n333), .B1(new_n332), .B2(KEYINPUT10), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n331), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n293), .A2(new_n231), .A3(new_n294), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT7), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT7), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n293), .A2(new_n339), .A3(new_n231), .A4(new_n294), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(G68), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G58), .A2(G68), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n204), .A2(new_n205), .A3(new_n342), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n343), .A2(G20), .B1(G159), .B2(new_n264), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT16), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n341), .A2(KEYINPUT16), .A3(new_n344), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(new_n278), .A3(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n278), .A2(new_n280), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n268), .A2(new_n271), .A3(KEYINPUT80), .A4(new_n283), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT8), .B(G58), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n267), .B1(new_n353), .B2(KEYINPUT72), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT80), .B1(new_n354), .B2(new_n283), .ZN(new_n355));
  INV_X1    g0155(.A(new_n280), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n352), .A2(new_n355), .B1(new_n356), .B2(new_n354), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n349), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT82), .ZN(new_n360));
  OR2_X1    g0160(.A1(G223), .A2(G1698), .ZN(new_n361));
  INV_X1    g0161(.A(G226), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G1698), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n361), .B(new_n363), .C1(new_n299), .C2(new_n300), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n292), .A2(new_n213), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n307), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT81), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI211_X1 g0169(.A(KEYINPUT81), .B(new_n307), .C1(new_n364), .C2(new_n366), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n314), .A2(new_n315), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n307), .A2(G232), .A3(new_n308), .ZN(new_n372));
  INV_X1    g0172(.A(G179), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n369), .A2(new_n370), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G169), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n371), .A2(new_n372), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(new_n367), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n360), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n374), .ZN(new_n381));
  NOR2_X1   g0181(.A1(G223), .A2(G1698), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n362), .B2(G1698), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n365), .B1(new_n383), .B2(new_n295), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT81), .B1(new_n384), .B2(new_n307), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n364), .A2(new_n366), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(new_n368), .A3(new_n304), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n381), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n388), .A2(KEYINPUT82), .A3(new_n378), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n359), .A2(new_n380), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT18), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT18), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n359), .A2(new_n380), .A3(new_n392), .A4(new_n389), .ZN(new_n393));
  INV_X1    g0193(.A(G190), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n371), .A2(new_n372), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n385), .A2(new_n395), .A3(new_n387), .ZN(new_n396));
  INV_X1    g0196(.A(G200), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n377), .B2(new_n367), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n349), .A2(new_n399), .A3(new_n358), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT17), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n349), .A2(new_n358), .A3(new_n399), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT17), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n391), .A2(new_n393), .A3(new_n402), .A4(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n353), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n406), .A2(new_n264), .B1(G20), .B2(G77), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n231), .A2(G33), .ZN(new_n408));
  XNOR2_X1  g0208(.A(KEYINPUT15), .B(G87), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(G77), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n410), .A2(new_n278), .B1(new_n411), .B2(new_n280), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n276), .A2(new_n230), .A3(new_n277), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(G77), .A3(new_n283), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n309), .A2(G244), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n371), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n295), .A2(G232), .A3(new_n296), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n295), .A2(G238), .A3(G1698), .ZN(new_n420));
  INV_X1    g0220(.A(G107), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n419), .B(new_n420), .C1(new_n421), .C2(new_n295), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n418), .B1(new_n304), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G190), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n416), .B(new_n424), .C1(new_n397), .C2(new_n423), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n373), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n415), .B(new_n426), .C1(G169), .C2(new_n423), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n405), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n373), .B1(new_n322), .B2(new_n323), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n319), .A2(new_n376), .A3(new_n320), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n279), .A2(new_n286), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n295), .A2(G232), .A3(G1698), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n295), .A2(G226), .A3(new_n296), .ZN(new_n435));
  NAND2_X1  g0235(.A1(G33), .A2(G97), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n304), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n309), .A2(G238), .B1(new_n314), .B2(new_n315), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT13), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n440), .B1(new_n438), .B2(new_n439), .ZN(new_n443));
  OAI21_X1  g0243(.A(G200), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n443), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n445), .A2(G190), .A3(new_n441), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n350), .A2(G68), .A3(new_n283), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT78), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT12), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n203), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI22_X1  g0250(.A1(new_n356), .A2(new_n450), .B1(KEYINPUT78), .B2(KEYINPUT12), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n280), .A2(new_n448), .A3(new_n449), .A4(new_n203), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n447), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT77), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n264), .A2(new_n455), .A3(G50), .ZN(new_n456));
  OAI221_X1 g0256(.A(new_n456), .B1(new_n231), .B2(G68), .C1(new_n411), .C2(new_n408), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n455), .B1(new_n264), .B2(G50), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n278), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n459), .A2(KEYINPUT11), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(KEYINPUT11), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n454), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n444), .A2(new_n446), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(KEYINPUT79), .A2(KEYINPUT14), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n442), .A2(new_n443), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n465), .B1(new_n466), .B2(new_n376), .ZN(new_n467));
  OAI211_X1 g0267(.A(G169), .B(new_n464), .C1(new_n442), .C2(new_n443), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(G179), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n462), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n463), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND4_X1   g0272(.A1(new_n336), .A2(new_n429), .A3(new_n433), .A4(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT21), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n356), .A2(G116), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n282), .A2(G33), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n413), .A2(new_n356), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G116), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(G20), .B1(new_n292), .B2(G97), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G283), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT86), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n479), .A2(G20), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n278), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n484), .B1(new_n278), .B2(new_n485), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n483), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT20), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n278), .A2(new_n485), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT86), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n486), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n494), .A2(KEYINPUT20), .A3(new_n483), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n480), .B1(new_n491), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n295), .A2(G264), .A3(G1698), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n295), .A2(G257), .A3(new_n296), .ZN(new_n498));
  INV_X1    g0298(.A(G303), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n497), .B(new_n498), .C1(new_n499), .C2(new_n295), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n304), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n310), .A2(G1), .ZN(new_n502));
  AND2_X1   g0302(.A1(KEYINPUT5), .A2(G41), .ZN(new_n503));
  NOR2_X1   g0303(.A1(KEYINPUT5), .A2(G41), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(G270), .A3(new_n307), .ZN(new_n506));
  XNOR2_X1  g0306(.A(KEYINPUT5), .B(G41), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n507), .A2(new_n307), .A3(G274), .A4(new_n502), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT85), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT85), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n501), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G169), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n474), .B1(new_n496), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n480), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT20), .B1(new_n494), .B2(new_n483), .ZN(new_n515));
  INV_X1    g0315(.A(new_n483), .ZN(new_n516));
  AOI211_X1 g0316(.A(new_n490), .B(new_n516), .C1(new_n493), .C2(new_n486), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n514), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  OR2_X1    g0318(.A1(new_n510), .A2(new_n509), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n376), .B1(new_n519), .B2(new_n501), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n520), .A3(KEYINPUT21), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n501), .B(G179), .C1(new_n509), .C2(new_n510), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n513), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n519), .A2(G190), .A3(new_n501), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n511), .A2(G200), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n496), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT87), .ZN(new_n530));
  XNOR2_X1  g0330(.A(new_n529), .B(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(G238), .B(new_n296), .C1(new_n299), .C2(new_n300), .ZN(new_n532));
  OAI211_X1 g0332(.A(G244), .B(G1698), .C1(new_n299), .C2(new_n300), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G116), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n304), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n502), .A2(G274), .ZN(new_n537));
  OAI21_X1  g0337(.A(G250), .B1(new_n310), .B2(G1), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n304), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G200), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT19), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n231), .B1(new_n436), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(G97), .A2(G107), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n213), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n231), .B(G68), .C1(new_n299), .C2(new_n300), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n543), .B1(new_n408), .B2(new_n215), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n278), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n413), .A2(G87), .A3(new_n356), .A4(new_n477), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n409), .A2(new_n280), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n539), .B1(new_n535), .B2(new_n304), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G190), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n542), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n373), .ZN(new_n558));
  INV_X1    g0358(.A(new_n409), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n413), .A2(new_n356), .A3(new_n477), .A4(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n551), .A2(new_n560), .A3(new_n553), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n558), .B(new_n561), .C1(G169), .C2(new_n555), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT84), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n295), .A2(G250), .A3(new_n296), .ZN(new_n565));
  OAI211_X1 g0365(.A(G257), .B(G1698), .C1(new_n299), .C2(new_n300), .ZN(new_n566));
  NAND2_X1  g0366(.A1(G33), .A2(G294), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n304), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n304), .B1(new_n502), .B2(new_n507), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G264), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n508), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n376), .ZN(new_n573));
  AOI21_X1  g0373(.A(G20), .B1(new_n293), .B2(new_n294), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n574), .A2(KEYINPUT88), .A3(KEYINPUT22), .A4(G87), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n231), .B(G87), .C1(new_n299), .C2(new_n300), .ZN(new_n576));
  OR2_X1    g0376(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n577));
  NAND2_X1  g0377(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n534), .A2(G20), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT23), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n231), .B2(G107), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n421), .A2(KEYINPUT23), .A3(G20), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n580), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n575), .A2(new_n579), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT24), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT24), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n575), .A2(new_n579), .A3(new_n587), .A4(new_n584), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n413), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n280), .A2(new_n421), .ZN(new_n590));
  XOR2_X1   g0390(.A(new_n590), .B(KEYINPUT25), .Z(new_n591));
  NAND3_X1  g0391(.A1(new_n350), .A2(G107), .A3(new_n477), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI221_X1 g0393(.A(new_n573), .B1(G179), .B2(new_n572), .C1(new_n589), .C2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT84), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n557), .A2(new_n562), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n564), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n505), .A2(new_n307), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n508), .B1(new_n598), .B2(new_n216), .ZN(new_n599));
  OAI211_X1 g0399(.A(G244), .B(new_n296), .C1(new_n299), .C2(new_n300), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT4), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n295), .A2(KEYINPUT4), .A3(G244), .A4(new_n296), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n295), .A2(G250), .A3(G1698), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n602), .A2(new_n603), .A3(new_n482), .A4(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n599), .B1(new_n605), .B2(new_n304), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G190), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT6), .ZN(new_n608));
  AND2_X1   g0408(.A1(G97), .A2(G107), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n608), .B1(new_n609), .B2(new_n545), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n421), .A2(KEYINPUT6), .A3(G97), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n612), .A2(G20), .B1(G77), .B2(new_n264), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n338), .A2(G107), .A3(new_n340), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n413), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n356), .A2(G97), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n478), .B2(new_n215), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(G200), .B1(new_n606), .B2(KEYINPUT83), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT83), .ZN(new_n621));
  AOI211_X1 g0421(.A(new_n621), .B(new_n599), .C1(new_n304), .C2(new_n605), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n607), .B(new_n619), .C1(new_n620), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n605), .A2(new_n304), .ZN(new_n624));
  INV_X1    g0424(.A(new_n599), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n376), .ZN(new_n627));
  OR2_X1    g0427(.A1(new_n615), .A2(new_n618), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n606), .A2(new_n373), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n586), .A2(new_n588), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n278), .ZN(new_n632));
  INV_X1    g0432(.A(new_n593), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n568), .A2(new_n304), .B1(G264), .B2(new_n570), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(G190), .A3(new_n508), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n572), .A2(G200), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n632), .A2(new_n633), .A3(new_n635), .A4(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n623), .A2(new_n630), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n597), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n473), .A2(new_n526), .A3(new_n531), .A4(new_n639), .ZN(new_n640));
  XOR2_X1   g0440(.A(new_n640), .B(KEYINPUT89), .Z(G372));
  NAND4_X1  g0441(.A1(new_n513), .A2(new_n521), .A3(new_n594), .A4(new_n524), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n623), .A2(new_n630), .A3(new_n637), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n554), .A2(new_n556), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT90), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n535), .A2(new_n645), .A3(new_n304), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n645), .B1(new_n535), .B2(new_n304), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n540), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n644), .B1(G200), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n536), .A2(KEYINPUT90), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n535), .A2(new_n645), .A3(new_n304), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n539), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT91), .B1(new_n652), .B2(G169), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT91), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n648), .A2(new_n654), .A3(new_n376), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n558), .A2(new_n561), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n649), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n642), .A2(new_n643), .A3(new_n659), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n652), .A2(KEYINPUT91), .A3(G169), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n654), .B1(new_n648), .B2(new_n376), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n658), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT92), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n627), .A2(new_n628), .A3(new_n664), .A4(new_n629), .ZN(new_n665));
  OAI22_X1  g0465(.A1(new_n606), .A2(G169), .B1(new_n615), .B2(new_n618), .ZN(new_n666));
  AOI211_X1 g0466(.A(G179), .B(new_n599), .C1(new_n304), .C2(new_n605), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT92), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(KEYINPUT26), .B1(new_n669), .B2(new_n659), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n557), .A2(new_n562), .A3(new_n595), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n595), .B1(new_n557), .B2(new_n562), .ZN(new_n672));
  XOR2_X1   g0472(.A(KEYINPUT93), .B(KEYINPUT26), .Z(new_n673));
  NOR4_X1   g0473(.A1(new_n671), .A2(new_n672), .A3(new_n630), .A4(new_n673), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n660), .B(new_n663), .C1(new_n670), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n473), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n433), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n391), .A2(new_n393), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n463), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n404), .A2(new_n680), .A3(new_n402), .ZN(new_n681));
  INV_X1    g0481(.A(new_n427), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n470), .B2(new_n471), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n679), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n677), .B1(new_n684), .B2(new_n336), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n676), .A2(new_n685), .ZN(G369));
  NOR2_X1   g0486(.A1(new_n236), .A2(G20), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n282), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT94), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G213), .A3(new_n691), .ZN(new_n692));
  XOR2_X1   g0492(.A(KEYINPUT95), .B(G343), .Z(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n531), .B(new_n526), .C1(new_n496), .C2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n525), .A2(new_n518), .A3(new_n694), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n589), .A2(new_n593), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n637), .B1(new_n695), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n594), .ZN(new_n702));
  INV_X1    g0502(.A(new_n594), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n695), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n525), .A2(new_n695), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT96), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT96), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n525), .A2(new_n710), .A3(new_n695), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n705), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n707), .A2(new_n704), .A3(new_n714), .ZN(G399));
  INV_X1    g0515(.A(new_n238), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G41), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n546), .A2(G116), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(G1), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n228), .B2(new_n718), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT28), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT29), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n675), .A2(new_n723), .A3(new_n695), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n657), .B1(new_n653), .B2(new_n655), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n638), .A2(new_n649), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(new_n642), .ZN(new_n727));
  INV_X1    g0527(.A(new_n649), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n663), .A2(new_n728), .A3(new_n668), .A4(new_n665), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT26), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n671), .A2(new_n672), .A3(new_n630), .ZN(new_n731));
  INV_X1    g0531(.A(new_n673), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n729), .A2(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n694), .B1(new_n727), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n724), .B1(new_n734), .B2(new_n723), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G330), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n639), .A2(new_n531), .A3(new_n526), .A4(new_n695), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n606), .A2(new_n634), .A3(new_n555), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(new_n523), .A3(KEYINPUT30), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n624), .A2(new_n625), .B1(new_n634), .B2(new_n508), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(new_n373), .A3(new_n511), .A4(new_n648), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT30), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(new_n739), .B2(new_n522), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n741), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n694), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(KEYINPUT31), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT31), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n746), .A2(new_n749), .A3(new_n694), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n737), .B1(new_n738), .B2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n736), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n722), .B1(new_n755), .B2(G1), .ZN(G364));
  AOI21_X1  g0556(.A(new_n230), .B1(G20), .B2(new_n376), .ZN(new_n757));
  XOR2_X1   g0557(.A(KEYINPUT33), .B(G317), .Z(new_n758));
  NOR2_X1   g0558(.A1(new_n373), .A2(new_n397), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n231), .A2(G190), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n373), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(new_n760), .ZN(new_n763));
  INV_X1    g0563(.A(G311), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n758), .A2(new_n761), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n231), .A2(new_n394), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n759), .A2(new_n766), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n295), .B(new_n765), .C1(G326), .C2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n397), .A2(G179), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n766), .A2(new_n762), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(G303), .A2(new_n771), .B1(new_n773), .B2(G322), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n760), .A2(new_n769), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G179), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n760), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(G283), .A2(new_n776), .B1(new_n779), .B2(G329), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n777), .A2(G190), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G294), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n768), .A2(new_n774), .A3(new_n780), .A4(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT100), .ZN(new_n785));
  INV_X1    g0585(.A(new_n763), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G58), .A2(new_n773), .B1(new_n786), .B2(G77), .ZN(new_n787));
  INV_X1    g0587(.A(new_n767), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n207), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT98), .ZN(new_n790));
  INV_X1    g0590(.A(new_n782), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n215), .ZN(new_n792));
  INV_X1    g0592(.A(new_n761), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n792), .B1(G68), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT99), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n779), .A2(G159), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT32), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n775), .A2(new_n421), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n770), .A2(new_n213), .ZN(new_n799));
  NOR4_X1   g0599(.A1(new_n797), .A2(new_n301), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  AND3_X1   g0600(.A1(new_n790), .A2(new_n795), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n757), .B1(new_n785), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n282), .B1(new_n687), .B2(G45), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n717), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n238), .A2(new_n295), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT97), .Z(new_n808));
  AOI22_X1  g0608(.A1(new_n808), .A2(G355), .B1(new_n479), .B2(new_n716), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n716), .A2(new_n295), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n311), .A2(new_n313), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n810), .B1(new_n257), .B2(new_n310), .C1(new_n228), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(G13), .A2(G33), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(G20), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n757), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n806), .B1(new_n814), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n817), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n802), .B(new_n819), .C1(new_n698), .C2(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT101), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n698), .A2(G330), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n699), .A2(new_n806), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(G396));
  NAND2_X1  g0625(.A1(new_n682), .A2(new_n695), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n694), .A2(new_n415), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n425), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n827), .B1(new_n427), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n675), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n831), .B1(new_n832), .B2(new_n694), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n660), .A2(new_n663), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n729), .A2(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n695), .B(new_n830), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n805), .B1(new_n837), .B2(new_n753), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n753), .B2(new_n837), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G150), .A2(new_n793), .B1(new_n767), .B2(G137), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT102), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G143), .A2(new_n773), .B1(new_n786), .B2(G159), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT34), .Z(new_n844));
  NOR2_X1   g0644(.A1(new_n791), .A2(new_n202), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n295), .B1(new_n770), .B2(new_n207), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n776), .A2(G68), .ZN(new_n847));
  INV_X1    g0647(.A(G132), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n847), .B1(new_n848), .B2(new_n778), .ZN(new_n849));
  NOR4_X1   g0649(.A1(new_n844), .A2(new_n845), .A3(new_n846), .A4(new_n849), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n767), .A2(G303), .B1(new_n779), .B2(G311), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n851), .B(new_n301), .C1(new_n421), .C2(new_n770), .ZN(new_n852));
  INV_X1    g0652(.A(G283), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n761), .A2(new_n853), .B1(new_n763), .B2(new_n479), .ZN(new_n854));
  INV_X1    g0654(.A(G294), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n772), .A2(new_n855), .B1(new_n775), .B2(new_n213), .ZN(new_n856));
  NOR4_X1   g0656(.A1(new_n852), .A2(new_n792), .A3(new_n854), .A4(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n757), .B1(new_n850), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n757), .A2(new_n815), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n806), .B1(new_n411), .B2(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n858), .B(new_n860), .C1(new_n816), .C2(new_n830), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n839), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(G384));
  NAND2_X1  g0663(.A1(new_n738), .A2(new_n751), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n695), .A2(new_n462), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n472), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n470), .A2(new_n865), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n864), .A2(new_n830), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT104), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n346), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n341), .A2(new_n344), .A3(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n873), .A2(new_n278), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n345), .A2(new_n871), .A3(new_n346), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n357), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n876), .A2(new_n692), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n405), .A2(new_n877), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n388), .A2(KEYINPUT82), .A3(new_n378), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT82), .B1(new_n388), .B2(new_n378), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n876), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n400), .B1(new_n876), .B2(new_n692), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT37), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n692), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n359), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT37), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n390), .A2(new_n885), .A3(new_n886), .A4(new_n400), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT38), .B1(new_n878), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n878), .A2(KEYINPUT38), .A3(new_n888), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT40), .B1(new_n870), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n879), .A2(new_n880), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n403), .B1(new_n894), .B2(new_n359), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n895), .A2(KEYINPUT105), .A3(new_n886), .A4(new_n885), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT105), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n887), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n390), .A2(new_n400), .A3(new_n885), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT37), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n896), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n405), .A2(new_n359), .A3(new_n884), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT38), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT106), .ZN(new_n906));
  AND4_X1   g0706(.A1(new_n906), .A2(new_n878), .A3(KEYINPUT38), .A4(new_n888), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n405), .A2(new_n877), .B1(new_n883), .B2(new_n887), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n906), .B1(new_n908), .B2(KEYINPUT38), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n905), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(KEYINPUT40), .A3(new_n870), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT107), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n910), .A2(new_n870), .A3(KEYINPUT107), .A4(KEYINPUT40), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n893), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n915), .A2(new_n473), .A3(new_n864), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n915), .B1(new_n473), .B2(new_n864), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n916), .A2(new_n917), .A3(new_n737), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n470), .A2(new_n471), .A3(new_n695), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n890), .A2(KEYINPUT39), .A3(new_n891), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n891), .A2(KEYINPUT106), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n908), .A2(new_n906), .A3(KEYINPUT38), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n922), .A2(new_n923), .B1(new_n904), .B2(new_n903), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n920), .B(new_n921), .C1(new_n924), .C2(KEYINPUT39), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n679), .A2(new_n884), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n865), .B(new_n463), .C1(new_n470), .C2(new_n471), .ZN(new_n928));
  INV_X1    g0728(.A(new_n868), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n836), .B2(new_n826), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT103), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n892), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI211_X1 g0733(.A(KEYINPUT103), .B(new_n930), .C1(new_n836), .C2(new_n826), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n925), .B(new_n927), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  AND3_X1   g0735(.A1(new_n675), .A2(new_n723), .A3(new_n695), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n733), .A2(new_n663), .A3(new_n660), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n723), .B1(new_n937), .B2(new_n695), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n473), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n685), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n935), .B(new_n940), .Z(new_n941));
  OAI22_X1  g0741(.A1(new_n918), .A2(new_n941), .B1(new_n282), .B2(new_n687), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n941), .B2(new_n918), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n612), .A2(KEYINPUT35), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n612), .A2(KEYINPUT35), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n944), .A2(G116), .A3(new_n232), .A4(new_n945), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT36), .Z(new_n947));
  NAND3_X1  g0747(.A1(new_n229), .A2(G77), .A3(new_n342), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n207), .A2(G68), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n282), .B(G13), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  OR3_X1    g0750(.A1(new_n943), .A2(new_n947), .A3(new_n950), .ZN(G367));
  OAI211_X1 g0751(.A(new_n623), .B(new_n630), .C1(new_n695), .C2(new_n619), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n695), .A2(new_n630), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n712), .A2(new_n713), .A3(new_n954), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(KEYINPUT42), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n703), .A2(new_n623), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n694), .B1(new_n957), .B2(new_n630), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(new_n955), .B2(KEYINPUT42), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n695), .A2(new_n554), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n961), .A2(new_n725), .A3(new_n649), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(new_n725), .B2(new_n961), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT43), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n963), .A2(new_n964), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n960), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n956), .A2(new_n959), .A3(new_n964), .A4(new_n963), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n706), .A2(new_n954), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n969), .B(new_n970), .Z(new_n971));
  XOR2_X1   g0771(.A(new_n717), .B(KEYINPUT41), .Z(new_n972));
  AOI21_X1  g0772(.A(new_n954), .B1(new_n714), .B2(new_n704), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT44), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n714), .A2(new_n704), .A3(new_n954), .ZN(new_n976));
  XOR2_X1   g0776(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n976), .B(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n706), .B1(new_n975), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n712), .B(new_n713), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(new_n699), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n982), .A2(new_n754), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n973), .B(KEYINPUT44), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n976), .B(new_n977), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n984), .A2(new_n707), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n980), .A2(new_n983), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n972), .B1(new_n987), .B2(new_n755), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n971), .B1(new_n988), .B2(new_n804), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n810), .A2(new_n249), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n818), .B1(new_n238), .B2(new_n409), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n788), .A2(new_n764), .B1(new_n775), .B2(new_n215), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n295), .B(new_n992), .C1(G317), .C2(new_n779), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n782), .A2(G107), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n771), .A2(G116), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT46), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n855), .A2(new_n761), .B1(new_n772), .B2(new_n499), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G283), .B2(new_n786), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n993), .A2(new_n994), .A3(new_n996), .A4(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n782), .A2(G68), .ZN(new_n1000));
  INV_X1    g0800(.A(G150), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1000), .B1(new_n1001), .B2(new_n772), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1002), .A2(KEYINPUT109), .ZN(new_n1003));
  INV_X1    g0803(.A(G137), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n775), .A2(new_n411), .B1(new_n778), .B2(new_n1004), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n301), .B(new_n1005), .C1(G58), .C2(new_n771), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1002), .A2(KEYINPUT109), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n767), .A2(G143), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G159), .A2(new_n793), .B1(new_n786), .B2(G50), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n999), .B1(new_n1003), .B2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT47), .Z(new_n1012));
  INV_X1    g0812(.A(new_n757), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n805), .B1(new_n990), .B2(new_n991), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT110), .Z(new_n1015));
  NAND2_X1  g0815(.A1(new_n963), .A2(new_n817), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n989), .A2(new_n1017), .ZN(G387));
  OAI22_X1  g0818(.A1(new_n772), .A2(new_n207), .B1(new_n778), .B2(new_n1001), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n301), .B(new_n1019), .C1(G97), .C2(new_n776), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n791), .A2(new_n409), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n354), .A2(new_n793), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n763), .A2(new_n203), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n770), .A2(new_n411), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(G159), .C2(new_n767), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1020), .A2(new_n1022), .A3(new_n1023), .A4(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(G317), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n772), .A2(new_n1028), .B1(new_n763), .B2(new_n499), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1029), .A2(KEYINPUT111), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(KEYINPUT111), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G311), .A2(new_n793), .B1(new_n767), .B2(G322), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT48), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n791), .A2(new_n853), .B1(new_n770), .B2(new_n855), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(KEYINPUT49), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n295), .B1(new_n779), .B2(G326), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(new_n479), .C2(new_n775), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1038), .A2(KEYINPUT49), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1027), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT112), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1013), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n1044), .B2(new_n1043), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n808), .B1(G116), .B2(new_n546), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n246), .A2(new_n811), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n406), .A2(new_n207), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT50), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n719), .B(new_n310), .C1(new_n203), .C2(new_n411), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n810), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1047), .B1(G107), .B2(new_n238), .C1(new_n1048), .C2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n806), .B1(new_n1053), .B2(new_n818), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1046), .B(new_n1054), .C1(new_n713), .C2(new_n820), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n717), .B1(new_n754), .B2(new_n982), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n982), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1057), .A2(new_n755), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1055), .B1(new_n803), .B2(new_n982), .C1(new_n1056), .C2(new_n1058), .ZN(G393));
  NAND3_X1  g0859(.A1(new_n980), .A2(new_n986), .A3(new_n804), .ZN(new_n1060));
  NOR3_X1   g0860(.A1(new_n254), .A2(new_n716), .A3(new_n295), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n818), .B1(new_n215), .B2(new_n238), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n805), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n788), .A2(new_n1028), .B1(new_n772), .B2(new_n764), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT52), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G303), .A2(new_n793), .B1(new_n786), .B2(G294), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G283), .A2(new_n771), .B1(new_n779), .B2(G322), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n295), .B(new_n798), .C1(G116), .C2(new_n782), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G68), .A2(new_n771), .B1(new_n779), .B2(G143), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1070), .B(new_n295), .C1(new_n213), .C2(new_n775), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT114), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G50), .A2(new_n793), .B1(new_n786), .B2(new_n406), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1072), .B(new_n1073), .C1(new_n411), .C2(new_n791), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n773), .A2(G159), .B1(new_n767), .B2(G150), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT113), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT51), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1069), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1063), .B1(new_n1078), .B2(new_n757), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n954), .B2(new_n820), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n987), .A2(new_n717), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n983), .B1(new_n980), .B2(new_n986), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1060), .B(new_n1080), .C1(new_n1081), .C2(new_n1082), .ZN(G390));
  NAND2_X1  g0883(.A1(new_n829), .A2(new_n427), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n827), .B1(new_n734), .B2(new_n1084), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n928), .A2(KEYINPUT115), .A3(new_n929), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT115), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n867), .B2(new_n868), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n910), .B(new_n919), .C1(new_n1085), .C2(new_n1089), .ZN(new_n1090));
  AND3_X1   g0890(.A1(new_n878), .A2(KEYINPUT38), .A3(new_n888), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT39), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n1091), .A2(new_n889), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n910), .B2(new_n1092), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n931), .A2(new_n920), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1090), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n752), .A2(new_n830), .A3(new_n869), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1090), .B(new_n1097), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1099), .A2(new_n804), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n354), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n806), .B1(new_n1102), .B2(new_n859), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n799), .A2(new_n295), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1104), .B(new_n847), .C1(new_n215), .C2(new_n763), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n791), .A2(new_n411), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n788), .A2(new_n853), .B1(new_n772), .B2(new_n479), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n761), .A2(new_n421), .B1(new_n778), .B2(new_n855), .ZN(new_n1108));
  NOR4_X1   g0908(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n295), .B1(new_n775), .B2(new_n207), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT118), .Z(new_n1111));
  AOI22_X1  g0911(.A1(new_n773), .A2(G132), .B1(new_n767), .B2(G128), .ZN(new_n1112));
  INV_X1    g0912(.A(G125), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1112), .B1(new_n1113), .B2(new_n778), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n770), .A2(new_n1001), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  NOR3_X1   g0917(.A1(new_n1111), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT54), .B(G143), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n761), .A2(new_n1004), .B1(new_n763), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G159), .B2(new_n782), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT117), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1109), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1103), .B1(new_n1013), .B2(new_n1123), .C1(new_n1094), .C2(new_n816), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1101), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1089), .B1(new_n753), .B2(new_n831), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1127), .A2(new_n1097), .A3(new_n1085), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n836), .A2(new_n826), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n869), .B1(new_n752), .B2(new_n830), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1129), .B1(new_n1098), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(KEYINPUT116), .B1(new_n473), .B2(new_n752), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n473), .A2(new_n752), .A3(KEYINPUT116), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n939), .B(new_n685), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n718), .B1(new_n1126), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1135), .B1(new_n1131), .B2(new_n1128), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1139), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1125), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(G378));
  NAND2_X1  g0942(.A1(new_n915), .A2(G330), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n336), .A2(new_n433), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n884), .A2(new_n432), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1145), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1150), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1152), .A2(new_n1148), .A3(new_n1144), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n935), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n926), .B1(new_n1094), .B2(new_n920), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1129), .A2(new_n869), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(KEYINPUT103), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n931), .A2(new_n932), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(new_n1160), .A3(new_n892), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1154), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1143), .B1(new_n1156), .B2(new_n1162), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n737), .B(new_n893), .C1(new_n913), .C2(new_n914), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1157), .A2(new_n1161), .A3(new_n1154), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n935), .A2(new_n1155), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n803), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1155), .A2(new_n815), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n757), .A2(G50), .A3(new_n815), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n788), .A2(new_n1113), .B1(new_n761), .B2(new_n848), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1119), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n771), .A2(new_n1172), .B1(new_n786), .B2(G137), .ZN(new_n1173));
  INV_X1    g0973(.A(G128), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1173), .B1(new_n1174), .B2(new_n772), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1171), .B(new_n1175), .C1(G150), .C2(new_n782), .ZN(new_n1176));
  XOR2_X1   g0976(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  OR2_X1    g0978(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n776), .A2(G159), .ZN(new_n1181));
  AOI211_X1 g0981(.A(G33), .B(G41), .C1(new_n779), .C2(G124), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  NOR3_X1   g0983(.A1(new_n1025), .A2(G41), .A3(new_n295), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n776), .A2(G58), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n779), .A2(G283), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1184), .A2(new_n1000), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n788), .A2(new_n479), .B1(new_n763), .B2(new_n409), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n215), .A2(new_n761), .B1(new_n772), .B2(new_n421), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(KEYINPUT58), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1190), .A2(KEYINPUT58), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n207), .B1(new_n299), .B2(G41), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1183), .A2(new_n1191), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n806), .B(new_n1170), .C1(new_n1194), .C2(new_n757), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1169), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1168), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1140), .A2(new_n1136), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1166), .A2(new_n1165), .B1(new_n915), .B2(G330), .ZN(new_n1201));
  OAI211_X1 g1001(.A(KEYINPUT57), .B(new_n1199), .C1(new_n1200), .C2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n717), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1204));
  AOI21_X1  g1004(.A(KEYINPUT57), .B1(new_n1204), .B2(new_n1199), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1198), .B1(new_n1203), .B2(new_n1205), .ZN(G375));
  NAND2_X1  g1006(.A1(new_n1132), .A2(new_n804), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1089), .A2(new_n815), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n806), .B1(new_n203), .B2(new_n859), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n767), .A2(G294), .B1(new_n779), .B2(G303), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n215), .B2(new_n770), .C1(new_n853), .C2(new_n772), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n301), .B1(new_n775), .B2(new_n411), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n761), .A2(new_n479), .B1(new_n763), .B2(new_n421), .ZN(new_n1213));
  NOR4_X1   g1013(.A1(new_n1211), .A2(new_n1021), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G159), .A2(new_n771), .B1(new_n786), .B2(G150), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1174), .B2(new_n778), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1185), .B(new_n295), .C1(new_n207), .C2(new_n791), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT121), .Z(new_n1219));
  OAI22_X1  g1019(.A1(new_n788), .A2(new_n848), .B1(new_n772), .B2(new_n1004), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n793), .B2(new_n1172), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1214), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1208), .B(new_n1209), .C1(new_n1013), .C2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1207), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n972), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1135), .A2(new_n1128), .A3(new_n1131), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1137), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1225), .A2(new_n1228), .ZN(G381));
  NOR3_X1   g1029(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT122), .Z(new_n1231));
  NOR4_X1   g1031(.A1(new_n1231), .A2(G387), .A3(G390), .A4(G381), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n804), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n1196), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1202), .A2(new_n717), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT57), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1234), .B1(new_n1235), .B2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1232), .A2(new_n1141), .A3(new_n1239), .ZN(G407));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1141), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n693), .A2(G213), .ZN(new_n1242));
  OAI211_X1 g1042(.A(G407), .B(G213), .C1(new_n1241), .C2(new_n1242), .ZN(G409));
  NAND3_X1  g1043(.A1(new_n989), .A2(new_n1017), .A3(G390), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(KEYINPUT125), .ZN(new_n1245));
  XOR2_X1   g1045(.A(G393), .B(G396), .Z(new_n1246));
  INV_X1    g1046(.A(G390), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(G387), .A2(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1248), .A4(new_n1244), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1245), .A2(new_n1246), .B1(new_n1248), .B2(new_n1244), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1242), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1168), .A2(KEYINPUT123), .A3(new_n1197), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1226), .B(new_n1199), .C1(new_n1200), .C2(new_n1201), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1141), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(KEYINPUT123), .B1(new_n1168), .B2(new_n1197), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1254), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT62), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1227), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT60), .B1(new_n1227), .B2(KEYINPUT124), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1137), .A2(new_n717), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G384), .B(new_n1225), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1227), .A2(KEYINPUT124), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT60), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1266), .B1(new_n1270), .B2(new_n1262), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n862), .B1(new_n1271), .B2(new_n1224), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1267), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G375), .A2(G378), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1260), .A2(new_n1261), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1254), .A2(G2897), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1267), .A2(new_n1272), .A3(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1276), .B1(new_n1267), .B2(new_n1272), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT123), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1233), .A2(new_n1280), .A3(new_n1196), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1259), .A2(new_n1281), .A3(new_n1141), .A4(new_n1256), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1242), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1238), .A2(new_n717), .A3(new_n1202), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1141), .B1(new_n1284), .B2(new_n1198), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1279), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT61), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1275), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  XOR2_X1   g1088(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1289));
  NOR2_X1   g1089(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1289), .B1(new_n1290), .B2(new_n1273), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1253), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT63), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1274), .A2(new_n1242), .A3(new_n1282), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1273), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1293), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT61), .B1(new_n1294), .B2(new_n1279), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1290), .A2(KEYINPUT63), .A3(new_n1273), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1296), .A2(new_n1297), .A3(new_n1298), .A4(new_n1252), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1292), .A2(new_n1299), .ZN(G405));
  OAI211_X1 g1100(.A(KEYINPUT127), .B(new_n1273), .C1(new_n1250), .C2(new_n1251), .ZN(new_n1301));
  OR2_X1    g1101(.A1(new_n1273), .A2(KEYINPUT127), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1241), .A2(new_n1302), .A3(new_n1274), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1248), .A2(new_n1244), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1273), .A2(KEYINPUT127), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1306), .A2(new_n1249), .A3(new_n1307), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1301), .A2(new_n1303), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1303), .B1(new_n1301), .B2(new_n1308), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(G402));
endmodule


