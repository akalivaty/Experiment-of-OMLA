//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n555, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  XNOR2_X1  g029(.A(G325), .B(KEYINPUT64), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI21_X1  g032(.A(new_n456), .B1(new_n457), .B2(new_n452), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT65), .Z(G319));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n460), .A2(new_n461), .A3(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT66), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n461), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(new_n464), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n463), .A2(G2105), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n475), .A2(G2105), .B1(G101), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n470), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NAND4_X1  g054(.A1(new_n467), .A2(new_n462), .A3(G2105), .A4(new_n464), .ZN(new_n480));
  INV_X1    g055(.A(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n466), .A2(G112), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  OAI22_X1  g058(.A1(new_n480), .A2(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(new_n469), .B2(G136), .ZN(G162));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n467), .A2(new_n462), .A3(new_n464), .A4(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n473), .ZN(new_n489));
  NOR3_X1   g064(.A1(new_n486), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n488), .A2(KEYINPUT4), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G126), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT67), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G114), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n466), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  OAI22_X1  g073(.A1(new_n480), .A2(new_n492), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n491), .A2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G50), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G651), .ZN(new_n503));
  XNOR2_X1  g078(.A(new_n503), .B(KEYINPUT68), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT6), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n504), .A2(G543), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(KEYINPUT69), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n504), .A2(new_n513), .A3(new_n506), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n501), .A2(new_n507), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(new_n513), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G651), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n516), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  INV_X1    g099(.A(new_n507), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G51), .ZN(new_n526));
  INV_X1    g101(.A(new_n514), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G89), .ZN(new_n528));
  AND2_X1   g103(.A1(G63), .A2(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n513), .A2(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n526), .A2(new_n528), .A3(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n536), .A2(new_n507), .B1(new_n514), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n505), .ZN(new_n540));
  OR3_X1    g115(.A1(new_n538), .A2(KEYINPUT70), .A3(new_n540), .ZN(new_n541));
  OAI21_X1  g116(.A(KEYINPUT70), .B1(new_n538), .B2(new_n540), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(G171));
  AOI22_X1  g118(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n505), .ZN(new_n545));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n546), .A2(new_n507), .B1(new_n514), .B2(new_n547), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n548), .A2(KEYINPUT71), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(KEYINPUT71), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n545), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g129(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n555));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n507), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT73), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n513), .B(KEYINPUT74), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g141(.A1(G78), .A2(G543), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT75), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n569), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n570), .A2(new_n571), .B1(G91), .B2(new_n527), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n563), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  NAND4_X1  g149(.A1(new_n504), .A2(G49), .A3(G543), .A4(new_n506), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n504), .A2(G87), .A3(new_n513), .A4(new_n506), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT76), .ZN(G288));
  AOI22_X1  g154(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n505), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n504), .A2(G86), .A3(new_n513), .A4(new_n506), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n504), .A2(G48), .A3(G543), .A4(new_n506), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G305));
  AOI22_X1  g160(.A1(G47), .A2(new_n525), .B1(new_n527), .B2(G85), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n505), .B2(new_n587), .ZN(G290));
  INV_X1    g163(.A(G92), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n514), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT10), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n564), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g168(.A1(G79), .A2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n525), .A2(G54), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n591), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(G868), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g174(.A(new_n598), .B1(G868), .B2(G171), .ZN(G321));
  NAND2_X1  g175(.A1(G286), .A2(G868), .ZN(new_n601));
  INV_X1    g176(.A(G299), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G297));
  OAI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G280));
  INV_X1    g179(.A(G860), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n597), .B1(G559), .B2(new_n605), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT77), .Z(G148));
  NOR2_X1   g182(.A1(new_n597), .A2(G559), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n489), .A2(new_n476), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT12), .Z(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(G2100), .Z(new_n616));
  AND2_X1   g191(.A1(new_n469), .A2(G135), .ZN(new_n617));
  INV_X1    g192(.A(G123), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n466), .A2(G111), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  OAI22_X1  g195(.A1(new_n480), .A2(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G2096), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(G2096), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n616), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT78), .Z(G156));
  INV_X1    g202(.A(KEYINPUT14), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2427), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n631), .B2(new_n630), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n633), .B(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(G14), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n641), .B2(new_n639), .ZN(G401));
  XNOR2_X1  g218(.A(G2072), .B(G2078), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT17), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT79), .Z(new_n651));
  NAND3_X1  g226(.A1(new_n648), .A2(new_n644), .A3(new_n646), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT18), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n645), .A2(new_n646), .ZN(new_n654));
  INV_X1    g229(.A(new_n644), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n648), .B1(new_n655), .B2(new_n647), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n653), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2096), .B(G2100), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(G1971), .B(G1976), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  AND2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT20), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n663), .A2(new_n664), .ZN(new_n668));
  NOR3_X1   g243(.A1(new_n662), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n662), .B2(new_n668), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n671), .B(new_n672), .Z(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1981), .B(G1986), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G229));
  MUX2_X1   g253(.A(G6), .B(G305), .S(G16), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT32), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G1981), .ZN(new_n681));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G22), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT82), .Z(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(G166), .B2(new_n682), .ZN(new_n685));
  INV_X1    g260(.A(G1971), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n578), .A2(KEYINPUT81), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT81), .ZN(new_n689));
  NAND4_X1  g264(.A1(new_n575), .A2(new_n576), .A3(new_n689), .A4(new_n577), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G16), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G16), .B2(G23), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT33), .B(G1976), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n687), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(KEYINPUT34), .B1(new_n681), .B2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT83), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NOR3_X1   g275(.A1(new_n681), .A2(new_n697), .A3(KEYINPUT34), .ZN(new_n701));
  OR2_X1    g276(.A1(G25), .A2(G29), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n703));
  INV_X1    g278(.A(G107), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(G2105), .ZN(new_n705));
  INV_X1    g280(.A(new_n480), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(G119), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT80), .ZN(new_n708));
  AND3_X1   g283(.A1(new_n469), .A2(new_n708), .A3(G131), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n708), .B1(new_n469), .B2(G131), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n707), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n702), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT35), .B(G1991), .Z(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  MUX2_X1   g290(.A(G24), .B(G290), .S(G16), .Z(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(G1986), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n713), .A2(new_n714), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR3_X1   g294(.A1(new_n701), .A2(new_n715), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n700), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT84), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(KEYINPUT36), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n721), .A2(new_n722), .ZN(new_n725));
  OAI221_X1 g300(.A(KEYINPUT85), .B1(KEYINPUT36), .B2(new_n721), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  OR3_X1    g301(.A1(new_n724), .A2(KEYINPUT85), .A3(new_n725), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n469), .A2(G139), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT25), .ZN(new_n730));
  NAND2_X1  g305(.A1(G115), .A2(G2104), .ZN(new_n731));
  INV_X1    g306(.A(G127), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n473), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n730), .B1(G2105), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n728), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n735), .A2(new_n712), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n712), .B2(G33), .ZN(new_n737));
  INV_X1    g312(.A(G2072), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n623), .A2(new_n712), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT31), .B(G11), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT30), .B(G28), .Z(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(G29), .ZN(new_n744));
  OR4_X1    g319(.A1(new_n739), .A2(new_n740), .A3(new_n741), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT27), .B(G1996), .ZN(new_n746));
  OAI21_X1  g321(.A(KEYINPUT91), .B1(G29), .B2(G32), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT26), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n750), .A2(new_n751), .B1(G105), .B2(new_n476), .ZN(new_n752));
  INV_X1    g327(.A(G129), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n480), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n469), .B2(G141), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G29), .ZN(new_n756));
  MUX2_X1   g331(.A(KEYINPUT91), .B(new_n747), .S(new_n756), .Z(new_n757));
  AOI21_X1  g332(.A(new_n745), .B1(new_n746), .B2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G2084), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT89), .B(KEYINPUT24), .Z(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(G29), .B1(new_n761), .B2(G34), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G34), .B2(new_n761), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G160), .B2(new_n712), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT90), .ZN(new_n765));
  OAI221_X1 g340(.A(new_n758), .B1(new_n759), .B2(new_n765), .C1(new_n746), .C2(new_n757), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n759), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT92), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n682), .A2(G21), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G168), .B2(new_n682), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(G1966), .ZN(new_n772));
  NOR2_X1   g347(.A1(G164), .A2(new_n712), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G27), .B2(new_n712), .ZN(new_n774));
  INV_X1    g349(.A(G2078), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n771), .A2(G1966), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n774), .A2(new_n775), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n772), .A2(new_n776), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G29), .A2(G35), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G162), .B2(G29), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT29), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(G2090), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n782), .A2(G2090), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n779), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(G5), .A2(G16), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G171), .B2(G16), .ZN(new_n787));
  INV_X1    g362(.A(G1961), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n769), .A2(new_n785), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n682), .A2(G20), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT23), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n602), .B2(new_n682), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT93), .B(G1956), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G104), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n796), .A2(new_n466), .A3(KEYINPUT86), .ZN(new_n797));
  AOI21_X1  g372(.A(KEYINPUT86), .B1(new_n796), .B2(new_n466), .ZN(new_n798));
  OAI221_X1 g373(.A(G2104), .B1(G116), .B2(new_n466), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(G128), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n480), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G140), .B2(new_n469), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n802), .A2(new_n712), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT87), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n712), .A2(G26), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT28), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G2067), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n682), .A2(G19), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n552), .B2(new_n682), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G1341), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n682), .A2(G4), .ZN(new_n813));
  INV_X1    g388(.A(new_n597), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(new_n682), .ZN(new_n815));
  INV_X1    g390(.A(G1348), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n809), .A2(new_n812), .A3(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT88), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n790), .A2(new_n795), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n726), .A2(new_n727), .A3(new_n820), .ZN(G150));
  INV_X1    g396(.A(G150), .ZN(G311));
  NAND2_X1  g397(.A1(new_n814), .A2(G559), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT94), .B(KEYINPUT38), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(G55), .ZN(new_n826));
  INV_X1    g401(.A(G93), .ZN(new_n827));
  OAI22_X1  g402(.A1(new_n826), .A2(new_n507), .B1(new_n514), .B2(new_n827), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n829), .A2(new_n505), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n551), .B(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n825), .B(new_n832), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n833), .A2(KEYINPUT39), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(KEYINPUT39), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n834), .A2(new_n605), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n831), .A2(new_n605), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT37), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(G145));
  XNOR2_X1  g414(.A(new_n802), .B(G164), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n840), .A2(new_n755), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n755), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n841), .A2(new_n735), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n842), .ZN(new_n844));
  INV_X1    g419(.A(new_n735), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n711), .B(KEYINPUT95), .ZN(new_n847));
  INV_X1    g422(.A(new_n614), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n848), .ZN(new_n850));
  OR2_X1    g425(.A1(G106), .A2(G2105), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n851), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n852));
  INV_X1    g427(.A(G130), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n480), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(new_n469), .B2(G142), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n849), .A2(new_n850), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n855), .B1(new_n849), .B2(new_n850), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n843), .B(new_n846), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n846), .A2(new_n843), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n849), .A2(new_n850), .ZN(new_n860));
  INV_X1    g435(.A(new_n855), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n849), .A2(new_n850), .A3(new_n855), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n859), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n858), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n622), .B(new_n478), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G162), .ZN(new_n867));
  AOI21_X1  g442(.A(G37), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT96), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n858), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n856), .A2(new_n857), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n867), .B1(new_n871), .B2(new_n859), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n862), .A2(new_n863), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n873), .A2(KEYINPUT96), .A3(new_n843), .A4(new_n846), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n870), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n868), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT97), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n868), .A2(new_n875), .A3(KEYINPUT97), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(G395));
  XOR2_X1   g457(.A(new_n691), .B(G305), .Z(new_n883));
  XNOR2_X1  g458(.A(G166), .B(G290), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(KEYINPUT42), .Z(new_n886));
  XNOR2_X1  g461(.A(new_n568), .B(new_n569), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n527), .A2(G91), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n561), .B(KEYINPUT73), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n597), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n563), .A2(new_n572), .A3(new_n814), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(KEYINPUT41), .A3(new_n892), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n891), .A2(KEYINPUT99), .A3(new_n892), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT99), .B1(new_n891), .B2(new_n892), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n831), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n551), .B(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(new_n609), .ZN(new_n903));
  MUX2_X1   g478(.A(new_n897), .B(new_n900), .S(new_n903), .Z(new_n904));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n886), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n906), .B(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(G868), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(G868), .B2(new_n831), .ZN(G295));
  OAI21_X1  g485(.A(new_n909), .B1(G868), .B2(new_n831), .ZN(G331));
  INV_X1    g486(.A(KEYINPUT101), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n541), .A2(new_n912), .A3(new_n542), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(G286), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n912), .B1(new_n541), .B2(new_n542), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR3_X1   g491(.A1(G301), .A2(new_n912), .A3(G286), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n902), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n919));
  INV_X1    g494(.A(new_n915), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n920), .A2(G286), .A3(new_n913), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n914), .A2(new_n915), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n832), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n918), .A2(new_n919), .A3(new_n923), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n921), .A2(new_n832), .A3(KEYINPUT102), .A4(new_n922), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n918), .A2(new_n923), .ZN(new_n927));
  OAI22_X1  g502(.A1(new_n926), .A2(new_n897), .B1(new_n900), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n885), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT103), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n931));
  INV_X1    g506(.A(new_n893), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n891), .A2(KEYINPUT41), .A3(new_n892), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT41), .B1(new_n891), .B2(new_n892), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI22_X1  g510(.A1(new_n926), .A2(new_n932), .B1(new_n935), .B2(new_n927), .ZN(new_n936));
  INV_X1    g511(.A(new_n885), .ZN(new_n937));
  AOI21_X1  g512(.A(G37), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT103), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n928), .A2(new_n939), .A3(new_n885), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n930), .A2(new_n931), .A3(new_n938), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n936), .A2(new_n937), .ZN(new_n942));
  INV_X1    g517(.A(G37), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n927), .A2(new_n895), .A3(new_n896), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n893), .B1(new_n924), .B2(new_n925), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n885), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n942), .A2(new_n943), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n941), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n931), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n930), .A2(new_n938), .A3(new_n940), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n951), .B1(new_n952), .B2(new_n931), .ZN(new_n953));
  MUX2_X1   g528(.A(new_n950), .B(new_n953), .S(KEYINPUT44), .Z(G397));
  NAND2_X1  g529(.A1(G303), .A2(G8), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT55), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n955), .B(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G1384), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(new_n491), .B2(new_n499), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT45), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n470), .A2(G40), .A3(new_n477), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT45), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n959), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n961), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n686), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n962), .B1(KEYINPUT50), .B2(new_n959), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n959), .A2(KEYINPUT106), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n971), .B(new_n958), .C1(new_n491), .C2(new_n499), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n968), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n967), .B1(G2090), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n957), .A2(new_n975), .A3(G8), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT107), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n977), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n583), .A2(new_n584), .ZN(new_n982));
  OAI21_X1  g557(.A(G1981), .B1(new_n982), .B2(new_n581), .ZN(new_n983));
  INV_X1    g558(.A(G1981), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n582), .A2(new_n984), .A3(new_n583), .A4(new_n584), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT49), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n987), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT109), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n986), .A2(new_n991), .A3(new_n987), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n988), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n489), .A2(new_n490), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n706), .A2(G126), .ZN(new_n997));
  OR2_X1    g572(.A1(new_n497), .A2(new_n498), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n971), .B1(new_n999), .B2(new_n958), .ZN(new_n1000));
  INV_X1    g575(.A(new_n972), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n1000), .A2(new_n1001), .A3(new_n962), .ZN(new_n1002));
  INV_X1    g577(.A(G8), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n993), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n688), .A2(G1976), .A3(new_n690), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n1006), .A2(KEYINPUT108), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(KEYINPUT108), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1004), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT52), .ZN(new_n1010));
  INV_X1    g585(.A(G1976), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT52), .B1(G288), .B2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1004), .A2(new_n1012), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1005), .A2(new_n1010), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G288), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1005), .A2(new_n1011), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n985), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n981), .A2(new_n1015), .B1(new_n1004), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n957), .B1(new_n975), .B2(G8), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1020), .B1(new_n1014), .B2(new_n1021), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1004), .A2(new_n993), .B1(new_n1009), .B2(KEYINPUT52), .ZN(new_n1023));
  INV_X1    g598(.A(new_n957), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n975), .A2(G8), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1023), .A2(new_n1026), .A3(KEYINPUT114), .A4(new_n1013), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n974), .ZN(new_n1029));
  XNOR2_X1  g604(.A(KEYINPUT113), .B(G2084), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n964), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT111), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(new_n963), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT45), .B1(new_n969), .B2(new_n972), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT111), .B1(new_n1036), .B2(new_n962), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n1037), .A3(new_n961), .ZN(new_n1038));
  INV_X1    g613(.A(G1966), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1032), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1038), .A2(KEYINPUT112), .A3(new_n1039), .ZN(new_n1043));
  AOI211_X1 g618(.A(new_n1003), .B(G286), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT63), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(new_n978), .B2(new_n979), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1028), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT115), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT110), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n962), .B1(new_n960), .B2(new_n970), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1050), .B1(new_n1051), .B2(new_n970), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(G2090), .ZN(new_n1053));
  INV_X1    g628(.A(new_n967), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1049), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G8), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1053), .A2(new_n1049), .A3(new_n1054), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1024), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n980), .A2(new_n1058), .A3(new_n1015), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1060), .A2(new_n1043), .A3(new_n1031), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(G8), .A3(G168), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1045), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1048), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1047), .A2(KEYINPUT115), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1019), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n561), .A2(KEYINPUT57), .ZN(new_n1067));
  AOI22_X1  g642(.A1(G299), .A2(KEYINPUT57), .B1(new_n572), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1956), .ZN(new_n1069));
  INV_X1    g644(.A(new_n966), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT56), .B(G2072), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1052), .A2(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1068), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1068), .A2(new_n1072), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n974), .A2(new_n816), .B1(new_n1002), .B2(new_n808), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(new_n597), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1073), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT116), .B(KEYINPUT58), .ZN(new_n1078));
  XOR2_X1   g653(.A(new_n1078), .B(G1341), .Z(new_n1079));
  OR2_X1    g654(.A1(new_n1002), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1996), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1070), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n551), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  XOR2_X1   g658(.A(new_n1083), .B(KEYINPUT59), .Z(new_n1084));
  NAND2_X1  g659(.A1(new_n1073), .A2(KEYINPUT61), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1075), .A2(KEYINPUT60), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n597), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT61), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1068), .A2(new_n1088), .A3(new_n1072), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .A4(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1075), .A2(KEYINPUT60), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1086), .A2(new_n1091), .A3(new_n597), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1077), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT54), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1070), .A2(new_n775), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1095), .A2(new_n1096), .B1(new_n788), .B2(new_n974), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n775), .A2(KEYINPUT53), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(new_n1098), .B2(new_n966), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(G171), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1038), .A2(new_n1098), .ZN(new_n1101));
  AOI21_X1  g676(.A(G301), .B1(new_n1101), .B2(new_n1097), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1094), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  OR2_X1    g678(.A1(new_n1103), .A2(KEYINPUT120), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(KEYINPUT120), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1099), .A2(G171), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1101), .A2(G301), .A3(new_n1097), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(KEYINPUT54), .A3(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1093), .A2(new_n1104), .A3(new_n1105), .A4(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1059), .B(KEYINPUT121), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n1112));
  XOR2_X1   g687(.A(KEYINPUT117), .B(KEYINPUT51), .Z(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(G286), .A2(G8), .ZN(new_n1115));
  XOR2_X1   g690(.A(new_n1115), .B(KEYINPUT118), .Z(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1038), .A2(KEYINPUT112), .A3(new_n1039), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT112), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1118), .A2(new_n1119), .A3(new_n1032), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1117), .B1(new_n1120), .B2(new_n1003), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1114), .B1(new_n1121), .B2(new_n1062), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1061), .A2(G8), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1112), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1116), .B1(new_n1061), .B2(G8), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1113), .B1(new_n1044), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1129), .A2(KEYINPUT119), .A3(new_n1125), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1066), .B1(new_n1111), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1127), .A2(new_n1133), .A3(new_n1130), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1059), .A2(KEYINPUT121), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1059), .A2(KEYINPUT121), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1135), .A2(new_n1102), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1134), .A2(KEYINPUT122), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1131), .A2(KEYINPUT62), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT122), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1132), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n802), .B(new_n808), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1143), .B(KEYINPUT105), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n755), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1145), .B1(G1996), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n965), .A2(new_n962), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n1148), .B(KEYINPUT104), .Z(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1081), .ZN(new_n1151));
  OAI22_X1  g726(.A1(new_n1147), .A2(new_n1150), .B1(new_n1146), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n711), .B(new_n714), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1153), .B1(new_n1154), .B2(new_n1150), .ZN(new_n1155));
  XNOR2_X1  g730(.A(G290), .B(G1986), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1155), .B1(new_n1148), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1142), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n714), .ZN(new_n1159));
  OR3_X1    g734(.A1(new_n1152), .A2(new_n711), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n802), .A2(new_n808), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1150), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1149), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1151), .B(KEYINPUT46), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT47), .ZN(new_n1169));
  NOR2_X1   g744(.A1(G290), .A2(G1986), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n1148), .ZN(new_n1171));
  XOR2_X1   g746(.A(new_n1171), .B(KEYINPUT124), .Z(new_n1172));
  XNOR2_X1  g747(.A(new_n1172), .B(KEYINPUT48), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1169), .B1(new_n1155), .B2(new_n1173), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1164), .A2(new_n1165), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1158), .A2(new_n1175), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n1178));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n1179));
  NOR3_X1   g753(.A1(G401), .A2(new_n458), .A3(G227), .ZN(new_n1180));
  INV_X1    g754(.A(KEYINPUT125), .ZN(new_n1181));
  OR2_X1    g755(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1183));
  NAND3_X1  g757(.A1(new_n677), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  AOI21_X1  g758(.A(new_n1184), .B1(new_n878), .B2(new_n879), .ZN(new_n1185));
  AND3_X1   g759(.A1(new_n950), .A2(new_n1179), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g760(.A(new_n1179), .B1(new_n950), .B2(new_n1185), .ZN(new_n1187));
  OAI21_X1  g761(.A(new_n1178), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g762(.A1(new_n950), .A2(new_n1185), .ZN(new_n1189));
  NAND2_X1  g763(.A1(new_n1189), .A2(KEYINPUT126), .ZN(new_n1190));
  NAND3_X1  g764(.A1(new_n950), .A2(new_n1179), .A3(new_n1185), .ZN(new_n1191));
  NAND3_X1  g765(.A1(new_n1190), .A2(KEYINPUT127), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n1188), .A2(new_n1192), .ZN(G308));
  NAND2_X1  g767(.A1(new_n1190), .A2(new_n1191), .ZN(G225));
endmodule


