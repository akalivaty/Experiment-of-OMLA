//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1250, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n202), .B(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G97), .A2(G257), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G87), .A2(G250), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT66), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AND2_X1   g0014(.A1(new_n212), .A2(new_n213), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n214), .B(new_n215), .C1(G77), .C2(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G116), .ZN(new_n219));
  INV_X1    g0019(.A(G270), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AND2_X1   g0021(.A1(KEYINPUT65), .A2(G68), .ZN(new_n222));
  NOR2_X1   g0022(.A1(KEYINPUT65), .A2(G68), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AND2_X1   g0024(.A1(new_n224), .A2(G238), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n208), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT1), .Z(new_n227));
  NOR2_X1   g0027(.A1(new_n208), .A2(G13), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT0), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G20), .ZN(new_n233));
  NOR2_X1   g0033(.A1(G58), .A2(G68), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n235), .A2(G50), .ZN(new_n236));
  OAI211_X1 g0036(.A(new_n227), .B(new_n230), .C1(new_n233), .C2(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(KEYINPUT67), .Z(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G226), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G264), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n220), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT69), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G68), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G107), .B(G116), .Z(new_n252));
  XNOR2_X1  g0052(.A(G87), .B(G97), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n251), .B(new_n254), .Z(G351));
  NAND2_X1  g0055(.A1(G33), .A2(G97), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n257), .B1(G232), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G226), .A2(G1698), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n232), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n261), .A2(new_n262), .B1(G238), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT13), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g0072(.A(new_n272), .B(KEYINPUT75), .Z(new_n273));
  AND3_X1   g0073(.A1(new_n269), .A2(new_n270), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n270), .B1(new_n269), .B2(new_n273), .ZN(new_n275));
  OAI211_X1 g0075(.A(KEYINPUT77), .B(G169), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT14), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n269), .A2(new_n273), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT13), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n269), .A2(new_n270), .A3(new_n273), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT14), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n281), .A2(KEYINPUT77), .A3(new_n282), .A4(G169), .ZN(new_n283));
  INV_X1    g0083(.A(G179), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n277), .B(new_n283), .C1(new_n284), .C2(new_n281), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT72), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n287), .A2(new_n231), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n286), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AND4_X1   g0090(.A1(new_n286), .A2(new_n289), .A3(new_n231), .A4(new_n287), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n292), .B1(new_n205), .B2(G20), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT12), .ZN(new_n294));
  OAI21_X1  g0094(.A(G68), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n289), .A2(new_n294), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n205), .A2(G13), .ZN(new_n298));
  OR4_X1    g0098(.A1(new_n294), .A2(new_n224), .A3(new_n206), .A4(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT70), .B1(new_n263), .B2(G20), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT70), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(new_n206), .A3(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(G20), .A2(G33), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n303), .A2(G77), .B1(G50), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(new_n206), .B2(new_n224), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n287), .A2(new_n231), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT76), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT76), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n306), .A2(new_n310), .A3(new_n307), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n309), .A2(KEYINPUT11), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT11), .B1(new_n309), .B2(new_n311), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n297), .B(new_n299), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n285), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G200), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n279), .B2(new_n280), .ZN(new_n317));
  INV_X1    g0117(.A(G190), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n281), .A2(new_n318), .ZN(new_n319));
  OR3_X1    g0119(.A1(new_n314), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT78), .ZN(new_n322));
  OR2_X1    g0122(.A1(KEYINPUT65), .A2(G68), .ZN(new_n323));
  NAND2_X1  g0123(.A1(KEYINPUT65), .A2(G68), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n323), .A2(G58), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n206), .B1(new_n325), .B2(new_n235), .ZN(new_n326));
  INV_X1    g0126(.A(new_n304), .ZN(new_n327));
  INV_X1    g0127(.A(G159), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n322), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n329), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n234), .B1(new_n224), .B2(G58), .ZN(new_n332));
  OAI211_X1 g0132(.A(KEYINPUT78), .B(new_n331), .C1(new_n332), .C2(new_n206), .ZN(new_n333));
  AND2_X1   g0133(.A1(KEYINPUT3), .A2(G33), .ZN(new_n334));
  NOR2_X1   g0134(.A1(KEYINPUT3), .A2(G33), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT7), .B1(new_n336), .B2(new_n206), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT7), .ZN(new_n338));
  NOR4_X1   g0138(.A1(new_n334), .A2(new_n335), .A3(new_n338), .A4(G20), .ZN(new_n339));
  OAI21_X1  g0139(.A(G68), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n330), .A2(new_n333), .A3(KEYINPUT16), .A4(new_n340), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n341), .A2(new_n307), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n224), .B1(new_n337), .B2(new_n339), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n330), .A2(new_n333), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT16), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  XOR2_X1   g0147(.A(KEYINPUT8), .B(G58), .Z(new_n348));
  NAND2_X1  g0148(.A1(new_n205), .A2(G20), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n289), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(new_n307), .ZN(new_n353));
  INV_X1    g0153(.A(new_n348), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n351), .A2(new_n353), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n218), .A2(G1698), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n257), .B(new_n356), .C1(G223), .C2(G1698), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G87), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n265), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G232), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n267), .A2(new_n360), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n359), .A2(new_n361), .A3(new_n272), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n318), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n362), .B2(G200), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n347), .A2(new_n355), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT17), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n355), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n342), .B2(new_n346), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(KEYINPUT17), .A3(new_n364), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT18), .ZN(new_n371));
  NOR4_X1   g0171(.A1(new_n359), .A2(new_n361), .A3(new_n284), .A4(new_n272), .ZN(new_n372));
  OR3_X1    g0172(.A1(new_n359), .A2(new_n361), .A3(new_n272), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n372), .B1(G169), .B2(new_n373), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n369), .A2(new_n371), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n346), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n341), .A2(new_n307), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n355), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n372), .ZN(new_n379));
  INV_X1    g0179(.A(G169), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n379), .B1(new_n380), .B2(new_n362), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT18), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n367), .B(new_n370), .C1(new_n375), .C2(new_n382), .ZN(new_n383));
  OR2_X1    g0183(.A1(KEYINPUT15), .A2(G87), .ZN(new_n384));
  NAND2_X1  g0184(.A1(KEYINPUT15), .A2(G87), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n303), .ZN(new_n388));
  INV_X1    g0188(.A(G77), .ZN(new_n389));
  XOR2_X1   g0189(.A(new_n348), .B(KEYINPUT71), .Z(new_n390));
  OAI221_X1 g0190(.A(new_n388), .B1(new_n206), .B2(new_n389), .C1(new_n390), .C2(new_n327), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n391), .A2(new_n307), .B1(G77), .B2(new_n293), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n352), .A2(new_n389), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(G238), .A2(G1698), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n257), .B(new_n395), .C1(new_n360), .C2(G1698), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n396), .B(new_n262), .C1(G107), .C2(new_n257), .ZN(new_n397));
  INV_X1    g0197(.A(new_n272), .ZN(new_n398));
  INV_X1    g0198(.A(G244), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n397), .B(new_n398), .C1(new_n399), .C2(new_n267), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G200), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n400), .A2(new_n318), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n394), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  OR3_X1    g0204(.A1(new_n321), .A2(new_n383), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n353), .A2(G50), .A3(new_n349), .ZN(new_n406));
  INV_X1    g0206(.A(G150), .ZN(new_n407));
  NOR3_X1   g0207(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n407), .A2(new_n327), .B1(new_n408), .B2(new_n206), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(new_n348), .B2(new_n303), .ZN(new_n410));
  OAI221_X1 g0210(.A(new_n406), .B1(G50), .B2(new_n289), .C1(new_n410), .C2(new_n288), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT73), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n411), .B(new_n412), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n413), .B(KEYINPUT9), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n258), .A2(G222), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G223), .A2(G1698), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n257), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n417), .B(new_n262), .C1(G77), .C2(new_n257), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n418), .B(new_n398), .C1(new_n218), .C2(new_n267), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n419), .A2(new_n318), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(G200), .B2(new_n419), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n414), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT74), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT10), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n424), .ZN(new_n426));
  NAND2_X1  g0226(.A1(KEYINPUT74), .A2(KEYINPUT10), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n414), .A2(new_n426), .A3(new_n427), .A4(new_n421), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n419), .A2(new_n380), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(new_n411), .C1(G179), .C2(new_n419), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n400), .A2(new_n380), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n394), .B(new_n431), .C1(G179), .C2(new_n400), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n425), .A2(new_n428), .A3(new_n430), .A4(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n405), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT82), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n386), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n384), .A2(KEYINPUT82), .A3(new_n385), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n205), .A2(G33), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n288), .A2(new_n289), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT83), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n439), .A2(new_n441), .A3(KEYINPUT83), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT81), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT19), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n206), .B1(new_n256), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G87), .ZN(new_n449));
  INV_X1    g0249(.A(G97), .ZN(new_n450));
  INV_X1    g0250(.A(G107), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n206), .B(G68), .C1(new_n334), .C2(new_n335), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n450), .B1(new_n300), .B2(new_n302), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n453), .B(new_n454), .C1(new_n455), .C2(KEYINPUT19), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n307), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n387), .A2(new_n289), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n446), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  AOI211_X1 g0260(.A(KEYINPUT81), .B(new_n458), .C1(new_n456), .C2(new_n307), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n445), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n399), .A2(G1698), .ZN(new_n463));
  OAI221_X1 g0263(.A(new_n463), .B1(G238), .B2(G1698), .C1(new_n334), .C2(new_n335), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G116), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n265), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n205), .A2(G45), .A3(G274), .ZN(new_n467));
  INV_X1    g0267(.A(G45), .ZN(new_n468));
  OAI21_X1  g0268(.A(G250), .B1(new_n468), .B2(G1), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n262), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NOR3_X1   g0270(.A1(new_n466), .A2(G179), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n470), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n464), .A2(new_n465), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(new_n265), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n471), .B1(new_n380), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n462), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n316), .B1(new_n466), .B2(new_n470), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n474), .B2(G190), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n441), .A2(G87), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n478), .B(new_n479), .C1(new_n461), .C2(new_n460), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n206), .B(G87), .C1(new_n334), .C2(new_n335), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT22), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT22), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n257), .A2(new_n483), .A3(new_n206), .A4(G87), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n206), .A2(G107), .ZN(new_n486));
  XNOR2_X1  g0286(.A(new_n486), .B(KEYINPUT23), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n465), .A2(G20), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT24), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n488), .B1(new_n482), .B2(new_n484), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(KEYINPUT24), .A3(new_n487), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n307), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n441), .A2(G107), .ZN(new_n496));
  INV_X1    g0296(.A(G13), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(G1), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n486), .ZN(new_n499));
  XNOR2_X1  g0299(.A(new_n499), .B(KEYINPUT25), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  XNOR2_X1  g0301(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT80), .B1(new_n502), .B2(G41), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT80), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT5), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n505), .A2(KEYINPUT79), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n505), .A2(KEYINPUT79), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n504), .B(new_n264), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  AOI211_X1 g0308(.A(G1), .B(new_n468), .C1(new_n505), .C2(G41), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n503), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(G264), .A3(new_n265), .ZN(new_n511));
  XOR2_X1   g0311(.A(KEYINPUT87), .B(G294), .Z(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G33), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n257), .B1(G257), .B2(new_n258), .ZN(new_n514));
  NOR2_X1   g0314(.A1(G250), .A2(G1698), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n262), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n467), .B1(new_n505), .B2(G41), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n503), .A2(new_n508), .A3(new_n265), .A4(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n511), .A2(new_n517), .A3(G190), .A4(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n495), .A2(new_n496), .A3(new_n501), .A4(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n511), .A2(new_n517), .A3(new_n519), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G200), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n476), .B(new_n480), .C1(new_n521), .C2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT6), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n526), .A2(new_n450), .A3(G107), .ZN(new_n527));
  XNOR2_X1  g0327(.A(G97), .B(G107), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n527), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  OAI22_X1  g0329(.A1(new_n529), .A2(new_n206), .B1(new_n389), .B2(new_n327), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n338), .B1(new_n257), .B2(G20), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n336), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n451), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n307), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n441), .A2(G97), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n289), .A2(G97), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G33), .A2(G283), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n258), .A2(KEYINPUT4), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n257), .A2(G244), .A3(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n336), .A2(new_n399), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n540), .B(new_n542), .C1(new_n543), .C2(KEYINPUT4), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n257), .A2(G250), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n258), .B1(new_n545), .B2(KEYINPUT4), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n262), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n510), .A2(G257), .A3(new_n265), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(new_n519), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G200), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n547), .A2(G190), .A3(new_n519), .A4(new_n548), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n539), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(new_n380), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n547), .A2(new_n284), .A3(new_n519), .A4(new_n548), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n538), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n525), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n510), .A2(G270), .A3(new_n265), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n258), .A2(G257), .ZN(new_n559));
  NAND2_X1  g0359(.A1(G264), .A2(G1698), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n257), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n561), .B(new_n262), .C1(G303), .C2(new_n257), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n558), .A2(new_n562), .A3(new_n519), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n563), .A2(KEYINPUT21), .A3(G169), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n558), .A2(G179), .A3(new_n562), .A4(new_n519), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(G116), .B(new_n440), .C1(new_n290), .C2(new_n291), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n498), .A2(G20), .A3(new_n219), .ZN(new_n568));
  XNOR2_X1  g0368(.A(new_n568), .B(KEYINPUT84), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n540), .B(new_n206), .C1(G33), .C2(new_n450), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n219), .A2(G20), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n570), .A2(new_n307), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT20), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n570), .A2(KEYINPUT20), .A3(new_n307), .A4(new_n571), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n567), .A2(new_n569), .A3(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT85), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n567), .A2(new_n576), .A3(KEYINPUT85), .A4(new_n569), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n566), .A2(KEYINPUT86), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT86), .B1(new_n566), .B2(new_n581), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n522), .A2(G169), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n511), .A2(new_n517), .A3(G179), .A4(new_n519), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(KEYINPUT88), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n495), .A2(new_n496), .A3(new_n501), .ZN(new_n588));
  OR2_X1    g0388(.A1(new_n586), .A2(KEYINPUT88), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT21), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n579), .A2(new_n580), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n563), .A2(G169), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n563), .A2(G200), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n318), .B2(new_n563), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n597), .A2(new_n581), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n557), .A2(new_n584), .A3(new_n595), .A4(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n435), .A2(new_n600), .ZN(G372));
  NOR3_X1   g0401(.A1(new_n314), .A2(new_n317), .A3(new_n319), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n315), .B1(new_n602), .B2(new_n432), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n603), .A2(new_n367), .A3(new_n370), .ZN(new_n604));
  OR2_X1    g0404(.A1(new_n375), .A2(new_n382), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n425), .A2(new_n428), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n608), .A2(new_n430), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n566), .A2(new_n581), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n595), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n557), .ZN(new_n612));
  INV_X1    g0412(.A(new_n476), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT26), .ZN(new_n614));
  INV_X1    g0414(.A(new_n444), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n615), .A2(new_n442), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n457), .A2(new_n459), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT81), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n457), .A2(new_n446), .A3(new_n459), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n475), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n480), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n614), .B1(new_n622), .B2(new_n555), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n553), .A2(new_n538), .A3(new_n554), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n624), .A2(KEYINPUT26), .A3(new_n476), .A4(new_n480), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n613), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n612), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n609), .B1(new_n435), .B2(new_n628), .ZN(G369));
  INV_X1    g0429(.A(new_n593), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT21), .B1(new_n630), .B2(new_n581), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n564), .A2(new_n565), .B1(new_n579), .B2(new_n580), .ZN(new_n632));
  OR3_X1    g0432(.A1(new_n298), .A2(KEYINPUT27), .A3(G20), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT27), .B1(new_n298), .B2(G20), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(G213), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(G343), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n581), .A2(new_n637), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n631), .A2(new_n632), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT86), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n610), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n632), .A2(KEYINPUT86), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(new_n642), .A3(new_n594), .ZN(new_n643));
  AOI211_X1 g0443(.A(new_n598), .B(new_n639), .C1(new_n643), .C2(new_n638), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n590), .A2(new_n637), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n493), .A2(KEYINPUT24), .A3(new_n487), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT24), .B1(new_n493), .B2(new_n487), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n500), .B1(new_n648), .B2(new_n307), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n649), .A2(new_n496), .A3(new_n523), .A4(new_n520), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n588), .A2(new_n637), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n645), .B1(new_n590), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n644), .A2(G330), .A3(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n645), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n521), .A2(new_n524), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n588), .A2(new_n589), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n656), .B1(new_n657), .B2(new_n587), .ZN(new_n658));
  INV_X1    g0458(.A(new_n637), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n643), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n654), .A2(new_n655), .A3(new_n660), .ZN(G399));
  INV_X1    g0461(.A(new_n228), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(G41), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n452), .A2(G116), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G1), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n236), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT28), .ZN(new_n668));
  INV_X1    g0468(.A(new_n479), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n618), .B2(new_n619), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n670), .A2(new_n478), .B1(new_n462), .B2(new_n475), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n650), .A2(new_n671), .A3(new_n555), .A4(new_n552), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n672), .B1(new_n584), .B2(new_n595), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n622), .A2(new_n614), .A3(new_n555), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT26), .B1(new_n671), .B2(new_n624), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n476), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n659), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT91), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n641), .A2(new_n642), .A3(new_n594), .A4(new_n590), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n557), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n626), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT91), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(new_n682), .A3(new_n659), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n678), .A2(KEYINPUT29), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n637), .B1(new_n612), .B2(new_n626), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT29), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT30), .ZN(new_n688));
  INV_X1    g0488(.A(new_n549), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT90), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n466), .A2(new_n470), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n511), .A2(new_n691), .A3(new_n517), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n689), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n690), .ZN(new_n694));
  INV_X1    g0494(.A(new_n565), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n688), .B1(new_n693), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n689), .A2(G179), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n698), .A2(new_n563), .A3(new_n522), .A4(new_n474), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n565), .B1(new_n690), .B2(new_n692), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n692), .A2(new_n690), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n700), .A2(new_n701), .A3(KEYINPUT30), .A4(new_n689), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n697), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n637), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT31), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g0506(.A(KEYINPUT89), .B(KEYINPUT31), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n703), .A2(new_n637), .A3(new_n707), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n706), .B(new_n708), .C1(new_n600), .C2(new_n637), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(G330), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n684), .A2(new_n687), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n668), .B1(new_n712), .B2(G1), .ZN(G364));
  INV_X1    g0513(.A(new_n644), .ZN(new_n714));
  NOR2_X1   g0514(.A1(G13), .A2(G33), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G20), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n231), .B1(G20), .B2(new_n380), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g0520(.A(new_n720), .B(KEYINPUT94), .Z(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n228), .A2(new_n257), .ZN(new_n723));
  OAI22_X1  g0523(.A1(new_n723), .A2(new_n203), .B1(G116), .B2(new_n228), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n724), .B(KEYINPUT93), .Z(new_n725));
  NOR2_X1   g0525(.A1(new_n662), .A2(new_n257), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(G45), .B2(new_n236), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n727), .B1(new_n251), .B2(G45), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n722), .B1(new_n725), .B2(new_n728), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n497), .A2(new_n468), .A3(G20), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n730), .A2(KEYINPUT92), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(KEYINPUT92), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n731), .A2(G1), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n663), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n735), .A2(KEYINPUT96), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(KEYINPUT96), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n736), .A2(new_n318), .A3(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  XOR2_X1   g0539(.A(KEYINPUT33), .B(G317), .Z(new_n740));
  INV_X1    g0540(.A(G322), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n206), .A2(new_n318), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n284), .A2(G200), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n739), .A2(new_n740), .B1(new_n741), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g0546(.A(new_n746), .B(KEYINPUT101), .Z(new_n747));
  NOR2_X1   g0547(.A1(new_n316), .A2(G179), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n742), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n747), .B1(G303), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G179), .A2(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G190), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n512), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n736), .A2(G190), .A3(new_n737), .ZN(new_n756));
  INV_X1    g0556(.A(G326), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT99), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G283), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n206), .A2(G190), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n762), .A2(KEYINPUT97), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(KEYINPUT97), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n763), .A2(new_n764), .A3(new_n748), .ZN(new_n765));
  OAI221_X1 g0565(.A(new_n336), .B1(new_n761), .B2(new_n765), .C1(new_n758), .C2(new_n759), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n763), .A2(new_n752), .A3(new_n764), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT100), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n766), .B1(G329), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n751), .A2(new_n760), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n743), .A2(new_n762), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n771), .B1(G311), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n767), .A2(new_n328), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT32), .ZN(new_n776));
  INV_X1    g0576(.A(G58), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n745), .A2(new_n777), .B1(new_n389), .B2(new_n772), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT95), .ZN(new_n779));
  INV_X1    g0579(.A(new_n765), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n778), .A2(new_n779), .B1(new_n780), .B2(G107), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n776), .B(new_n781), .C1(new_n217), .C2(new_n756), .ZN(new_n782));
  INV_X1    g0582(.A(new_n754), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n450), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n778), .A2(new_n779), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT98), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n749), .A2(new_n449), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(new_n787), .B2(new_n336), .ZN(new_n788));
  OAI211_X1 g0588(.A(KEYINPUT98), .B(new_n257), .C1(new_n749), .C2(new_n449), .ZN(new_n789));
  INV_X1    g0589(.A(G68), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n788), .B(new_n789), .C1(new_n739), .C2(new_n790), .ZN(new_n791));
  NOR4_X1   g0591(.A1(new_n782), .A2(new_n784), .A3(new_n785), .A4(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n719), .B1(new_n774), .B2(new_n792), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n718), .A2(new_n729), .A3(new_n734), .A4(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G330), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n714), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n598), .B1(new_n643), .B2(new_n638), .ZN(new_n797));
  INV_X1    g0597(.A(new_n639), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n797), .A2(G330), .A3(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n734), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n796), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n794), .A2(new_n801), .ZN(G396));
  OR2_X1    g0602(.A1(new_n432), .A2(new_n637), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n659), .B1(new_n392), .B2(new_n393), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n432), .B1(new_n404), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n716), .ZN(new_n808));
  INV_X1    g0608(.A(new_n719), .ZN(new_n809));
  INV_X1    g0609(.A(G311), .ZN(new_n810));
  XNOR2_X1  g0610(.A(KEYINPUT102), .B(G283), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n768), .A2(new_n810), .B1(new_n739), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n765), .A2(new_n449), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n772), .A2(new_n219), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n336), .B1(new_n749), .B2(new_n451), .C1(new_n783), .C2(new_n450), .ZN(new_n816));
  NOR4_X1   g0616(.A1(new_n813), .A2(new_n814), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G294), .ZN(new_n818));
  INV_X1    g0618(.A(G303), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n817), .B1(new_n818), .B2(new_n745), .C1(new_n819), .C2(new_n756), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n738), .A2(G150), .B1(G143), .B2(new_n744), .ZN(new_n821));
  INV_X1    g0621(.A(G137), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n821), .B1(new_n822), .B2(new_n756), .C1(new_n328), .C2(new_n772), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT34), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n780), .A2(G68), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n825), .B(new_n257), .C1(new_n217), .C2(new_n749), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n769), .B2(G132), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n824), .B(new_n827), .C1(new_n777), .C2(new_n783), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n809), .B1(new_n820), .B2(new_n828), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n808), .A2(new_n800), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n719), .A2(new_n715), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n830), .B1(G77), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n685), .B(new_n806), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(new_n710), .Z(new_n835));
  OAI21_X1  g0635(.A(new_n833), .B1(new_n835), .B2(new_n734), .ZN(G384));
  INV_X1    g0636(.A(KEYINPUT35), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n233), .B1(new_n529), .B2(new_n837), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n838), .B(G116), .C1(new_n837), .C2(new_n529), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT36), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n325), .A2(G50), .A3(G77), .A4(new_n235), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(G50), .B2(new_n790), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(G1), .A3(new_n497), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n315), .A2(new_n637), .ZN(new_n844));
  AND3_X1   g0644(.A1(new_n330), .A2(new_n333), .A3(new_n340), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n342), .B1(KEYINPUT16), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n635), .B1(new_n846), .B2(new_n355), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n383), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n635), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n378), .B1(new_n381), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n365), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT37), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n846), .A2(new_n355), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n381), .B2(new_n849), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n855), .A2(KEYINPUT37), .A3(new_n365), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n848), .A2(KEYINPUT38), .A3(new_n853), .A4(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT39), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT38), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n369), .A2(new_n635), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n383), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT104), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT104), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n383), .A2(new_n864), .A3(new_n861), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n347), .A2(new_n355), .B1(new_n374), .B2(new_n635), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT37), .B1(new_n866), .B2(KEYINPUT103), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n851), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n850), .A2(KEYINPUT103), .A3(new_n365), .A4(KEYINPUT37), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n863), .A2(new_n865), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n859), .B1(new_n860), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n848), .A2(new_n853), .A3(new_n856), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n860), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n858), .B1(new_n874), .B2(new_n857), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n872), .A2(new_n875), .A3(KEYINPUT105), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT105), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n871), .A2(new_n860), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n857), .A2(new_n858), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n857), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n383), .A2(new_n847), .B1(new_n852), .B2(new_n851), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT38), .B1(new_n882), .B2(new_n856), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT39), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n877), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n844), .B1(new_n876), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n605), .A2(new_n849), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n881), .A2(new_n883), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n803), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(new_n685), .B2(new_n807), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n314), .A2(new_n637), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n315), .A2(new_n320), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n285), .A2(new_n314), .A3(new_n637), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n887), .B1(new_n889), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n886), .A2(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n685), .A2(new_n686), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n682), .B1(new_n681), .B2(new_n659), .ZN(new_n900));
  AOI211_X1 g0700(.A(KEYINPUT91), .B(new_n637), .C1(new_n680), .C2(new_n626), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n899), .B1(new_n902), .B2(KEYINPUT29), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n903), .A2(new_n435), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n608), .A2(new_n430), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n898), .B(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n865), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n864), .B1(new_n383), .B2(new_n861), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n868), .A2(new_n869), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n857), .B1(new_n911), .B2(KEYINPUT38), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n806), .B1(new_n894), .B2(new_n893), .ZN(new_n913));
  INV_X1    g0713(.A(new_n707), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n704), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n703), .A2(KEYINPUT31), .A3(new_n637), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n915), .B(new_n916), .C1(new_n600), .C2(new_n637), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n912), .A2(new_n918), .A3(KEYINPUT40), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n913), .A2(new_n917), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n920), .B1(new_n888), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n434), .A2(new_n917), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n923), .B(new_n924), .Z(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(G330), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n907), .B(new_n926), .Z(new_n927));
  AOI21_X1  g0727(.A(new_n205), .B1(G13), .B2(new_n206), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n840), .B(new_n843), .C1(new_n927), .C2(new_n928), .ZN(G367));
  NAND2_X1  g0729(.A1(new_n624), .A2(new_n637), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n538), .A2(new_n637), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n552), .A2(new_n555), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n654), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n637), .B1(new_n584), .B2(new_n594), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n936), .A2(KEYINPUT42), .A3(new_n658), .A4(new_n933), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n643), .A2(new_n658), .A3(new_n933), .A4(new_n659), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT42), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n555), .B1(new_n932), .B2(new_n590), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n659), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT106), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n670), .A2(new_n659), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n613), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n622), .B2(new_n946), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n944), .A2(new_n945), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n948), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n937), .A2(new_n940), .B1(new_n659), .B2(new_n942), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n950), .B1(new_n951), .B2(KEYINPUT106), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n953));
  AND3_X1   g0753(.A1(new_n949), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT43), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n949), .B2(new_n952), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n935), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n948), .B1(new_n944), .B2(new_n945), .ZN(new_n958));
  NOR3_X1   g0758(.A1(new_n951), .A2(KEYINPUT106), .A3(new_n950), .ZN(new_n959));
  OAI21_X1  g0759(.A(KEYINPUT43), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n935), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n949), .A2(new_n952), .A3(new_n953), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n957), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n663), .B(KEYINPUT41), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n660), .A2(new_n655), .A3(new_n933), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT45), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n660), .A2(KEYINPUT45), .A3(new_n655), .A4(new_n933), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n660), .A2(new_n655), .ZN(new_n972));
  XOR2_X1   g0772(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n973));
  NAND3_X1  g0773(.A1(new_n972), .A2(new_n934), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n934), .ZN(new_n975));
  INV_X1    g0775(.A(new_n973), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n971), .A2(new_n974), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n654), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(KEYINPUT108), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n660), .B1(new_n936), .B2(new_n653), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n982), .A2(G330), .A3(new_n644), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n652), .A2(new_n590), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n655), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n643), .A2(new_n659), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n799), .A2(new_n987), .A3(new_n660), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n983), .A2(new_n988), .ZN(new_n989));
  AND4_X1   g0789(.A1(new_n710), .A2(new_n684), .A3(new_n687), .A4(new_n989), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n971), .A2(new_n977), .A3(new_n654), .A4(new_n974), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT108), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n978), .A2(new_n992), .A3(new_n979), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n981), .A2(new_n990), .A3(new_n991), .A4(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n966), .B1(new_n994), .B2(new_n712), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n964), .B1(new_n995), .B2(new_n733), .ZN(new_n996));
  INV_X1    g0796(.A(G317), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n336), .B1(new_n756), .B2(new_n810), .C1(new_n767), .C2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(new_n512), .B2(new_n738), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n749), .A2(new_n219), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT46), .Z(new_n1001));
  NOR2_X1   g0801(.A1(new_n765), .A2(new_n450), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G107), .B2(new_n754), .ZN(new_n1003));
  AND3_X1   g0803(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n819), .B2(new_n745), .C1(new_n772), .C2(new_n812), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n783), .A2(new_n790), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(G150), .B2(new_n744), .ZN(new_n1007));
  INV_X1    g0807(.A(G143), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1007), .B1(new_n1008), .B2(new_n756), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT109), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n765), .A2(new_n389), .B1(new_n777), .B2(new_n749), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n1010), .A2(new_n336), .A3(new_n1011), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n217), .B2(new_n772), .C1(new_n328), .C2(new_n739), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n767), .A2(new_n822), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1005), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n1016));
  XNOR2_X1  g0816(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n719), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n726), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n722), .B1(new_n228), .B2(new_n386), .C1(new_n246), .C2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n950), .A2(new_n717), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1018), .A2(new_n734), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n996), .A2(new_n1022), .ZN(G387));
  INV_X1    g0823(.A(new_n989), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n711), .A2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n684), .A2(new_n989), .A3(new_n710), .A4(new_n687), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1025), .A2(new_n663), .A3(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n738), .A2(G311), .B1(G317), .B2(new_n744), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n819), .B2(new_n772), .C1(new_n741), .C2(new_n756), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT48), .Z(new_n1030));
  NOR2_X1   g0830(.A1(new_n783), .A2(new_n812), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n750), .A2(new_n512), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1033), .A2(KEYINPUT49), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1033), .A2(KEYINPUT49), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n336), .B1(new_n767), .B2(new_n757), .C1(new_n219), .C2(new_n765), .ZN(new_n1036));
  OR3_X1    g0836(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n767), .A2(new_n407), .B1(new_n389), .B2(new_n749), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT111), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n439), .A2(new_n754), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(new_n328), .C2(new_n756), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1041), .A2(new_n336), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n772), .A2(new_n790), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1043), .B(new_n1002), .C1(G50), .C2(new_n744), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1042), .B(new_n1044), .C1(new_n354), .C2(new_n739), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n809), .B1(new_n1037), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n726), .B1(new_n243), .B2(new_n468), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n665), .B2(new_n723), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n390), .A2(G50), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT50), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1050), .B(new_n468), .C1(new_n790), .C2(new_n389), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n665), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1048), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n662), .A2(new_n451), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n721), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1046), .A2(new_n800), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n985), .A2(new_n717), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1056), .A2(new_n1057), .B1(new_n733), .B2(new_n989), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1027), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT112), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1027), .A2(new_n1058), .A3(KEYINPUT112), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(G393));
  AND3_X1   g0863(.A1(new_n978), .A2(new_n992), .A3(new_n979), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n992), .B1(new_n978), .B2(new_n979), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n991), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1026), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n980), .A2(new_n991), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1066), .A2(new_n1068), .B1(new_n1026), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n663), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n980), .A2(new_n733), .A3(new_n991), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n810), .A2(new_n745), .B1(new_n756), .B2(new_n997), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT52), .Z(new_n1074));
  NOR2_X1   g0874(.A1(new_n1074), .A2(new_n257), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n819), .B2(new_n739), .C1(new_n749), .C2(new_n812), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n783), .A2(new_n219), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n767), .A2(new_n741), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n765), .A2(new_n451), .B1(new_n818), .B2(new_n772), .ZN(new_n1079));
  NOR4_X1   g0879(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n756), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1081), .A2(G150), .B1(G159), .B2(new_n744), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT51), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n783), .A2(new_n389), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n224), .B2(new_n750), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1085), .B(new_n257), .C1(new_n390), .C2(new_n772), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n739), .A2(new_n217), .B1(new_n1008), .B2(new_n767), .ZN(new_n1087));
  NOR4_X1   g0887(.A1(new_n1083), .A2(new_n1086), .A3(new_n814), .A4(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n719), .B1(new_n1080), .B2(new_n1088), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n722), .B1(new_n450), .B2(new_n228), .C1(new_n254), .C2(new_n1019), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT113), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n934), .A2(new_n717), .B1(new_n1091), .B2(new_n1090), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1089), .A2(new_n734), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1072), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(KEYINPUT114), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT114), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1072), .A2(new_n1097), .A3(new_n1094), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1071), .A2(new_n1099), .ZN(G390));
  OAI21_X1  g0900(.A(KEYINPUT105), .B1(new_n872), .B2(new_n875), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n880), .A2(new_n877), .A3(new_n884), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1101), .A2(new_n1102), .A3(new_n715), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n780), .A2(G50), .B1(G132), .B2(new_n744), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1081), .A2(G128), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1104), .B(new_n1105), .C1(new_n328), .C2(new_n783), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n750), .A2(G150), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT53), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(KEYINPUT54), .B(G143), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n772), .A2(new_n1109), .ZN(new_n1110));
  NOR4_X1   g0910(.A1(new_n1106), .A2(new_n336), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(G125), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n1111), .B1(new_n1112), .B2(new_n768), .C1(new_n822), .C2(new_n739), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT116), .Z(new_n1114));
  OAI22_X1  g0914(.A1(new_n739), .A2(new_n451), .B1(new_n761), .B2(new_n756), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n769), .B2(G294), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n787), .B(new_n1084), .C1(G97), .C2(new_n773), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n825), .A3(new_n1117), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n257), .B(new_n1118), .C1(G116), .C2(new_n744), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n719), .B1(new_n1114), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n831), .A2(new_n354), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1103), .A2(new_n734), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n1122), .A2(KEYINPUT117), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(KEYINPUT117), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n844), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n891), .B2(new_n895), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1101), .A2(new_n1102), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n678), .A2(new_n683), .A3(new_n803), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n805), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n912), .B(new_n1125), .C1(new_n1129), .C2(new_n895), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT115), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n913), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1131), .B1(new_n1132), .B2(new_n710), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n913), .A2(new_n709), .A3(KEYINPUT115), .A4(G330), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1127), .A2(new_n1130), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n913), .A2(G330), .A3(new_n917), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n733), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1123), .B(new_n1124), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n609), .B1(new_n924), .B2(new_n795), .C1(new_n435), .C2(new_n903), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n917), .A2(G330), .A3(new_n807), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1128), .A2(new_n805), .B1(new_n1145), .B2(new_n895), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n895), .B1(new_n710), .B2(new_n806), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n1138), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n891), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1135), .A2(new_n1146), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1144), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1150), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n924), .A2(new_n795), .ZN(new_n1154));
  NOR3_X1   g0954(.A1(new_n904), .A2(new_n1154), .A3(new_n905), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n664), .B1(new_n1141), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1143), .B1(new_n1152), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(G378));
  NAND3_X1  g0959(.A1(new_n919), .A2(G330), .A3(new_n922), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n886), .A2(new_n897), .A3(new_n1160), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n919), .A2(G330), .A3(new_n922), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1125), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n897), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1162), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n607), .A2(new_n430), .ZN(new_n1166));
  XOR2_X1   g0966(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT119), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1166), .B(new_n1168), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n413), .A2(new_n849), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1169), .B(new_n1170), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n1161), .A2(new_n1165), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1171), .B1(new_n1161), .B2(new_n1165), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1172), .A2(new_n1173), .A3(new_n1142), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1171), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n715), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n756), .A2(new_n219), .B1(new_n389), .B2(new_n749), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n780), .A2(G58), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT118), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1177), .B(new_n1179), .C1(G283), .C2(new_n769), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n264), .B(new_n336), .C1(new_n739), .C2(new_n450), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1006), .B(new_n1181), .C1(new_n439), .C2(new_n773), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1180), .B(new_n1182), .C1(new_n451), .C2(new_n745), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT58), .Z(new_n1184));
  OAI21_X1  g0984(.A(new_n217), .B1(new_n334), .B2(G41), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n756), .A2(new_n1112), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n773), .A2(G137), .B1(new_n744), .B2(G128), .ZN(new_n1187));
  INV_X1    g0987(.A(G132), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1187), .B1(new_n749), .B2(new_n1109), .C1(new_n739), .C2(new_n1188), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1186), .B(new_n1189), .C1(G150), .C2(new_n754), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT59), .ZN(new_n1191));
  AOI21_X1  g0991(.A(G33), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n767), .ZN(new_n1193));
  AOI21_X1  g0993(.A(G41), .B1(new_n1193), .B2(G124), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1192), .B(new_n1194), .C1(new_n328), .C2(new_n765), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1185), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n719), .B1(new_n1184), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n831), .A2(new_n217), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1176), .A2(new_n734), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1174), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1161), .A2(new_n1165), .A3(new_n1171), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1160), .B1(new_n886), .B2(new_n897), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1175), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1203), .A2(KEYINPUT57), .A3(new_n1204), .A4(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n663), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1210));
  AOI21_X1  g1010(.A(KEYINPUT57), .B1(new_n1210), .B2(new_n1203), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1202), .B1(new_n1209), .B2(new_n1211), .ZN(G375));
  OAI21_X1  g1012(.A(new_n734), .B1(G68), .B2(new_n832), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT120), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n769), .A2(G128), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n257), .B1(new_n756), .B2(new_n1188), .C1(new_n739), .C2(new_n1109), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n745), .A2(new_n822), .B1(new_n407), .B2(new_n772), .ZN(new_n1217));
  NOR4_X1   g1017(.A1(new_n1215), .A2(new_n1179), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n217), .B2(new_n783), .C1(new_n328), .C2(new_n749), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n768), .A2(new_n819), .B1(new_n450), .B2(new_n749), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT121), .Z(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G294), .B2(new_n1081), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n738), .A2(G116), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n780), .A2(G77), .B1(G283), .B2(new_n744), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1222), .A2(new_n1040), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n336), .B1(new_n772), .B2(new_n451), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1219), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1227), .A2(new_n719), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1214), .B(new_n1228), .C1(new_n715), .C2(new_n895), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1153), .B2(new_n733), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1144), .A2(new_n1150), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n965), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1230), .B1(new_n1232), .B2(new_n1151), .ZN(G381));
  INV_X1    g1033(.A(KEYINPUT57), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1207), .A2(new_n1204), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1127), .A2(new_n1130), .A3(new_n1136), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1236), .B1(new_n1237), .B2(new_n1139), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1144), .B1(new_n1238), .B2(new_n1151), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1234), .B1(new_n1235), .B2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1240), .A2(new_n663), .A3(new_n1208), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1241), .A2(new_n1158), .A3(new_n1202), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1070), .A2(new_n663), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n996), .A2(new_n1243), .A3(new_n1022), .ZN(new_n1244));
  INV_X1    g1044(.A(G396), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1061), .A2(new_n1245), .A3(new_n1062), .ZN(new_n1246));
  NOR4_X1   g1046(.A1(new_n1244), .A2(G381), .A3(G384), .A4(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1242), .A2(new_n1247), .ZN(G407));
  NAND3_X1  g1048(.A1(new_n1241), .A2(new_n1158), .A3(new_n1202), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1247), .A2(new_n636), .ZN(new_n1250));
  OAI21_X1  g1050(.A(G213), .B1(new_n1249), .B2(new_n1250), .ZN(G409));
  AND3_X1   g1051(.A1(new_n1027), .A2(KEYINPUT112), .A3(new_n1058), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT112), .B1(new_n1027), .B2(new_n1058), .ZN(new_n1253));
  OAI21_X1  g1053(.A(G396), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1254), .A2(new_n1246), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT126), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1255), .B1(new_n1256), .B2(G387), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1022), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n903), .A2(new_n710), .A3(new_n989), .A4(new_n991), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1259), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n965), .B1(new_n1260), .B2(new_n711), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1142), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1258), .B1(new_n1262), .B2(new_n964), .ZN(new_n1263));
  OAI211_X1 g1063(.A(KEYINPUT126), .B(G390), .C1(new_n1263), .C2(KEYINPUT125), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT125), .B1(new_n996), .B2(new_n1022), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1243), .B1(new_n1265), .B2(new_n1256), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1257), .A2(new_n1264), .A3(new_n1266), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n996), .A2(new_n1243), .A3(new_n1022), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1243), .B1(new_n996), .B2(new_n1022), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT124), .B1(new_n1270), .B2(new_n1255), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n957), .A2(new_n963), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n1261), .B2(new_n1142), .ZN(new_n1273));
  OAI21_X1  g1073(.A(G390), .B1(new_n1273), .B2(new_n1258), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1274), .A2(KEYINPUT124), .A3(new_n1255), .A4(new_n1244), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1267), .B1(new_n1271), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(KEYINPUT127), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1274), .A2(new_n1244), .A3(new_n1255), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT124), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1275), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT127), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1282), .A2(new_n1283), .A3(new_n1267), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1278), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT60), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1231), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1144), .A2(new_n1150), .A3(KEYINPUT60), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1287), .A2(new_n663), .A3(new_n1156), .A4(new_n1288), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1289), .A2(G384), .A3(new_n1230), .ZN(new_n1290));
  AOI21_X1  g1090(.A(G384), .B1(new_n1289), .B2(new_n1230), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT123), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1290), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1292), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n636), .A2(G213), .ZN(new_n1295));
  INV_X1    g1095(.A(G2897), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1294), .A2(new_n1297), .ZN(new_n1298));
  OAI221_X1 g1098(.A(new_n1292), .B1(new_n1296), .B2(new_n1295), .C1(new_n1290), .C2(new_n1291), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1293), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(KEYINPUT122), .B1(new_n1174), .B2(new_n1201), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT122), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1302), .B(new_n1200), .C1(new_n1235), .C2(new_n1142), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1210), .A2(new_n965), .A3(new_n1203), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1301), .A2(new_n1158), .A3(new_n1303), .A4(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1295), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1158), .B1(new_n1241), .B2(new_n1202), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1300), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n1306), .A2(new_n1307), .A3(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT62), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1308), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT61), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(G375), .A2(G378), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1315), .A2(new_n1309), .A3(new_n1295), .A4(new_n1305), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1314), .B1(new_n1316), .B2(KEYINPUT62), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1285), .B1(new_n1313), .B2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(KEYINPUT61), .B1(new_n1282), .B2(new_n1267), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1311), .A2(KEYINPUT63), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT63), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1315), .A2(new_n1295), .A3(new_n1305), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1321), .B1(new_n1322), .B2(new_n1300), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n1319), .B(new_n1320), .C1(new_n1323), .C2(new_n1311), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1318), .A2(new_n1324), .ZN(G405));
  NOR2_X1   g1125(.A1(new_n1242), .A2(new_n1307), .ZN(new_n1326));
  AND3_X1   g1126(.A1(new_n1282), .A2(new_n1283), .A3(new_n1267), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1283), .B1(new_n1282), .B2(new_n1267), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1326), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1315), .A2(new_n1249), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1278), .A2(new_n1284), .A3(new_n1330), .ZN(new_n1331));
  AND3_X1   g1131(.A1(new_n1329), .A2(new_n1309), .A3(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1309), .B1(new_n1329), .B2(new_n1331), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1332), .A2(new_n1333), .ZN(G402));
endmodule


