

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579;

  NOR2_X1 U322 ( .A1(n564), .A2(n395), .ZN(n396) );
  XNOR2_X1 U323 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n404) );
  XNOR2_X1 U324 ( .A(n405), .B(n404), .ZN(n533) );
  NOR2_X1 U325 ( .A1(n505), .A2(n441), .ZN(n555) );
  XOR2_X1 U326 ( .A(n548), .B(KEYINPUT77), .Z(n557) );
  XNOR2_X1 U327 ( .A(n442), .B(G176GAT), .ZN(n443) );
  XNOR2_X1 U328 ( .A(n444), .B(n443), .ZN(G1349GAT) );
  XOR2_X1 U329 ( .A(G176GAT), .B(KEYINPUT72), .Z(n411) );
  XOR2_X1 U330 ( .A(KEYINPUT31), .B(n411), .Z(n293) );
  XOR2_X1 U331 ( .A(G64GAT), .B(KEYINPUT13), .Z(n291) );
  XNOR2_X1 U332 ( .A(G71GAT), .B(G57GAT), .ZN(n290) );
  XNOR2_X1 U333 ( .A(n291), .B(n290), .ZN(n366) );
  XNOR2_X1 U334 ( .A(G120GAT), .B(n366), .ZN(n292) );
  XNOR2_X1 U335 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U336 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n295) );
  NAND2_X1 U337 ( .A1(G230GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U338 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U339 ( .A(n297), .B(n296), .Z(n302) );
  XOR2_X1 U340 ( .A(KEYINPUT71), .B(G92GAT), .Z(n299) );
  XNOR2_X1 U341 ( .A(G99GAT), .B(G85GAT), .ZN(n298) );
  XNOR2_X1 U342 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U343 ( .A(G106GAT), .B(n300), .Z(n390) );
  XNOR2_X1 U344 ( .A(n390), .B(KEYINPUT33), .ZN(n301) );
  XNOR2_X1 U345 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U346 ( .A(KEYINPUT69), .B(G204GAT), .Z(n304) );
  XNOR2_X1 U347 ( .A(G148GAT), .B(G78GAT), .ZN(n303) );
  XNOR2_X1 U348 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U349 ( .A(KEYINPUT70), .B(n305), .ZN(n344) );
  XNOR2_X1 U350 ( .A(n306), .B(n344), .ZN(n570) );
  XNOR2_X1 U351 ( .A(KEYINPUT41), .B(n570), .ZN(n539) );
  XNOR2_X1 U352 ( .A(KEYINPUT104), .B(n539), .ZN(n517) );
  XOR2_X1 U353 ( .A(G71GAT), .B(G176GAT), .Z(n308) );
  XNOR2_X1 U354 ( .A(G15GAT), .B(KEYINPUT82), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U356 ( .A(KEYINPUT83), .B(KEYINPUT87), .Z(n310) );
  XNOR2_X1 U357 ( .A(KEYINPUT86), .B(KEYINPUT84), .ZN(n309) );
  XNOR2_X1 U358 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U359 ( .A(n312), .B(n311), .Z(n325) );
  XOR2_X1 U360 ( .A(KEYINPUT81), .B(KEYINPUT0), .Z(n314) );
  XNOR2_X1 U361 ( .A(G134GAT), .B(KEYINPUT80), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U363 ( .A(n315), .B(G127GAT), .Z(n317) );
  XNOR2_X1 U364 ( .A(G113GAT), .B(G120GAT), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n317), .B(n316), .ZN(n425) );
  XOR2_X1 U366 ( .A(KEYINPUT20), .B(G99GAT), .Z(n319) );
  XNOR2_X1 U367 ( .A(G43GAT), .B(G190GAT), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U369 ( .A(G183GAT), .B(n320), .Z(n322) );
  NAND2_X1 U370 ( .A1(G227GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U372 ( .A(n425), .B(n323), .ZN(n324) );
  XNOR2_X1 U373 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U374 ( .A(KEYINPUT17), .B(KEYINPUT85), .Z(n327) );
  XNOR2_X1 U375 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n326) );
  XNOR2_X1 U376 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U377 ( .A(G169GAT), .B(n328), .ZN(n419) );
  XOR2_X1 U378 ( .A(n329), .B(n419), .Z(n514) );
  INV_X1 U379 ( .A(n514), .ZN(n505) );
  XOR2_X1 U380 ( .A(KEYINPUT22), .B(KEYINPUT89), .Z(n331) );
  NAND2_X1 U381 ( .A1(G228GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U382 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U383 ( .A(n332), .B(KEYINPUT24), .Z(n337) );
  XNOR2_X1 U384 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n333) );
  XNOR2_X1 U385 ( .A(n333), .B(KEYINPUT2), .ZN(n428) );
  XOR2_X1 U386 ( .A(G211GAT), .B(KEYINPUT21), .Z(n335) );
  XNOR2_X1 U387 ( .A(G197GAT), .B(KEYINPUT88), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n414) );
  XNOR2_X1 U389 ( .A(n428), .B(n414), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U391 ( .A(KEYINPUT90), .B(KEYINPUT23), .Z(n339) );
  XNOR2_X1 U392 ( .A(G218GAT), .B(G106GAT), .ZN(n338) );
  XNOR2_X1 U393 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U394 ( .A(n341), .B(n340), .Z(n343) );
  XOR2_X1 U395 ( .A(G50GAT), .B(G162GAT), .Z(n378) );
  XOR2_X1 U396 ( .A(G22GAT), .B(G155GAT), .Z(n365) );
  XNOR2_X1 U397 ( .A(n378), .B(n365), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n343), .B(n342), .ZN(n345) );
  XNOR2_X1 U399 ( .A(n345), .B(n344), .ZN(n452) );
  XOR2_X1 U400 ( .A(G197GAT), .B(G141GAT), .Z(n347) );
  XNOR2_X1 U401 ( .A(G169GAT), .B(G22GAT), .ZN(n346) );
  XNOR2_X1 U402 ( .A(n347), .B(n346), .ZN(n362) );
  XOR2_X1 U403 ( .A(G15GAT), .B(G1GAT), .Z(n373) );
  XOR2_X1 U404 ( .A(n373), .B(G50GAT), .Z(n351) );
  XOR2_X1 U405 ( .A(G29GAT), .B(G43GAT), .Z(n349) );
  XNOR2_X1 U406 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n379) );
  XNOR2_X1 U408 ( .A(G36GAT), .B(n379), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U410 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n353) );
  NAND2_X1 U411 ( .A1(G229GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U412 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U413 ( .A(n355), .B(n354), .Z(n360) );
  XOR2_X1 U414 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n357) );
  XNOR2_X1 U415 ( .A(G113GAT), .B(KEYINPUT30), .ZN(n356) );
  XNOR2_X1 U416 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n358), .B(G8GAT), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U419 ( .A(n362), .B(n361), .ZN(n536) );
  INV_X1 U420 ( .A(n536), .ZN(n564) );
  XOR2_X1 U421 ( .A(KEYINPUT12), .B(G211GAT), .Z(n364) );
  XNOR2_X1 U422 ( .A(G127GAT), .B(G78GAT), .ZN(n363) );
  XNOR2_X1 U423 ( .A(n364), .B(n363), .ZN(n377) );
  XOR2_X1 U424 ( .A(n366), .B(n365), .Z(n368) );
  NAND2_X1 U425 ( .A1(G231GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U426 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U427 ( .A(KEYINPUT78), .B(KEYINPUT15), .Z(n370) );
  XNOR2_X1 U428 ( .A(KEYINPUT14), .B(KEYINPUT79), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U430 ( .A(n372), .B(n371), .Z(n375) );
  XOR2_X1 U431 ( .A(G8GAT), .B(G183GAT), .Z(n413) );
  XNOR2_X1 U432 ( .A(n373), .B(n413), .ZN(n374) );
  XNOR2_X1 U433 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U434 ( .A(n377), .B(n376), .ZN(n574) );
  INV_X1 U435 ( .A(n574), .ZN(n397) );
  XOR2_X1 U436 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n381) );
  XNOR2_X1 U437 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U438 ( .A(n381), .B(n380), .ZN(n386) );
  XNOR2_X1 U439 ( .A(G36GAT), .B(G190GAT), .ZN(n382) );
  XNOR2_X1 U440 ( .A(n382), .B(G218GAT), .ZN(n408) );
  XOR2_X1 U441 ( .A(n408), .B(KEYINPUT65), .Z(n384) );
  NAND2_X1 U442 ( .A1(G232GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U444 ( .A(n386), .B(n385), .Z(n392) );
  XOR2_X1 U445 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n388) );
  XNOR2_X1 U446 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n387) );
  XNOR2_X1 U447 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U449 ( .A(n392), .B(n391), .ZN(n548) );
  XNOR2_X1 U450 ( .A(KEYINPUT36), .B(n557), .ZN(n577) );
  NOR2_X1 U451 ( .A1(n397), .A2(n577), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n393), .B(KEYINPUT45), .ZN(n394) );
  NAND2_X1 U453 ( .A1(n394), .A2(n570), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(KEYINPUT111), .ZN(n403) );
  XOR2_X1 U455 ( .A(KEYINPUT110), .B(n397), .Z(n552) );
  NAND2_X1 U456 ( .A1(n564), .A2(n539), .ZN(n398) );
  XNOR2_X1 U457 ( .A(KEYINPUT46), .B(n398), .ZN(n399) );
  NAND2_X1 U458 ( .A1(n399), .A2(n548), .ZN(n400) );
  NOR2_X1 U459 ( .A1(n552), .A2(n400), .ZN(n401) );
  XNOR2_X1 U460 ( .A(KEYINPUT47), .B(n401), .ZN(n402) );
  AND2_X1 U461 ( .A1(n403), .A2(n402), .ZN(n405) );
  XOR2_X1 U462 ( .A(KEYINPUT93), .B(G64GAT), .Z(n407) );
  XNOR2_X1 U463 ( .A(G204GAT), .B(G92GAT), .ZN(n406) );
  XNOR2_X1 U464 ( .A(n407), .B(n406), .ZN(n418) );
  XOR2_X1 U465 ( .A(n408), .B(KEYINPUT94), .Z(n410) );
  NAND2_X1 U466 ( .A1(G226GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n410), .B(n409), .ZN(n412) );
  XOR2_X1 U468 ( .A(n412), .B(n411), .Z(n416) );
  XNOR2_X1 U469 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U470 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U471 ( .A(n418), .B(n417), .ZN(n420) );
  XNOR2_X1 U472 ( .A(n420), .B(n419), .ZN(n503) );
  NOR2_X1 U473 ( .A1(n533), .A2(n503), .ZN(n421) );
  XNOR2_X1 U474 ( .A(n421), .B(KEYINPUT54), .ZN(n439) );
  XOR2_X1 U475 ( .A(KEYINPUT5), .B(G57GAT), .Z(n423) );
  XNOR2_X1 U476 ( .A(KEYINPUT4), .B(KEYINPUT92), .ZN(n422) );
  XNOR2_X1 U477 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n425), .B(n424), .ZN(n438) );
  XOR2_X1 U479 ( .A(G85GAT), .B(G155GAT), .Z(n427) );
  XNOR2_X1 U480 ( .A(G29GAT), .B(G162GAT), .ZN(n426) );
  XNOR2_X1 U481 ( .A(n427), .B(n426), .ZN(n436) );
  XOR2_X1 U482 ( .A(n428), .B(G1GAT), .Z(n430) );
  NAND2_X1 U483 ( .A1(G225GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U485 ( .A(KEYINPUT1), .B(KEYINPUT91), .Z(n432) );
  XNOR2_X1 U486 ( .A(G148GAT), .B(KEYINPUT6), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U488 ( .A(n434), .B(n433), .Z(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n438), .B(n437), .ZN(n532) );
  NAND2_X1 U491 ( .A1(n439), .A2(n532), .ZN(n562) );
  NOR2_X1 U492 ( .A1(n452), .A2(n562), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n440), .B(KEYINPUT55), .ZN(n441) );
  NAND2_X1 U494 ( .A1(n517), .A2(n555), .ZN(n444) );
  XOR2_X1 U495 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n442) );
  NAND2_X1 U496 ( .A1(n452), .A2(n505), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n445), .B(KEYINPUT26), .ZN(n563) );
  XNOR2_X1 U498 ( .A(KEYINPUT27), .B(n503), .ZN(n454) );
  NOR2_X1 U499 ( .A1(n563), .A2(n454), .ZN(n535) );
  XOR2_X1 U500 ( .A(n535), .B(KEYINPUT96), .Z(n450) );
  NOR2_X1 U501 ( .A1(n505), .A2(n503), .ZN(n446) );
  XOR2_X1 U502 ( .A(KEYINPUT97), .B(n446), .Z(n447) );
  NOR2_X1 U503 ( .A1(n452), .A2(n447), .ZN(n448) );
  XNOR2_X1 U504 ( .A(KEYINPUT25), .B(n448), .ZN(n449) );
  NAND2_X1 U505 ( .A1(n450), .A2(n449), .ZN(n451) );
  NAND2_X1 U506 ( .A1(n532), .A2(n451), .ZN(n459) );
  XOR2_X1 U507 ( .A(n452), .B(KEYINPUT28), .Z(n508) );
  INV_X1 U508 ( .A(n508), .ZN(n453) );
  NOR2_X1 U509 ( .A1(n532), .A2(n453), .ZN(n456) );
  INV_X1 U510 ( .A(n454), .ZN(n455) );
  NAND2_X1 U511 ( .A1(n456), .A2(n455), .ZN(n512) );
  XNOR2_X1 U512 ( .A(KEYINPUT95), .B(n512), .ZN(n457) );
  NAND2_X1 U513 ( .A1(n457), .A2(n505), .ZN(n458) );
  NAND2_X1 U514 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U515 ( .A(n460), .B(KEYINPUT98), .ZN(n475) );
  NAND2_X1 U516 ( .A1(n557), .A2(n574), .ZN(n461) );
  XOR2_X1 U517 ( .A(KEYINPUT16), .B(n461), .Z(n462) );
  AND2_X1 U518 ( .A1(n475), .A2(n462), .ZN(n489) );
  NAND2_X1 U519 ( .A1(n570), .A2(n564), .ZN(n463) );
  XOR2_X1 U520 ( .A(KEYINPUT74), .B(n463), .Z(n477) );
  NAND2_X1 U521 ( .A1(n489), .A2(n477), .ZN(n471) );
  NOR2_X1 U522 ( .A1(n532), .A2(n471), .ZN(n464) );
  XOR2_X1 U523 ( .A(KEYINPUT34), .B(n464), .Z(n465) );
  XNOR2_X1 U524 ( .A(G1GAT), .B(n465), .ZN(G1324GAT) );
  NOR2_X1 U525 ( .A1(n503), .A2(n471), .ZN(n467) );
  XNOR2_X1 U526 ( .A(G8GAT), .B(KEYINPUT99), .ZN(n466) );
  XNOR2_X1 U527 ( .A(n467), .B(n466), .ZN(G1325GAT) );
  NOR2_X1 U528 ( .A1(n505), .A2(n471), .ZN(n469) );
  XNOR2_X1 U529 ( .A(KEYINPUT35), .B(KEYINPUT100), .ZN(n468) );
  XNOR2_X1 U530 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U531 ( .A(G15GAT), .B(n470), .ZN(G1326GAT) );
  NOR2_X1 U532 ( .A1(n508), .A2(n471), .ZN(n473) );
  XNOR2_X1 U533 ( .A(G22GAT), .B(KEYINPUT101), .ZN(n472) );
  XNOR2_X1 U534 ( .A(n473), .B(n472), .ZN(G1327GAT) );
  NOR2_X1 U535 ( .A1(n574), .A2(n577), .ZN(n474) );
  NAND2_X1 U536 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X1 U537 ( .A(KEYINPUT37), .B(n476), .ZN(n501) );
  NAND2_X1 U538 ( .A1(n477), .A2(n501), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n478), .B(KEYINPUT38), .ZN(n486) );
  NOR2_X1 U540 ( .A1(n486), .A2(n532), .ZN(n481) );
  XNOR2_X1 U541 ( .A(G29GAT), .B(KEYINPUT102), .ZN(n479) );
  XNOR2_X1 U542 ( .A(n479), .B(KEYINPUT39), .ZN(n480) );
  XNOR2_X1 U543 ( .A(n481), .B(n480), .ZN(G1328GAT) );
  NOR2_X1 U544 ( .A1(n486), .A2(n503), .ZN(n483) );
  XNOR2_X1 U545 ( .A(G36GAT), .B(KEYINPUT103), .ZN(n482) );
  XNOR2_X1 U546 ( .A(n483), .B(n482), .ZN(G1329GAT) );
  NOR2_X1 U547 ( .A1(n505), .A2(n486), .ZN(n484) );
  XOR2_X1 U548 ( .A(KEYINPUT40), .B(n484), .Z(n485) );
  XNOR2_X1 U549 ( .A(G43GAT), .B(n485), .ZN(G1330GAT) );
  NOR2_X1 U550 ( .A1(n508), .A2(n486), .ZN(n487) );
  XOR2_X1 U551 ( .A(G50GAT), .B(n487), .Z(G1331GAT) );
  NAND2_X1 U552 ( .A1(n536), .A2(n517), .ZN(n488) );
  XNOR2_X1 U553 ( .A(n488), .B(KEYINPUT105), .ZN(n500) );
  NAND2_X1 U554 ( .A1(n500), .A2(n489), .ZN(n496) );
  NOR2_X1 U555 ( .A1(n532), .A2(n496), .ZN(n491) );
  XNOR2_X1 U556 ( .A(KEYINPUT42), .B(KEYINPUT106), .ZN(n490) );
  XNOR2_X1 U557 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U558 ( .A(G57GAT), .B(n492), .Z(G1332GAT) );
  NOR2_X1 U559 ( .A1(n503), .A2(n496), .ZN(n493) );
  XOR2_X1 U560 ( .A(G64GAT), .B(n493), .Z(G1333GAT) );
  NOR2_X1 U561 ( .A1(n505), .A2(n496), .ZN(n495) );
  XNOR2_X1 U562 ( .A(G71GAT), .B(KEYINPUT107), .ZN(n494) );
  XNOR2_X1 U563 ( .A(n495), .B(n494), .ZN(G1334GAT) );
  NOR2_X1 U564 ( .A1(n508), .A2(n496), .ZN(n498) );
  XNOR2_X1 U565 ( .A(KEYINPUT43), .B(KEYINPUT108), .ZN(n497) );
  XNOR2_X1 U566 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U567 ( .A(G78GAT), .B(n499), .ZN(G1335GAT) );
  NAND2_X1 U568 ( .A1(n501), .A2(n500), .ZN(n507) );
  NOR2_X1 U569 ( .A1(n532), .A2(n507), .ZN(n502) );
  XOR2_X1 U570 ( .A(G85GAT), .B(n502), .Z(G1336GAT) );
  NOR2_X1 U571 ( .A1(n503), .A2(n507), .ZN(n504) );
  XOR2_X1 U572 ( .A(G92GAT), .B(n504), .Z(G1337GAT) );
  NOR2_X1 U573 ( .A1(n505), .A2(n507), .ZN(n506) );
  XOR2_X1 U574 ( .A(G99GAT), .B(n506), .Z(G1338GAT) );
  NOR2_X1 U575 ( .A1(n508), .A2(n507), .ZN(n510) );
  XNOR2_X1 U576 ( .A(KEYINPUT44), .B(KEYINPUT109), .ZN(n509) );
  XNOR2_X1 U577 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U578 ( .A(G106GAT), .B(n511), .ZN(G1339GAT) );
  NOR2_X1 U579 ( .A1(n533), .A2(n512), .ZN(n513) );
  NAND2_X1 U580 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(KEYINPUT112), .B(n515), .ZN(n527) );
  INV_X1 U582 ( .A(n527), .ZN(n522) );
  NAND2_X1 U583 ( .A1(n564), .A2(n522), .ZN(n516) );
  XNOR2_X1 U584 ( .A(G113GAT), .B(n516), .ZN(G1340GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n519) );
  NAND2_X1 U586 ( .A1(n517), .A2(n522), .ZN(n518) );
  XNOR2_X1 U587 ( .A(n519), .B(n518), .ZN(n521) );
  XOR2_X1 U588 ( .A(G120GAT), .B(KEYINPUT113), .Z(n520) );
  XNOR2_X1 U589 ( .A(n521), .B(n520), .ZN(G1341GAT) );
  XNOR2_X1 U590 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n526) );
  XOR2_X1 U591 ( .A(KEYINPUT116), .B(KEYINPUT115), .Z(n524) );
  NAND2_X1 U592 ( .A1(n552), .A2(n522), .ZN(n523) );
  XNOR2_X1 U593 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U594 ( .A(n526), .B(n525), .ZN(G1342GAT) );
  NOR2_X1 U595 ( .A1(n527), .A2(n557), .ZN(n531) );
  XOR2_X1 U596 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n529) );
  XNOR2_X1 U597 ( .A(G134GAT), .B(KEYINPUT118), .ZN(n528) );
  XNOR2_X1 U598 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(G1343GAT) );
  NOR2_X1 U600 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n547) );
  NOR2_X1 U602 ( .A1(n536), .A2(n547), .ZN(n538) );
  XNOR2_X1 U603 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(G1344GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n541) );
  INV_X1 U606 ( .A(n547), .ZN(n545) );
  NAND2_X1 U607 ( .A1(n545), .A2(n539), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U609 ( .A(n542), .B(KEYINPUT52), .Z(n544) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(G1345GAT) );
  NAND2_X1 U612 ( .A1(n574), .A2(n545), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n546), .B(G155GAT), .ZN(G1346GAT) );
  NOR2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U615 ( .A(KEYINPUT122), .B(n549), .Z(n550) );
  XNOR2_X1 U616 ( .A(G162GAT), .B(n550), .ZN(G1347GAT) );
  NAND2_X1 U617 ( .A1(n564), .A2(n555), .ZN(n551) );
  XNOR2_X1 U618 ( .A(G169GAT), .B(n551), .ZN(G1348GAT) );
  XOR2_X1 U619 ( .A(G183GAT), .B(KEYINPUT123), .Z(n554) );
  NAND2_X1 U620 ( .A1(n555), .A2(n552), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1350GAT) );
  INV_X1 U622 ( .A(n555), .ZN(n556) );
  NOR2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n561) );
  XNOR2_X1 U624 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(KEYINPUT124), .ZN(n559) );
  XNOR2_X1 U626 ( .A(KEYINPUT125), .B(n559), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1351GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT127), .B(KEYINPUT60), .Z(n566) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n573) );
  NAND2_X1 U630 ( .A1(n573), .A2(n564), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(n567) );
  XOR2_X1 U632 ( .A(n567), .B(KEYINPUT59), .Z(n569) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .Z(n572) );
  INV_X1 U636 ( .A(n573), .ZN(n576) );
  OR2_X1 U637 ( .A1(n576), .A2(n570), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1353GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U642 ( .A(KEYINPUT62), .B(n578), .Z(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

