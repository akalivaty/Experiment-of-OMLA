//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n871, new_n872, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT31), .ZN(new_n188));
  XOR2_X1   g002(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G210), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n189), .B(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT26), .B(G101), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n193), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT68), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT67), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n197), .B1(G116), .B2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G116), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(new_n198), .ZN(new_n201));
  INV_X1    g015(.A(G116), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT66), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G116), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(new_n197), .A3(G119), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT2), .B(G113), .ZN(new_n208));
  AND3_X1   g022(.A1(new_n201), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n208), .B1(new_n201), .B2(new_n207), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n196), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n208), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT67), .B1(new_n202), .B2(G119), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n213), .B1(new_n206), .B2(G119), .ZN(new_n214));
  AOI211_X1 g028(.A(KEYINPUT67), .B(new_n198), .C1(new_n203), .C2(new_n205), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n212), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n201), .A2(new_n207), .A3(new_n208), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(KEYINPUT68), .A3(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n211), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n220));
  INV_X1    g034(.A(G143), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(G146), .ZN(new_n223));
  INV_X1    g037(.A(G146), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(KEYINPUT64), .A3(G143), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT1), .B1(new_n221), .B2(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G128), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(G143), .B(G146), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT11), .ZN(new_n235));
  INV_X1    g049(.A(G134), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(G137), .ZN(new_n237));
  INV_X1    g051(.A(G137), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT11), .A3(G134), .ZN(new_n239));
  INV_X1    g053(.A(G131), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n236), .A2(G137), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n237), .A2(new_n239), .A3(new_n240), .A4(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n238), .A2(G134), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n236), .A2(G137), .ZN(new_n244));
  OAI21_X1  g058(.A(G131), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT65), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n234), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n226), .A2(new_n228), .B1(new_n230), .B2(new_n232), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n242), .A2(new_n245), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT65), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n237), .A2(new_n241), .A3(new_n239), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G131), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n242), .ZN(new_n254));
  AND2_X1   g068(.A1(KEYINPUT0), .A2(G128), .ZN(new_n255));
  NOR2_X1   g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n226), .A2(new_n257), .B1(new_n230), .B2(new_n255), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n248), .A2(new_n251), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT30), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n234), .A2(new_n246), .A3(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT69), .B1(new_n249), .B2(new_n250), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n264), .A2(new_n265), .A3(new_n259), .A4(KEYINPUT30), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n219), .A2(new_n262), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n211), .A2(new_n218), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n264), .A2(new_n265), .A3(new_n259), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT70), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT70), .B1(new_n268), .B2(new_n269), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n195), .B(new_n267), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT72), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n264), .A2(new_n265), .A3(new_n259), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n274), .B1(new_n219), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT70), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n278), .A2(new_n279), .A3(new_n195), .A4(new_n267), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n188), .B1(new_n273), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n219), .A2(new_n260), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n282), .B1(new_n270), .B2(new_n271), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT28), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n234), .A2(new_n246), .B1(new_n254), .B2(new_n258), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT28), .B1(new_n268), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n195), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n272), .A2(KEYINPUT31), .ZN(new_n289));
  NOR3_X1   g103(.A1(new_n281), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(G472), .A2(G902), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n187), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n273), .A2(new_n280), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT31), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n284), .A2(new_n287), .ZN(new_n296));
  INV_X1    g110(.A(new_n195), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n289), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n295), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(KEYINPUT32), .A3(new_n291), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n293), .A2(KEYINPUT73), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n291), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(new_n187), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n278), .A2(new_n267), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n297), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT29), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n308), .B(new_n309), .C1(new_n296), .C2(new_n297), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n276), .A2(new_n277), .B1(new_n219), .B2(new_n275), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT28), .ZN(new_n312));
  OAI211_X1 g126(.A(KEYINPUT29), .B(new_n287), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT74), .B1(new_n313), .B2(new_n297), .ZN(new_n314));
  INV_X1    g128(.A(G902), .ZN(new_n315));
  OAI22_X1  g129(.A1(new_n270), .A2(new_n271), .B1(new_n268), .B2(new_n269), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n286), .B1(new_n316), .B2(KEYINPUT28), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT74), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT29), .A4(new_n195), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n310), .A2(new_n314), .A3(new_n315), .A4(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G472), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n306), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(G214), .B1(G237), .B2(G902), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT5), .B1(new_n214), .B2(new_n215), .ZN(new_n325));
  NOR3_X1   g139(.A1(new_n202), .A2(KEYINPUT5), .A3(G119), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(G113), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT86), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n325), .A2(KEYINPUT86), .A3(G113), .A4(new_n327), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT82), .B(G104), .ZN(new_n332));
  INV_X1    g146(.A(G107), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT3), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n332), .A2(new_n333), .ZN(new_n336));
  INV_X1    g150(.A(G101), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT3), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(new_n333), .A3(G104), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n335), .A2(new_n336), .A3(new_n337), .A4(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n334), .B1(G104), .B2(new_n333), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G101), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n330), .A2(new_n331), .A3(new_n216), .A4(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT87), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n335), .A2(new_n336), .A3(new_n339), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n347), .A3(G101), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(G101), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(KEYINPUT4), .A3(new_n340), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n219), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n210), .B1(new_n328), .B2(new_n329), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT87), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n352), .A2(new_n353), .A3(new_n343), .A4(new_n331), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n345), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  XOR2_X1   g169(.A(G110), .B(G122), .Z(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n356), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n345), .A2(new_n358), .A3(new_n351), .A4(new_n354), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n357), .A2(KEYINPUT6), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G125), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT77), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT77), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G125), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n249), .A2(new_n365), .ZN(new_n366));
  XOR2_X1   g180(.A(new_n366), .B(KEYINPUT88), .Z(new_n367));
  OR2_X1    g181(.A1(new_n258), .A2(new_n365), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G224), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(G953), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n369), .B(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT6), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n355), .A2(new_n373), .A3(new_n356), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n360), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n367), .A2(KEYINPUT89), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n368), .B1(new_n367), .B2(KEYINPUT89), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT7), .ZN(new_n378));
  OAI22_X1  g192(.A1(new_n376), .A2(new_n377), .B1(new_n378), .B2(new_n371), .ZN(new_n379));
  OR3_X1    g193(.A1(new_n369), .A2(new_n378), .A3(new_n371), .ZN(new_n380));
  INV_X1    g194(.A(new_n328), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n343), .B1(new_n381), .B2(new_n210), .ZN(new_n382));
  XOR2_X1   g196(.A(new_n356), .B(KEYINPUT8), .Z(new_n383));
  NAND2_X1  g197(.A1(new_n352), .A2(new_n331), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n382), .B(new_n383), .C1(new_n384), .C2(new_n343), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n379), .A2(new_n380), .A3(new_n359), .A4(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n375), .A2(new_n315), .A3(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(G210), .B1(G237), .B2(G902), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n375), .A2(new_n315), .A3(new_n388), .A4(new_n386), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n324), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G221), .ZN(new_n393));
  XOR2_X1   g207(.A(KEYINPUT9), .B(G234), .Z(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n394), .B2(new_n315), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n350), .A2(new_n258), .A3(new_n348), .ZN(new_n396));
  INV_X1    g210(.A(new_n254), .ZN(new_n397));
  MUX2_X1   g211(.A(new_n228), .B(new_n232), .S(new_n230), .Z(new_n398));
  NAND3_X1  g212(.A1(new_n340), .A2(new_n342), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT10), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n343), .A2(KEYINPUT10), .A3(new_n234), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n396), .A2(new_n397), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n397), .A2(KEYINPUT83), .ZN(new_n404));
  INV_X1    g218(.A(new_n399), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n234), .B1(new_n340), .B2(new_n342), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT12), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT12), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n409), .B(new_n404), .C1(new_n405), .C2(new_n406), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n403), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(G110), .B(G140), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n191), .A2(G227), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT84), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n396), .A2(new_n401), .A3(new_n402), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n254), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n403), .A3(new_n414), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n416), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n417), .B1(new_n416), .B2(new_n420), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n315), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G469), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n411), .A2(new_n415), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n414), .B1(new_n419), .B2(new_n403), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT85), .ZN(new_n428));
  INV_X1    g242(.A(G469), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n428), .A2(new_n429), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n427), .A2(new_n315), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n395), .B1(new_n424), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n191), .A2(G952), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(G234), .B2(G237), .ZN(new_n436));
  XOR2_X1   g250(.A(KEYINPUT21), .B(G898), .Z(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(KEYINPUT96), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AOI211_X1 g253(.A(new_n315), .B(new_n191), .C1(G234), .C2(G237), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n436), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n392), .A2(new_n434), .A3(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT24), .B(G110), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n444), .B(KEYINPUT75), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n198), .A2(G128), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n231), .A2(G119), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(KEYINPUT23), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT23), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n231), .A3(G119), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n450), .A2(new_n452), .B1(new_n198), .B2(G128), .ZN(new_n453));
  INV_X1    g267(.A(G110), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n449), .A2(new_n455), .ZN(new_n456));
  NOR3_X1   g270(.A1(new_n365), .A2(KEYINPUT16), .A3(G140), .ZN(new_n457));
  NOR2_X1   g271(.A1(G125), .A2(G140), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G140), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n459), .B1(new_n365), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n457), .B1(new_n461), .B2(KEYINPUT16), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G146), .ZN(new_n463));
  XNOR2_X1  g277(.A(G125), .B(G140), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n224), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n456), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT78), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n466), .B(new_n467), .ZN(new_n468));
  OR2_X1    g282(.A1(new_n462), .A2(G146), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n463), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n453), .A2(new_n454), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(KEYINPUT76), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n470), .B(new_n472), .C1(new_n448), .C2(new_n445), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(KEYINPUT22), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(G137), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n468), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n476), .B1(new_n468), .B2(new_n473), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT80), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT80), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n478), .B2(new_n479), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G234), .ZN(new_n485));
  AOI21_X1  g299(.A(G902), .B1(new_n485), .B2(G217), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT81), .ZN(new_n487));
  OAI21_X1  g301(.A(G217), .B1(new_n485), .B2(G902), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n468), .A2(new_n473), .ZN(new_n489));
  INV_X1    g303(.A(new_n476), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(new_n315), .A3(new_n477), .ZN(new_n492));
  AND2_X1   g306(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n488), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n480), .A2(new_n315), .A3(new_n496), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n484), .A2(new_n487), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G122), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n200), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n202), .A2(G122), .ZN(new_n501));
  OAI21_X1  g315(.A(G107), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n206), .A2(G122), .ZN(new_n503));
  INV_X1    g317(.A(new_n501), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n333), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n221), .A2(G128), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n231), .A2(G143), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(G134), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT13), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n231), .B2(G143), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT93), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n507), .A2(KEYINPUT93), .A3(new_n511), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n221), .A2(KEYINPUT13), .A3(G128), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n514), .A2(new_n515), .A3(new_n508), .A4(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n510), .B1(new_n517), .B2(G134), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n506), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT94), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT94), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n506), .A2(new_n521), .A3(new_n518), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT14), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n503), .A2(new_n524), .A3(new_n504), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n525), .B(G107), .C1(new_n524), .C2(new_n503), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n509), .B(G134), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n526), .A2(new_n505), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n523), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n394), .A2(G217), .A3(new_n191), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n528), .B1(new_n520), .B2(new_n522), .ZN(new_n533));
  INV_X1    g347(.A(new_n531), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(G902), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT95), .ZN(new_n537));
  INV_X1    g351(.A(G478), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(KEYINPUT15), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n537), .B(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT90), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n461), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g356(.A(KEYINPUT90), .B(new_n459), .C1(new_n365), .C2(new_n460), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n543), .A3(G146), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(KEYINPUT91), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n190), .A2(new_n191), .A3(G214), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(new_n221), .ZN(new_n547));
  AND2_X1   g361(.A1(KEYINPUT18), .A2(G131), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n544), .A2(KEYINPUT91), .A3(new_n465), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  XOR2_X1   g366(.A(G113), .B(G122), .Z(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(G104), .ZN(new_n554));
  OR2_X1    g368(.A1(new_n547), .A2(G131), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n547), .A2(G131), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n547), .A2(KEYINPUT17), .A3(G131), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n469), .A2(new_n463), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n552), .A2(new_n554), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT19), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT92), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT19), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n464), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT92), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n542), .A2(new_n543), .A3(new_n566), .A4(KEYINPUT19), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n563), .A2(new_n224), .A3(new_n565), .A4(new_n567), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n557), .A2(new_n555), .B1(new_n462), .B2(G146), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n568), .A2(new_n569), .B1(new_n550), .B2(new_n551), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n561), .B1(new_n570), .B2(new_n554), .ZN(new_n571));
  INV_X1    g385(.A(G475), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n572), .A3(new_n315), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT20), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n561), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n554), .B1(new_n552), .B2(new_n560), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n315), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G475), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n571), .A2(KEYINPUT20), .A3(new_n572), .A4(new_n315), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n575), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n540), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n322), .A2(new_n443), .A3(new_n498), .A4(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(G101), .ZN(G3));
  INV_X1    g398(.A(new_n498), .ZN(new_n585));
  INV_X1    g399(.A(new_n303), .ZN(new_n586));
  INV_X1    g400(.A(G472), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n587), .B1(new_n300), .B2(new_n315), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n443), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n575), .A2(new_n579), .A3(new_n580), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n532), .A2(new_n535), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT97), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n593), .B1(new_n533), .B2(new_n534), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n592), .A2(KEYINPUT33), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT33), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n532), .B(new_n535), .C1(new_n593), .C2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n595), .A2(G478), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n536), .A2(new_n538), .ZN(new_n599));
  NAND2_X1  g413(.A1(G478), .A2(G902), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT98), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n591), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT98), .B1(new_n604), .B2(new_n581), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n590), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT34), .B(G104), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(KEYINPUT99), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n608), .B(new_n610), .ZN(G6));
  NAND2_X1  g425(.A1(new_n591), .A2(new_n540), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n590), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT35), .B(G107), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G9));
  NOR2_X1   g429(.A1(new_n586), .A2(new_n588), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n494), .A2(new_n497), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n490), .A2(KEYINPUT36), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n489), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n487), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n443), .A2(new_n582), .A3(new_n616), .A4(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT37), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(new_n454), .ZN(G12));
  INV_X1    g438(.A(new_n621), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n306), .B2(new_n321), .ZN(new_n626));
  INV_X1    g440(.A(G900), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n436), .B1(new_n440), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n612), .A2(new_n628), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n392), .A2(new_n434), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G128), .ZN(G30));
  AOI22_X1  g446(.A1(new_n273), .A2(new_n280), .B1(new_n297), .B2(new_n316), .ZN(new_n633));
  OAI21_X1  g447(.A(G472), .B1(new_n633), .B2(G902), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n306), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT100), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n628), .B(KEYINPUT39), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n434), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n636), .B1(KEYINPUT40), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(KEYINPUT40), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n540), .A2(new_n581), .ZN(new_n642));
  NOR4_X1   g456(.A1(new_n641), .A2(new_n324), .A3(new_n621), .A4(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n390), .A2(new_n391), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT38), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n640), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT101), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(new_n221), .ZN(G45));
  NOR3_X1   g462(.A1(new_n591), .A2(new_n601), .A3(new_n628), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n392), .A2(new_n434), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n322), .A2(new_n650), .A3(new_n621), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT102), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G146), .ZN(G48));
  AND3_X1   g467(.A1(new_n606), .A2(new_n392), .A3(new_n442), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n315), .B1(new_n425), .B2(new_n426), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(G469), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n433), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n395), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n654), .A2(new_n322), .A3(new_n498), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT41), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G113), .ZN(G15));
  INV_X1    g475(.A(new_n612), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n392), .A2(new_n442), .A3(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n322), .A2(new_n663), .A3(new_n498), .A4(new_n658), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G116), .ZN(G18));
  NAND2_X1  g479(.A1(new_n392), .A2(new_n658), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n626), .A2(new_n582), .A3(new_n442), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G119), .ZN(G21));
  OAI21_X1  g483(.A(G472), .B1(new_n290), .B2(G902), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n295), .B(new_n299), .C1(new_n195), .C2(new_n317), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n291), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n585), .A2(new_n673), .A3(new_n441), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n674), .A2(new_n667), .A3(new_n540), .A4(new_n581), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT103), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G122), .ZN(G24));
  NAND4_X1  g491(.A1(new_n649), .A2(new_n670), .A3(new_n621), .A4(new_n672), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n666), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(new_n361), .ZN(G27));
  NAND3_X1  g494(.A1(new_n321), .A2(new_n293), .A3(new_n301), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(KEYINPUT42), .A3(new_n498), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n416), .A2(KEYINPUT104), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n411), .A2(new_n684), .A3(new_n415), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n683), .A2(new_n420), .A3(new_n685), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n686), .A2(new_n315), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n433), .B1(new_n687), .B2(new_n429), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n395), .A2(new_n324), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n688), .A2(new_n390), .A3(new_n391), .A4(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n649), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n682), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n690), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n322), .A2(new_n498), .A3(new_n649), .A4(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT42), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n692), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n240), .ZN(G33));
  NAND4_X1  g511(.A1(new_n322), .A2(new_n498), .A3(new_n629), .A4(new_n693), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G134), .ZN(G36));
  INV_X1    g513(.A(KEYINPUT45), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n700), .B1(new_n421), .B2(new_n422), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n701), .B(G469), .C1(new_n700), .C2(new_n686), .ZN(new_n702));
  XOR2_X1   g516(.A(new_n702), .B(KEYINPUT105), .Z(new_n703));
  NAND2_X1  g517(.A1(G469), .A2(G902), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n703), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n705), .A2(new_n706), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n708), .A2(new_n710), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n433), .A3(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n395), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(new_n714), .A3(new_n638), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n601), .A2(new_n581), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT43), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n718), .B(new_n621), .C1(new_n586), .C2(new_n588), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n715), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n644), .A2(new_n324), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n720), .B(new_n721), .C1(new_n716), .C2(new_n719), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G137), .ZN(G39));
  NAND2_X1  g537(.A1(new_n713), .A2(new_n714), .ZN(new_n724));
  AND2_X1   g538(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n727), .B1(new_n713), .B2(new_n714), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n726), .B1(new_n728), .B2(new_n725), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n721), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n322), .A2(new_n731), .A3(new_n691), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n730), .A2(new_n585), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G140), .ZN(G42));
  NAND2_X1  g548(.A1(new_n498), .A2(new_n689), .ZN(new_n735));
  XOR2_X1   g549(.A(new_n735), .B(KEYINPUT108), .Z(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n717), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n645), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n737), .A2(new_n738), .ZN(new_n741));
  XOR2_X1   g555(.A(new_n657), .B(KEYINPUT49), .Z(new_n742));
  NAND4_X1  g556(.A1(new_n740), .A2(new_n636), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n324), .B(new_n642), .C1(new_n390), .C2(new_n391), .ZN(new_n744));
  INV_X1    g558(.A(new_n628), .ZN(new_n745));
  AND4_X1   g559(.A1(new_n714), .A2(new_n625), .A3(new_n688), .A4(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n635), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n679), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n631), .A2(new_n651), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n679), .B1(new_n626), .B2(new_n630), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(KEYINPUT52), .A3(new_n651), .A4(new_n747), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n690), .A2(new_n691), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n673), .A2(new_n625), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n698), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n756), .B1(new_n755), .B2(new_n757), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n696), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n668), .A2(new_n659), .A3(new_n664), .A4(new_n675), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n612), .B1(new_n591), .B2(new_n601), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n583), .B(new_n622), .C1(new_n590), .C2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n582), .A2(new_n745), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT110), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n626), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n767), .A2(KEYINPUT110), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n771), .A2(new_n434), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n769), .A2(new_n770), .A3(new_n721), .A4(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n772), .A2(new_n626), .A3(new_n721), .A4(new_n768), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT111), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n754), .A2(new_n761), .A3(new_n766), .A4(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n766), .A2(new_n761), .A3(new_n776), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n753), .A2(KEYINPUT114), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n751), .A2(KEYINPUT113), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n753), .A2(KEYINPUT114), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n783), .B1(new_n782), .B2(new_n784), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n781), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n779), .B1(new_n788), .B2(new_n778), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n790));
  OR3_X1    g604(.A1(new_n789), .A2(KEYINPUT115), .A3(new_n790), .ZN(new_n791));
  OAI211_X1 g605(.A(KEYINPUT53), .B(new_n781), .C1(new_n786), .C2(new_n787), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n793), .B1(new_n777), .B2(new_n778), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n777), .A2(new_n793), .A3(new_n778), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n792), .B(new_n790), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT115), .B1(new_n789), .B2(new_n790), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n791), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n718), .A2(new_n436), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n800), .A2(new_n585), .A3(new_n673), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n657), .A2(new_n714), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n721), .B(new_n801), .C1(new_n730), .C2(new_n802), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n644), .A2(new_n395), .A3(new_n324), .ZN(new_n804));
  INV_X1    g618(.A(new_n657), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n800), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n757), .ZN(new_n808));
  INV_X1    g622(.A(new_n806), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n636), .A2(new_n498), .A3(new_n436), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n591), .A2(new_n601), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n801), .A2(new_n658), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n812), .A2(new_n323), .A3(new_n645), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  OR2_X1    g628(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n815));
  OAI221_X1 g629(.A(new_n808), .B1(new_n810), .B2(new_n811), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n814), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n803), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(KEYINPUT51), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(KEYINPUT51), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n822), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n435), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n799), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n810), .A2(new_n607), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n681), .A2(new_n498), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n807), .A2(new_n829), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n830), .B(KEYINPUT48), .Z(new_n831));
  AND2_X1   g645(.A1(new_n801), .A2(new_n667), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n827), .A2(new_n828), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(G952), .A2(G953), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n743), .B1(new_n833), .B2(new_n834), .ZN(G75));
  OAI21_X1  g649(.A(new_n792), .B1(new_n794), .B2(new_n795), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(G902), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(G210), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT56), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n360), .A2(new_n374), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(new_n372), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT55), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n839), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n843), .B1(new_n839), .B2(new_n840), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n191), .A2(G952), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(G51));
  INV_X1    g661(.A(KEYINPUT121), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n795), .A2(new_n794), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n751), .A2(KEYINPUT113), .ZN(new_n850));
  INV_X1    g664(.A(new_n784), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n753), .A2(KEYINPUT114), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI211_X1 g667(.A(new_n778), .B(new_n780), .C1(new_n853), .C2(new_n785), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT54), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n855), .A2(new_n856), .A3(new_n796), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n836), .A2(KEYINPUT119), .A3(KEYINPUT54), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n704), .B(KEYINPUT57), .Z(new_n859));
  NAND3_X1  g673(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT120), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n857), .A2(new_n862), .A3(new_n858), .A4(new_n859), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n848), .B1(new_n864), .B2(new_n427), .ZN(new_n865));
  INV_X1    g679(.A(new_n427), .ZN(new_n866));
  AOI211_X1 g680(.A(KEYINPUT121), .B(new_n866), .C1(new_n861), .C2(new_n863), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n837), .A2(new_n703), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n846), .B1(new_n868), .B2(new_n869), .ZN(G54));
  NAND3_X1  g684(.A1(new_n838), .A2(KEYINPUT58), .A3(G475), .ZN(new_n871));
  INV_X1    g685(.A(new_n571), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n871), .A2(new_n872), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n873), .A2(new_n874), .A3(new_n846), .ZN(G60));
  NAND2_X1  g689(.A1(new_n595), .A2(new_n597), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n600), .B(KEYINPUT59), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n876), .B1(new_n798), .B2(new_n877), .ZN(new_n878));
  AND4_X1   g692(.A1(new_n876), .A2(new_n857), .A3(new_n858), .A4(new_n877), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n878), .A2(new_n846), .A3(new_n879), .ZN(G63));
  NAND2_X1  g694(.A1(G217), .A2(G902), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT122), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT60), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n836), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n884), .A2(new_n484), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n619), .B(KEYINPUT123), .Z(new_n886));
  AOI211_X1 g700(.A(new_n846), .B(new_n885), .C1(new_n884), .C2(new_n886), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT61), .ZN(G66));
  NOR2_X1   g702(.A1(new_n766), .A2(G953), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT124), .ZN(new_n890));
  OAI21_X1  g704(.A(G953), .B1(new_n439), .B2(new_n370), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n841), .B1(G898), .B2(new_n191), .ZN(new_n893));
  XNOR2_X1  g707(.A(KEYINPUT125), .B(KEYINPUT126), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n893), .B(new_n894), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n892), .B(new_n895), .ZN(G69));
  AND2_X1   g710(.A1(new_n733), .A2(new_n722), .ZN(new_n897));
  INV_X1    g711(.A(new_n715), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n898), .A2(new_n829), .A3(new_n744), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n752), .A2(new_n651), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n696), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n897), .A2(new_n698), .A3(new_n899), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n191), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n262), .A2(new_n266), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n563), .A2(new_n565), .A3(new_n567), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n904), .B(new_n905), .Z(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n903), .B(new_n907), .C1(G227), .C2(new_n191), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n646), .A2(new_n651), .A3(new_n752), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT62), .Z(new_n910));
  NOR2_X1   g724(.A1(new_n731), .A2(new_n639), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n911), .A2(new_n498), .A3(new_n322), .A4(new_n763), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n897), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  OR3_X1    g727(.A1(new_n913), .A2(G953), .A3(new_n907), .ZN(new_n914));
  OAI21_X1  g728(.A(G900), .B1(new_n907), .B2(G227), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(G953), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n908), .A2(new_n914), .A3(new_n916), .ZN(G72));
  NAND2_X1  g731(.A1(new_n913), .A2(new_n766), .ZN(new_n918));
  NAND2_X1  g732(.A1(G472), .A2(G902), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT63), .Z(new_n920));
  NAND2_X1  g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT127), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n918), .A2(KEYINPUT127), .A3(new_n920), .ZN(new_n924));
  AND4_X1   g738(.A1(new_n195), .A2(new_n923), .A3(new_n307), .A4(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n789), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n294), .A2(new_n308), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n926), .A2(new_n920), .A3(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n766), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n920), .B1(new_n902), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n297), .ZN(new_n931));
  OAI221_X1 g745(.A(new_n928), .B1(G952), .B2(new_n191), .C1(new_n931), .C2(new_n307), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n925), .A2(new_n932), .ZN(G57));
endmodule


