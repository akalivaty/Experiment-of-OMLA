//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 0 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G116), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT2), .A2(G113), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT71), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT71), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT2), .A3(G113), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(KEYINPUT2), .A2(G113), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n192), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n200));
  INV_X1    g014(.A(G113), .ZN(new_n201));
  AOI22_X1  g015(.A1(new_n194), .A2(new_n196), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n192), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AND2_X1   g018(.A1(new_n199), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT65), .A2(G146), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT65), .A2(G146), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(KEYINPUT64), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n215), .B1(KEYINPUT0), .B2(G128), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n214), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n212), .A2(new_n217), .A3(KEYINPUT66), .ZN(new_n218));
  OR2_X1    g032(.A1(KEYINPUT65), .A2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(KEYINPUT65), .A2(G146), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(G143), .A3(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n210), .A2(G143), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n221), .A2(KEYINPUT0), .A3(G128), .A4(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n218), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT66), .B1(new_n212), .B2(new_n217), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT67), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G137), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G134), .ZN(new_n229));
  NOR2_X1   g043(.A1(KEYINPUT68), .A2(KEYINPUT11), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT68), .A2(KEYINPUT11), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n229), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G134), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n232), .B1(new_n234), .B2(G137), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(G137), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(G131), .B1(new_n233), .B2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n234), .A2(G137), .ZN(new_n239));
  INV_X1    g053(.A(new_n232), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(new_n230), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT69), .B(G131), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n241), .A2(new_n236), .A3(new_n235), .A4(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n245));
  INV_X1    g059(.A(new_n211), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT65), .B(G146), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n246), .B1(new_n247), .B2(new_n206), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n216), .A2(new_n213), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n215), .A2(KEYINPUT0), .A3(G128), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n245), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n252), .A2(new_n218), .A3(new_n253), .A4(new_n224), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n227), .A2(new_n244), .A3(new_n254), .ZN(new_n255));
  NOR3_X1   g069(.A1(new_n207), .A2(new_n208), .A3(new_n206), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n257));
  OAI21_X1  g071(.A(G128), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n207), .A2(new_n208), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n222), .B1(new_n259), .B2(G143), .ZN(new_n260));
  INV_X1    g074(.A(G128), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(KEYINPUT1), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n258), .A2(new_n212), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n229), .A2(new_n236), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G131), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n264), .B1(new_n243), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n243), .A2(new_n266), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n264), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n205), .B1(new_n255), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n199), .A2(new_n204), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n221), .A2(new_n223), .A3(new_n262), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n261), .B1(new_n221), .B2(KEYINPUT1), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n274), .B1(new_n275), .B2(new_n248), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n273), .B1(new_n269), .B2(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n244), .A2(new_n252), .A3(new_n224), .A4(new_n218), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT28), .B1(new_n272), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT28), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(G237), .A2(G953), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G210), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n286), .B(KEYINPUT27), .ZN(new_n287));
  XNOR2_X1  g101(.A(KEYINPUT26), .B(G101), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n287), .B(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n187), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  AOI211_X1 g105(.A(KEYINPUT72), .B(new_n289), .C1(new_n281), .C2(new_n283), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT30), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n255), .A2(new_n293), .A3(new_n271), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n269), .A2(new_n276), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n293), .B1(new_n278), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n280), .B1(new_n298), .B2(new_n273), .ZN(new_n299));
  AOI21_X1  g113(.A(KEYINPUT31), .B1(new_n299), .B2(new_n289), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n205), .B1(new_n294), .B2(new_n297), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT31), .ZN(new_n302));
  NOR4_X1   g116(.A1(new_n301), .A2(new_n302), .A3(new_n280), .A4(new_n290), .ZN(new_n303));
  OAI22_X1  g117(.A1(new_n291), .A2(new_n292), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(G472), .A2(G902), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT32), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n283), .A2(KEYINPUT29), .A3(new_n289), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n252), .A2(new_n224), .A3(new_n218), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n238), .A2(new_n243), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n243), .A2(new_n266), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n205), .B1(new_n263), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT73), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n277), .A2(new_n278), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n278), .A2(new_n295), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n273), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n205), .B1(new_n278), .B2(new_n295), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT74), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n319), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n310), .B1(new_n326), .B2(KEYINPUT28), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT75), .B1(new_n327), .B2(G902), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n329));
  INV_X1    g143(.A(G902), .ZN(new_n330));
  AOI22_X1  g144(.A1(new_n316), .A2(new_n318), .B1(KEYINPUT74), .B2(new_n324), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n282), .B1(new_n331), .B2(new_n323), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n329), .B(new_n330), .C1(new_n332), .C2(new_n310), .ZN(new_n333));
  INV_X1    g147(.A(new_n283), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(new_n290), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT29), .B1(new_n281), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n290), .B1(new_n301), .B2(new_n280), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n328), .A2(new_n333), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G472), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n312), .B1(new_n311), .B2(KEYINPUT67), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n341), .A2(new_n254), .B1(new_n270), .B2(new_n268), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n279), .B1(new_n342), .B2(new_n205), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n334), .B1(new_n343), .B2(KEYINPUT28), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT72), .B1(new_n344), .B2(new_n289), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n284), .A2(new_n187), .A3(new_n290), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n296), .B1(new_n342), .B2(new_n293), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n279), .B(new_n289), .C1(new_n348), .C2(new_n205), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n302), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n299), .A2(KEYINPUT31), .A3(new_n289), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n306), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n309), .B(new_n340), .C1(new_n353), .C2(KEYINPUT32), .ZN(new_n354));
  INV_X1    g168(.A(G953), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(G221), .A3(G234), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(KEYINPUT79), .ZN(new_n357));
  XNOR2_X1  g171(.A(KEYINPUT22), .B(G137), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n357), .B(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT77), .ZN(new_n361));
  INV_X1    g175(.A(G140), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G125), .ZN(new_n363));
  INV_X1    g177(.A(G125), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G140), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT76), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n364), .A2(KEYINPUT76), .A3(G140), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(KEYINPUT16), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT16), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n363), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n361), .B1(new_n372), .B2(G146), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT23), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n374), .B1(new_n188), .B2(G128), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n261), .A2(KEYINPUT23), .A3(G119), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n375), .B(new_n376), .C1(G119), .C2(new_n261), .ZN(new_n377));
  XNOR2_X1  g191(.A(G119), .B(G128), .ZN(new_n378));
  XOR2_X1   g192(.A(KEYINPUT24), .B(G110), .Z(new_n379));
  OAI22_X1  g193(.A1(new_n377), .A2(G110), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(G125), .B(G140), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n259), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n382), .A2(KEYINPUT78), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT78), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n384), .B1(new_n259), .B2(new_n381), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n380), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  AOI211_X1 g200(.A(KEYINPUT77), .B(new_n210), .C1(new_n369), .C2(new_n371), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n373), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n377), .A2(G110), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n379), .A2(new_n378), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n372), .A2(G146), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n369), .A2(new_n210), .A3(new_n371), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n360), .B1(new_n388), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n392), .A2(KEYINPUT77), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n372), .A2(new_n361), .A3(G146), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n382), .B(KEYINPUT78), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n396), .A2(new_n397), .A3(new_n398), .A4(new_n380), .ZN(new_n399));
  INV_X1    g213(.A(new_n394), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n400), .A3(new_n359), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n395), .A2(new_n401), .A3(new_n330), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT25), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(KEYINPUT80), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(KEYINPUT80), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n395), .A2(new_n401), .A3(new_n330), .A4(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G217), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n408), .B1(G234), .B2(new_n330), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n409), .A2(G902), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT81), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n395), .A2(new_n401), .A3(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(KEYINPUT82), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G475), .ZN(new_n416));
  INV_X1    g230(.A(G237), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(new_n355), .A3(G214), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n206), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n285), .A2(G143), .A3(G214), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT18), .ZN(new_n421));
  INV_X1    g235(.A(G131), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n419), .B(new_n420), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n420), .ZN(new_n424));
  AOI21_X1  g238(.A(G143), .B1(new_n285), .B2(G214), .ZN(new_n425));
  OAI211_X1 g239(.A(KEYINPUT18), .B(G131), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n383), .A2(new_n385), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n367), .A2(new_n368), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n428), .A2(new_n210), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n423), .B(new_n426), .C1(new_n427), .C2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n242), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n424), .B2(new_n425), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT17), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n419), .A2(new_n242), .A3(new_n420), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(KEYINPUT17), .B(new_n431), .C1(new_n424), .C2(new_n425), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n392), .A2(new_n435), .A3(new_n393), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n430), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G113), .B(G122), .ZN(new_n439));
  INV_X1    g253(.A(G104), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n439), .B(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n430), .A2(new_n437), .A3(new_n441), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n416), .B1(new_n445), .B2(new_n330), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n426), .A2(new_n423), .ZN(new_n448));
  INV_X1    g262(.A(new_n429), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n448), .B1(new_n398), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n373), .A2(new_n387), .ZN(new_n451));
  OR2_X1    g265(.A1(new_n381), .A2(KEYINPUT19), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n364), .A2(KEYINPUT76), .A3(G140), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n381), .B2(new_n366), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT19), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n456), .A2(new_n259), .B1(new_n432), .B2(new_n434), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n450), .B1(new_n451), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n444), .B1(new_n458), .B2(new_n441), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT91), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT20), .ZN(new_n461));
  NOR2_X1   g275(.A1(G475), .A2(G902), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n459), .A2(new_n460), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n457), .A2(new_n396), .A3(new_n397), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n441), .B1(new_n465), .B2(new_n430), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n430), .A2(new_n441), .A3(new_n437), .ZN(new_n467));
  OAI21_X1  g281(.A(KEYINPUT91), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI22_X1  g282(.A1(new_n468), .A2(new_n461), .B1(new_n459), .B2(new_n462), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n447), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT92), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n432), .A2(new_n434), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n381), .A2(KEYINPUT19), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(new_n428), .B2(KEYINPUT19), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n474), .B1(new_n476), .B2(new_n247), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n477), .A2(new_n373), .A3(new_n387), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n442), .B1(new_n478), .B2(new_n450), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n460), .B1(new_n479), .B2(new_n444), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n473), .B1(new_n480), .B2(KEYINPUT20), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n463), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(KEYINPUT92), .A3(new_n447), .ZN(new_n483));
  NAND2_X1  g297(.A1(G234), .A2(G237), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(G952), .A3(new_n355), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n485), .B(KEYINPUT95), .Z(new_n486));
  XNOR2_X1  g300(.A(KEYINPUT21), .B(G898), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n487), .A2(G902), .A3(G953), .A4(new_n484), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G478), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(KEYINPUT15), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(G128), .B(G143), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n261), .A2(G143), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT13), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n234), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n493), .B(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G122), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G116), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n190), .A2(G122), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT93), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G116), .B(G122), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(KEYINPUT93), .ZN(new_n505));
  INV_X1    g319(.A(G107), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n501), .A2(new_n502), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n504), .A2(KEYINPUT93), .ZN(new_n509));
  AOI21_X1  g323(.A(G107), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n497), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n506), .B1(new_n503), .B2(new_n505), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n190), .A2(KEYINPUT14), .A3(G122), .ZN(new_n513));
  OAI211_X1 g327(.A(G107), .B(new_n513), .C1(new_n501), .C2(KEYINPUT14), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n493), .B(new_n234), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n512), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT9), .B(G234), .ZN(new_n518));
  NOR3_X1   g332(.A1(new_n518), .A2(new_n408), .A3(G953), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n511), .A2(new_n516), .A3(new_n519), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n492), .B1(new_n523), .B2(new_n330), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  AOI211_X1 g339(.A(G902), .B(new_n491), .C1(new_n521), .C2(new_n522), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n527), .A3(KEYINPUT94), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT94), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n529), .B1(new_n524), .B2(new_n526), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n489), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n472), .A2(new_n483), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G469), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT3), .B1(new_n440), .B2(G107), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT3), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(new_n506), .A3(G104), .ZN(new_n536));
  INV_X1    g350(.A(G101), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n440), .A2(G107), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n534), .A2(new_n536), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n440), .A2(G107), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n506), .A2(G104), .ZN(new_n541));
  OAI21_X1  g355(.A(G101), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT1), .B1(new_n206), .B2(G146), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n221), .A2(new_n223), .B1(G128), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n274), .B1(new_n546), .B2(KEYINPUT83), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT83), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n261), .B1(new_n211), .B2(KEYINPUT1), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n260), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n544), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n263), .A2(new_n543), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n312), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  XOR2_X1   g367(.A(KEYINPUT86), .B(KEYINPUT12), .Z(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(KEYINPUT86), .A2(KEYINPUT12), .ZN(new_n556));
  AOI211_X1 g370(.A(new_n312), .B(new_n556), .C1(new_n551), .C2(new_n552), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT10), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n551), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n218), .A2(new_n224), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n534), .A2(new_n536), .A3(new_n538), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT4), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n563), .A3(G101), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(G101), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(KEYINPUT4), .A3(new_n539), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n561), .A2(new_n252), .A3(new_n564), .A4(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT84), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n539), .B2(new_n542), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n539), .A2(new_n542), .A3(new_n568), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n276), .B(KEYINPUT10), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n238), .A2(KEYINPUT85), .A3(new_n243), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT85), .B1(new_n238), .B2(new_n243), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n560), .A2(new_n567), .A3(new_n571), .A4(new_n574), .ZN(new_n575));
  XOR2_X1   g389(.A(G110), .B(G140), .Z(new_n576));
  NAND2_X1  g390(.A1(new_n355), .A2(G227), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n558), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n560), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n566), .A2(new_n564), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n571), .B1(new_n311), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n244), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n579), .B1(new_n585), .B2(new_n575), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n533), .B(new_n330), .C1(new_n581), .C2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n579), .A3(new_n575), .ZN(new_n588));
  OR2_X1    g402(.A1(new_n553), .A2(new_n554), .ZN(new_n589));
  INV_X1    g403(.A(new_n557), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n582), .A2(new_n584), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n589), .A2(new_n590), .B1(new_n591), .B2(new_n574), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n588), .B(G469), .C1(new_n592), .C2(new_n579), .ZN(new_n593));
  NAND2_X1  g407(.A1(G469), .A2(G902), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n587), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(G214), .B1(G237), .B2(G902), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(G210), .B1(G237), .B2(G902), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n273), .A2(new_n564), .A3(new_n566), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n190), .A2(G119), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT5), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n201), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT5), .ZN(new_n604));
  AOI22_X1  g418(.A1(new_n202), .A2(new_n203), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n605), .B1(new_n570), .B2(new_n569), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n600), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n498), .A2(G110), .ZN(new_n608));
  INV_X1    g422(.A(G110), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(G122), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT87), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n608), .A2(new_n610), .A3(KEYINPUT87), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n607), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n600), .A2(new_n606), .A3(new_n614), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(KEYINPUT6), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT6), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n607), .A2(new_n619), .A3(new_n615), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n252), .A2(new_n218), .A3(G125), .A4(new_n224), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n276), .A2(new_n364), .ZN(new_n622));
  INV_X1    g436(.A(G224), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(G953), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n621), .A2(new_n622), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n625), .B1(new_n621), .B2(new_n622), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n618), .A2(new_n620), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n621), .A2(new_n622), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(KEYINPUT7), .A3(new_n625), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n625), .A2(KEYINPUT7), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n621), .A2(new_n622), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n631), .A2(new_n617), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT89), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n539), .A2(new_n542), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT88), .B(KEYINPUT8), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n612), .A2(new_n613), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n637), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n608), .A2(new_n610), .A3(KEYINPUT87), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n639), .B1(new_n640), .B2(new_n611), .ZN(new_n641));
  AOI22_X1  g455(.A1(new_n605), .A2(new_n636), .B1(new_n638), .B2(new_n641), .ZN(new_n642));
  OR2_X1    g456(.A1(new_n605), .A2(new_n636), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n642), .A2(KEYINPUT90), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT90), .B1(new_n642), .B2(new_n643), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n330), .B1(new_n634), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n599), .B1(new_n629), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n618), .A2(new_n620), .A3(new_n628), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n617), .A2(new_n633), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n650), .B(new_n631), .C1(new_n645), .C2(new_n644), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n649), .A2(new_n651), .A3(new_n330), .A4(new_n598), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n597), .B1(new_n648), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(G221), .B1(new_n518), .B2(G902), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n595), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n532), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n354), .A2(new_n415), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G101), .ZN(G3));
  INV_X1    g472(.A(G472), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n304), .B2(new_n330), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n595), .A2(new_n654), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n660), .A2(new_n353), .A3(new_n661), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n662), .A2(new_n415), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n472), .A2(new_n483), .ZN(new_n664));
  INV_X1    g478(.A(new_n489), .ZN(new_n665));
  AOI211_X1 g479(.A(G478), .B(G902), .C1(new_n521), .C2(new_n522), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n490), .A2(new_n330), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n523), .B(KEYINPUT33), .Z(new_n668));
  AOI211_X1 g482(.A(new_n666), .B(new_n667), .C1(new_n668), .C2(G478), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n664), .A2(new_n665), .A3(new_n653), .A4(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n663), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT34), .B(G104), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G6));
  AND2_X1   g488(.A1(new_n528), .A2(new_n530), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n473), .A2(KEYINPUT20), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n459), .A2(new_n461), .A3(new_n462), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n446), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n489), .B(KEYINPUT96), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n653), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n663), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT35), .B(G107), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G9));
  NAND2_X1  g499(.A1(new_n304), .A2(new_n330), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n353), .B1(new_n686), .B2(G472), .ZN(new_n687));
  INV_X1    g501(.A(new_n661), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n399), .A2(new_n400), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n689), .A2(KEYINPUT97), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n360), .A2(KEYINPUT36), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n689), .A2(KEYINPUT97), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n691), .B1(new_n690), .B2(new_n692), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n412), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n410), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n653), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n532), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n687), .A2(new_n688), .A3(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT37), .B(G110), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G12));
  INV_X1    g515(.A(new_n697), .ZN(new_n702));
  INV_X1    g516(.A(G900), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n484), .A2(new_n703), .A3(G902), .A4(G953), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT98), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n486), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT99), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n661), .A2(new_n679), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n354), .A2(new_n702), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G128), .ZN(G30));
  XOR2_X1   g524(.A(new_n707), .B(KEYINPUT39), .Z(new_n711));
  NAND2_X1  g525(.A1(new_n688), .A2(new_n711), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n712), .A2(KEYINPUT40), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n648), .A2(new_n652), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n715));
  XOR2_X1   g529(.A(new_n714), .B(new_n715), .Z(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n696), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n712), .A2(KEYINPUT40), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n528), .A2(new_n530), .A3(new_n596), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n664), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n713), .A2(new_n718), .A3(new_n719), .A4(new_n721), .ZN(new_n722));
  AOI22_X1  g536(.A1(new_n345), .A2(new_n346), .B1(new_n350), .B2(new_n351), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n307), .B1(new_n723), .B2(new_n306), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n326), .A2(new_n289), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(G902), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n289), .B1(new_n301), .B2(new_n280), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n659), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n728), .B1(new_n304), .B2(new_n308), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n724), .A2(new_n729), .A3(KEYINPUT101), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT101), .B1(new_n724), .B2(new_n729), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n722), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n206), .ZN(G45));
  INV_X1    g549(.A(new_n707), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT92), .B1(new_n482), .B2(new_n447), .ZN(new_n737));
  AOI211_X1 g551(.A(new_n471), .B(new_n446), .C1(new_n481), .C2(new_n463), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n669), .B(new_n736), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n661), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n354), .A2(new_n740), .A3(new_n702), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G146), .ZN(G48));
  NOR2_X1   g556(.A1(new_n581), .A2(new_n586), .ZN(new_n743));
  OAI21_X1  g557(.A(G469), .B1(new_n743), .B2(G902), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n415), .A2(new_n654), .A3(new_n587), .A4(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n671), .A2(new_n354), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(KEYINPUT41), .B(G113), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G15));
  NAND3_X1  g563(.A1(new_n354), .A2(new_n682), .A3(new_n746), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G116), .ZN(G18));
  NAND3_X1  g565(.A1(new_n744), .A2(new_n654), .A3(new_n587), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n532), .A2(new_n697), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n354), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G119), .ZN(G21));
  OAI211_X1 g569(.A(new_n714), .B(new_n720), .C1(new_n737), .C2(new_n738), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n744), .A2(new_n654), .A3(new_n587), .A4(new_n680), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g572(.A(new_n305), .B(KEYINPUT102), .Z(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT103), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n761), .B1(new_n332), .B2(new_n334), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n317), .B1(new_n277), .B2(new_n278), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n277), .A2(new_n317), .A3(new_n278), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n325), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n324), .A2(KEYINPUT74), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT28), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(KEYINPUT103), .A3(new_n283), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n762), .A2(new_n768), .A3(new_n290), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n760), .B1(new_n769), .B2(new_n352), .ZN(new_n770));
  XOR2_X1   g584(.A(KEYINPUT104), .B(G472), .Z(new_n771));
  AOI21_X1  g585(.A(new_n770), .B1(new_n686), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n410), .A2(new_n414), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT105), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n758), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G122), .ZN(G24));
  INV_X1    g590(.A(new_n739), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n744), .A2(new_n653), .A3(new_n654), .A4(new_n587), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n772), .A2(new_n696), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  XOR2_X1   g594(.A(KEYINPUT106), .B(G125), .Z(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G27));
  AND3_X1   g596(.A1(new_n648), .A2(new_n596), .A3(new_n652), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n595), .A2(new_n783), .A3(new_n654), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n739), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n354), .A2(new_n785), .A3(new_n774), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n739), .A2(KEYINPUT42), .A3(new_n784), .ZN(new_n787));
  AOI22_X1  g601(.A1(new_n304), .A2(new_n308), .B1(new_n339), .B2(G472), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n773), .B1(new_n788), .B2(new_n724), .ZN(new_n789));
  AOI22_X1  g603(.A1(new_n786), .A2(KEYINPUT42), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G131), .ZN(G33));
  INV_X1    g605(.A(new_n783), .ZN(new_n792));
  NOR4_X1   g606(.A1(new_n661), .A2(new_n792), .A3(new_n679), .A4(new_n707), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G134), .ZN(G36));
  INV_X1    g609(.A(KEYINPUT108), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n664), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n472), .A2(KEYINPUT108), .A3(new_n483), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n668), .A2(G478), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n666), .A2(new_n667), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT43), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n797), .A2(new_n798), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n472), .A2(new_n669), .A3(new_n483), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n805), .A2(KEYINPUT107), .A3(new_n802), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT107), .B1(new_n805), .B2(new_n802), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n804), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n696), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n687), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT44), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n783), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT109), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n813), .B(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n588), .B1(new_n592), .B2(new_n579), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT45), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n533), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n818), .B1(new_n817), .B2(new_n816), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n594), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT46), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(KEYINPUT46), .A3(new_n594), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(new_n587), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n654), .A3(new_n711), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n825), .B1(new_n811), .B2(new_n812), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n815), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G137), .ZN(G39));
  NAND2_X1  g642(.A1(new_n824), .A2(new_n654), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT47), .ZN(new_n830));
  INV_X1    g644(.A(new_n354), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n773), .A3(new_n777), .A4(new_n783), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(new_n362), .ZN(G42));
  NAND2_X1  g648(.A1(new_n717), .A2(new_n774), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n744), .A2(new_n587), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(KEYINPUT49), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n836), .A2(KEYINPUT49), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n669), .A2(new_n596), .A3(new_n654), .ZN(new_n839));
  NOR4_X1   g653(.A1(new_n835), .A2(new_n837), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n840), .A2(new_n733), .A3(new_n797), .A4(new_n798), .ZN(new_n841));
  NAND2_X1  g655(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n842));
  INV_X1    g656(.A(new_n808), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(new_n486), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n844), .A2(new_n774), .A3(new_n772), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n597), .B1(KEYINPUT116), .B2(KEYINPUT50), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n716), .A2(new_n752), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n842), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n752), .A2(new_n792), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n773), .A2(new_n486), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n733), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n851), .A2(new_n664), .A3(new_n669), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n836), .A2(new_n654), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n792), .B1(new_n830), .B2(new_n854), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n847), .A2(new_n842), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n845), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n771), .B1(new_n723), .B2(G902), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n769), .A2(new_n352), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n759), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n858), .A2(new_n696), .A3(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n844), .A2(KEYINPUT117), .A3(new_n849), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT117), .B1(new_n844), .B2(new_n849), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n853), .B(new_n857), .C1(new_n861), .C2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n354), .A2(new_n774), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(new_n862), .B2(new_n863), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT48), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n355), .A2(G952), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n669), .B1(new_n737), .B2(new_n738), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n851), .A2(new_n873), .ZN(new_n874));
  AOI211_X1 g688(.A(new_n872), .B(new_n874), .C1(new_n845), .C2(new_n779), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n867), .A2(new_n868), .A3(new_n871), .A4(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT111), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n595), .A2(new_n783), .A3(new_n654), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n801), .B1(new_n472), .B2(new_n483), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n880), .A3(new_n736), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n878), .B1(new_n861), .B2(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n785), .A2(new_n772), .A3(KEYINPUT111), .A4(new_n696), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n789), .A2(new_n656), .B1(new_n662), .B2(new_n698), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n524), .A2(new_n526), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n472), .A2(new_n483), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n681), .B1(new_n873), .B2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n889), .A2(new_n687), .A3(new_n415), .A4(new_n688), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n884), .A2(new_n885), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n678), .A2(new_n886), .A3(new_n736), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n784), .A2(new_n809), .A3(new_n892), .ZN(new_n893));
  AOI22_X1  g707(.A1(new_n789), .A2(new_n793), .B1(new_n354), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n786), .A2(KEYINPUT42), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n789), .A2(new_n787), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n747), .A2(new_n750), .A3(new_n775), .A4(new_n754), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT110), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n745), .B1(new_n788), .B2(new_n724), .ZN(new_n901));
  AOI22_X1  g715(.A1(new_n901), .A2(new_n671), .B1(new_n354), .B2(new_n753), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT110), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n902), .A2(new_n903), .A3(new_n750), .A4(new_n775), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n898), .A2(KEYINPUT112), .A3(new_n900), .A4(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT112), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n900), .A2(new_n904), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n890), .A2(new_n657), .A3(new_n699), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n908), .A2(new_n790), .A3(new_n894), .A4(new_n884), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n906), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n756), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n661), .A2(new_n696), .A3(new_n707), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n912), .B(new_n913), .C1(new_n731), .C2(new_n732), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n354), .B(new_n702), .C1(new_n740), .C2(new_n708), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n914), .A2(KEYINPUT113), .A3(new_n780), .A4(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT113), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n915), .A2(new_n780), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n913), .A2(new_n912), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n724), .A2(new_n729), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT101), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n919), .B1(new_n922), .B2(new_n730), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n917), .B1(new_n918), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n916), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT52), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n916), .A2(new_n924), .A3(KEYINPUT52), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n877), .B1(new_n911), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT54), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n918), .A2(new_n923), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n932), .A2(new_n926), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n925), .B2(new_n926), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n909), .A2(new_n877), .A3(new_n899), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n930), .A2(new_n931), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(KEYINPUT53), .B1(new_n911), .B2(new_n929), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n934), .A2(new_n905), .A3(new_n910), .A4(new_n877), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n938), .A2(KEYINPUT54), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n937), .A2(new_n940), .A3(KEYINPUT114), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT114), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n938), .A2(new_n942), .A3(KEYINPUT54), .A4(new_n939), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT115), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT115), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n941), .A2(new_n946), .A3(new_n943), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n876), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(G952), .A2(G953), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n841), .B1(new_n948), .B2(new_n949), .ZN(G75));
  INV_X1    g764(.A(KEYINPUT56), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n930), .A2(new_n936), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n952), .A2(new_n330), .ZN(new_n953));
  INV_X1    g767(.A(G210), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n618), .A2(new_n620), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(new_n628), .Z(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT55), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n958), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n951), .B(new_n960), .C1(new_n953), .C2(new_n954), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n355), .A2(G952), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n959), .A2(new_n961), .A3(new_n963), .ZN(G51));
  XOR2_X1   g778(.A(new_n594), .B(KEYINPUT57), .Z(new_n965));
  INV_X1    g779(.A(new_n937), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n931), .B1(new_n930), .B2(new_n936), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(KEYINPUT118), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT118), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n970), .B(new_n965), .C1(new_n966), .C2(new_n967), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n743), .B(KEYINPUT119), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n969), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n953), .A2(new_n819), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n962), .B1(new_n973), .B2(new_n974), .ZN(G54));
  NOR2_X1   g789(.A1(new_n952), .A2(new_n330), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n976), .A2(KEYINPUT58), .A3(G475), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n466), .A2(new_n467), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n977), .A2(new_n978), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n979), .A2(new_n980), .A3(new_n962), .ZN(G60));
  NOR2_X1   g795(.A1(new_n966), .A2(new_n967), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n667), .B(KEYINPUT59), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n668), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n963), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n983), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n945), .A2(new_n947), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n985), .B1(new_n987), .B2(new_n668), .ZN(G63));
  NAND2_X1  g802(.A1(G217), .A2(G902), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT60), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n952), .A2(new_n990), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n693), .A2(new_n694), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n395), .A2(new_n401), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n993), .B(new_n963), .C1(new_n994), .C2(new_n991), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT61), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n991), .A2(new_n994), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n998), .A2(KEYINPUT61), .A3(new_n963), .A4(new_n993), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n997), .A2(new_n999), .ZN(G66));
  OAI21_X1  g814(.A(G953), .B1(new_n487), .B2(new_n623), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n900), .A2(new_n904), .A3(new_n908), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1001), .B1(new_n1003), .B2(G953), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n956), .B1(G898), .B2(new_n355), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT120), .Z(new_n1006));
  XNOR2_X1  g820(.A(new_n1004), .B(new_n1006), .ZN(G69));
  AOI21_X1  g821(.A(new_n355), .B1(G227), .B2(G900), .ZN(new_n1008));
  OR2_X1    g822(.A1(new_n734), .A2(new_n918), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1009), .A2(KEYINPUT62), .ZN(new_n1010));
  INV_X1    g824(.A(new_n789), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n873), .A2(new_n888), .ZN(new_n1012));
  NOR4_X1   g826(.A1(new_n1011), .A2(new_n712), .A3(new_n792), .A4(new_n1012), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT121), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1015), .B1(new_n1009), .B2(KEYINPUT62), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1009), .A2(new_n1015), .A3(KEYINPUT62), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1014), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n833), .B1(new_n815), .B2(new_n826), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n355), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n298), .B(new_n456), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1008), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n703), .A2(G953), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1026), .B(KEYINPUT122), .ZN(new_n1027));
  INV_X1    g841(.A(new_n833), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n869), .A2(new_n912), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n794), .B1(new_n1029), .B2(new_n825), .ZN(new_n1030));
  INV_X1    g844(.A(new_n790), .ZN(new_n1031));
  NOR3_X1   g845(.A1(new_n1030), .A2(new_n1031), .A3(new_n918), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n827), .A2(new_n1028), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1027), .B1(new_n1033), .B2(new_n355), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1025), .B1(new_n1024), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1036));
  OAI21_X1  g850(.A(KEYINPUT123), .B1(new_n1034), .B2(new_n1024), .ZN(new_n1037));
  INV_X1    g851(.A(KEYINPUT123), .ZN(new_n1038));
  AOI21_X1  g852(.A(G953), .B1(new_n1020), .B2(new_n1032), .ZN(new_n1039));
  OAI211_X1 g853(.A(new_n1038), .B(new_n1023), .C1(new_n1039), .C2(new_n1027), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n1036), .A2(new_n1037), .A3(new_n1040), .ZN(new_n1041));
  AND3_X1   g855(.A1(new_n1041), .A2(KEYINPUT124), .A3(new_n1008), .ZN(new_n1042));
  AOI21_X1  g856(.A(KEYINPUT124), .B1(new_n1041), .B2(new_n1008), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n1035), .B1(new_n1042), .B2(new_n1043), .ZN(G72));
  NAND2_X1  g858(.A1(new_n337), .A2(new_n349), .ZN(new_n1045));
  XNOR2_X1  g859(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1046));
  NOR2_X1   g860(.A1(new_n659), .A2(new_n330), .ZN(new_n1047));
  XNOR2_X1  g861(.A(new_n1046), .B(new_n1047), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g863(.A(new_n1049), .B(KEYINPUT127), .ZN(new_n1050));
  NAND3_X1  g864(.A1(new_n938), .A2(new_n939), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1051), .A2(new_n963), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n299), .A2(new_n290), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n1048), .B1(new_n1033), .B2(new_n1002), .ZN(new_n1054));
  OR2_X1    g868(.A1(new_n1054), .A2(KEYINPUT126), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1054), .A2(KEYINPUT126), .ZN(new_n1056));
  AOI21_X1  g870(.A(new_n1053), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g871(.A(new_n727), .ZN(new_n1058));
  OR2_X1    g872(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1059));
  OAI21_X1  g873(.A(new_n1048), .B1(new_n1059), .B2(new_n1002), .ZN(new_n1060));
  AOI211_X1 g874(.A(new_n1052), .B(new_n1057), .C1(new_n1058), .C2(new_n1060), .ZN(G57));
endmodule


