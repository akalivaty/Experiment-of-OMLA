

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592;

  XNOR2_X1 U326 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U327 ( .A(KEYINPUT93), .B(KEYINPUT21), .Z(n294) );
  XNOR2_X1 U328 ( .A(n350), .B(n349), .ZN(n351) );
  NOR2_X1 U329 ( .A1(n586), .A2(n481), .ZN(n482) );
  XNOR2_X1 U330 ( .A(n352), .B(n351), .ZN(n357) );
  XNOR2_X1 U331 ( .A(n442), .B(n390), .ZN(n392) );
  XOR2_X1 U332 ( .A(n581), .B(n358), .Z(n565) );
  AND2_X1 U333 ( .A1(n461), .A2(n541), .ZN(n571) );
  INV_X1 U334 ( .A(G106GAT), .ZN(n487) );
  XOR2_X1 U335 ( .A(n398), .B(n397), .Z(n530) );
  XNOR2_X1 U336 ( .A(KEYINPUT124), .B(G183GAT), .ZN(n462) );
  XNOR2_X1 U337 ( .A(n487), .B(KEYINPUT44), .ZN(n488) );
  XNOR2_X1 U338 ( .A(n484), .B(KEYINPUT116), .ZN(n485) );
  XNOR2_X1 U339 ( .A(n463), .B(n462), .ZN(G1350GAT) );
  XNOR2_X1 U340 ( .A(n486), .B(n485), .ZN(G1336GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT14), .B(KEYINPUT87), .Z(n296) );
  XNOR2_X1 U342 ( .A(G155GAT), .B(KEYINPUT82), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U344 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n298) );
  XNOR2_X1 U345 ( .A(G22GAT), .B(G71GAT), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U347 ( .A(n300), .B(n299), .ZN(n315) );
  XOR2_X1 U348 ( .A(KEYINPUT86), .B(KEYINPUT84), .Z(n302) );
  XNOR2_X1 U349 ( .A(G127GAT), .B(KEYINPUT85), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U351 ( .A(G78GAT), .B(G64GAT), .Z(n304) );
  XOR2_X1 U352 ( .A(G15GAT), .B(G1GAT), .Z(n316) );
  XOR2_X1 U353 ( .A(G8GAT), .B(G183GAT), .Z(n396) );
  XNOR2_X1 U354 ( .A(n316), .B(n396), .ZN(n303) );
  XNOR2_X1 U355 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U356 ( .A(n306), .B(n305), .Z(n308) );
  NAND2_X1 U357 ( .A1(G231GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U358 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U359 ( .A(n309), .B(KEYINPUT83), .Z(n313) );
  XOR2_X1 U360 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n311) );
  XNOR2_X1 U361 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n355) );
  XNOR2_X1 U363 ( .A(n355), .B(G211GAT), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n315), .B(n314), .ZN(n586) );
  XOR2_X1 U366 ( .A(G36GAT), .B(G50GAT), .Z(n318) );
  XOR2_X1 U367 ( .A(G141GAT), .B(G22GAT), .Z(n430) );
  XNOR2_X1 U368 ( .A(n316), .B(n430), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U370 ( .A(n319), .B(G113GAT), .Z(n324) );
  XOR2_X1 U371 ( .A(KEYINPUT71), .B(KEYINPUT69), .Z(n321) );
  XNOR2_X1 U372 ( .A(G8GAT), .B(G197GAT), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U374 ( .A(G169GAT), .B(n322), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U376 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n326) );
  NAND2_X1 U377 ( .A1(G229GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U379 ( .A(n328), .B(n327), .Z(n333) );
  XOR2_X1 U380 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n330) );
  XNOR2_X1 U381 ( .A(G43GAT), .B(G29GAT), .ZN(n329) );
  XNOR2_X1 U382 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U383 ( .A(KEYINPUT72), .B(n331), .Z(n375) );
  XNOR2_X1 U384 ( .A(n375), .B(KEYINPUT70), .ZN(n332) );
  XNOR2_X1 U385 ( .A(n333), .B(n332), .ZN(n563) );
  INV_X1 U386 ( .A(G78GAT), .ZN(n334) );
  NAND2_X1 U387 ( .A1(n334), .A2(KEYINPUT76), .ZN(n337) );
  INV_X1 U388 ( .A(KEYINPUT76), .ZN(n335) );
  NAND2_X1 U389 ( .A1(n335), .A2(G78GAT), .ZN(n336) );
  NAND2_X1 U390 ( .A1(n337), .A2(n336), .ZN(n339) );
  XNOR2_X1 U391 ( .A(G148GAT), .B(G106GAT), .ZN(n338) );
  XNOR2_X1 U392 ( .A(n339), .B(n338), .ZN(n436) );
  INV_X1 U393 ( .A(n436), .ZN(n340) );
  XOR2_X1 U394 ( .A(G99GAT), .B(G85GAT), .Z(n363) );
  NAND2_X1 U395 ( .A1(n340), .A2(n363), .ZN(n343) );
  INV_X1 U396 ( .A(n363), .ZN(n341) );
  NAND2_X1 U397 ( .A1(n436), .A2(n341), .ZN(n342) );
  NAND2_X1 U398 ( .A1(n343), .A2(n342), .ZN(n345) );
  NAND2_X1 U399 ( .A1(G230GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U400 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U401 ( .A(n346), .B(KEYINPUT75), .Z(n352) );
  XOR2_X1 U402 ( .A(G120GAT), .B(G71GAT), .Z(n454) );
  XNOR2_X1 U403 ( .A(n454), .B(KEYINPUT33), .ZN(n350) );
  XOR2_X1 U404 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n348) );
  XNOR2_X1 U405 ( .A(KEYINPUT78), .B(KEYINPUT77), .ZN(n347) );
  XNOR2_X1 U406 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U407 ( .A(G204GAT), .B(G64GAT), .Z(n354) );
  XNOR2_X1 U408 ( .A(G176GAT), .B(G92GAT), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n391) );
  XNOR2_X1 U410 ( .A(n355), .B(n391), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n357), .B(n356), .ZN(n581) );
  XOR2_X1 U412 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n358) );
  NAND2_X1 U413 ( .A1(n563), .A2(n565), .ZN(n359) );
  XOR2_X1 U414 ( .A(n359), .B(KEYINPUT46), .Z(n360) );
  NOR2_X1 U415 ( .A1(n586), .A2(n360), .ZN(n376) );
  XOR2_X1 U416 ( .A(KEYINPUT81), .B(KEYINPUT9), .Z(n362) );
  XNOR2_X1 U417 ( .A(G106GAT), .B(G92GAT), .ZN(n361) );
  XNOR2_X1 U418 ( .A(n362), .B(n361), .ZN(n367) );
  XOR2_X1 U419 ( .A(G218GAT), .B(n363), .Z(n365) );
  XOR2_X1 U420 ( .A(G36GAT), .B(G190GAT), .Z(n389) );
  XNOR2_X1 U421 ( .A(G134GAT), .B(n389), .ZN(n364) );
  XNOR2_X1 U422 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U423 ( .A(n367), .B(n366), .Z(n369) );
  NAND2_X1 U424 ( .A1(G232GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U425 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U426 ( .A(n370), .B(KEYINPUT10), .Z(n373) );
  XNOR2_X1 U427 ( .A(G50GAT), .B(G162GAT), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n371), .B(KEYINPUT80), .ZN(n437) );
  XNOR2_X1 U429 ( .A(n437), .B(KEYINPUT11), .ZN(n372) );
  XNOR2_X1 U430 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n491) );
  NAND2_X1 U432 ( .A1(n376), .A2(n491), .ZN(n378) );
  XOR2_X1 U433 ( .A(KEYINPUT117), .B(KEYINPUT47), .Z(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n384) );
  XOR2_X1 U435 ( .A(KEYINPUT67), .B(KEYINPUT45), .Z(n380) );
  INV_X1 U436 ( .A(n491), .ZN(n570) );
  XNOR2_X1 U437 ( .A(n570), .B(KEYINPUT36), .ZN(n588) );
  NAND2_X1 U438 ( .A1(n586), .A2(n588), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n382) );
  INV_X1 U440 ( .A(n563), .ZN(n577) );
  NAND2_X1 U441 ( .A1(n581), .A2(n577), .ZN(n381) );
  NOR2_X1 U442 ( .A1(n382), .A2(n381), .ZN(n383) );
  NOR2_X1 U443 ( .A1(n384), .A2(n383), .ZN(n385) );
  XNOR2_X1 U444 ( .A(n385), .B(KEYINPUT48), .ZN(n536) );
  XNOR2_X1 U445 ( .A(G197GAT), .B(G218GAT), .ZN(n386) );
  XNOR2_X1 U446 ( .A(n294), .B(n386), .ZN(n387) );
  XNOR2_X1 U447 ( .A(G211GAT), .B(n387), .ZN(n442) );
  NAND2_X1 U448 ( .A1(G226GAT), .A2(G233GAT), .ZN(n388) );
  XOR2_X1 U449 ( .A(n392), .B(n391), .Z(n398) );
  XOR2_X1 U450 ( .A(KEYINPUT90), .B(KEYINPUT18), .Z(n394) );
  XNOR2_X1 U451 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U453 ( .A(KEYINPUT19), .B(n395), .Z(n458) );
  XNOR2_X1 U454 ( .A(n458), .B(n396), .ZN(n397) );
  XNOR2_X1 U455 ( .A(KEYINPUT122), .B(n530), .ZN(n399) );
  NOR2_X1 U456 ( .A1(n536), .A2(n399), .ZN(n400) );
  XNOR2_X1 U457 ( .A(n400), .B(KEYINPUT54), .ZN(n427) );
  XOR2_X1 U458 ( .A(G85GAT), .B(G162GAT), .Z(n403) );
  XNOR2_X1 U459 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n401), .B(KEYINPUT2), .ZN(n429) );
  XNOR2_X1 U461 ( .A(G57GAT), .B(n429), .ZN(n402) );
  XNOR2_X1 U462 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U463 ( .A(G29GAT), .B(n404), .ZN(n426) );
  XOR2_X1 U464 ( .A(KEYINPUT5), .B(KEYINPUT95), .Z(n406) );
  XNOR2_X1 U465 ( .A(KEYINPUT96), .B(KEYINPUT6), .ZN(n405) );
  XNOR2_X1 U466 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U467 ( .A(G148GAT), .B(G120GAT), .Z(n408) );
  XNOR2_X1 U468 ( .A(G1GAT), .B(G141GAT), .ZN(n407) );
  XNOR2_X1 U469 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n410), .B(n409), .ZN(n424) );
  XOR2_X1 U471 ( .A(KEYINPUT100), .B(KEYINPUT97), .Z(n412) );
  XNOR2_X1 U472 ( .A(KEYINPUT99), .B(KEYINPUT98), .ZN(n411) );
  XNOR2_X1 U473 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U474 ( .A(KEYINPUT101), .B(n413), .Z(n415) );
  NAND2_X1 U475 ( .A1(G225GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U476 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U477 ( .A(n416), .B(KEYINPUT1), .Z(n422) );
  XOR2_X1 U478 ( .A(G134GAT), .B(KEYINPUT0), .Z(n418) );
  XNOR2_X1 U479 ( .A(G113GAT), .B(KEYINPUT89), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U481 ( .A(G127GAT), .B(n419), .ZN(n459) );
  INV_X1 U482 ( .A(n459), .ZN(n420) );
  XNOR2_X1 U483 ( .A(n420), .B(KEYINPUT4), .ZN(n421) );
  XNOR2_X1 U484 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n426), .B(n425), .ZN(n535) );
  NAND2_X1 U487 ( .A1(n427), .A2(n535), .ZN(n428) );
  XNOR2_X1 U488 ( .A(n428), .B(KEYINPUT65), .ZN(n576) );
  XOR2_X1 U489 ( .A(KEYINPUT23), .B(G204GAT), .Z(n432) );
  XNOR2_X1 U490 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U491 ( .A(n432), .B(n431), .ZN(n441) );
  XOR2_X1 U492 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n434) );
  NAND2_X1 U493 ( .A1(G228GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U494 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U495 ( .A(n435), .B(KEYINPUT94), .Z(n439) );
  XNOR2_X1 U496 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U497 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n472) );
  NAND2_X1 U500 ( .A1(n576), .A2(n472), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n444), .B(KEYINPUT55), .ZN(n461) );
  XOR2_X1 U502 ( .A(G176GAT), .B(G99GAT), .Z(n446) );
  XNOR2_X1 U503 ( .A(G43GAT), .B(G190GAT), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U505 ( .A(KEYINPUT92), .B(KEYINPUT66), .Z(n448) );
  XNOR2_X1 U506 ( .A(G15GAT), .B(G183GAT), .ZN(n447) );
  XNOR2_X1 U507 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U508 ( .A(n450), .B(n449), .Z(n456) );
  XOR2_X1 U509 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n452) );
  NAND2_X1 U510 ( .A1(G227GAT), .A2(G233GAT), .ZN(n451) );
  XNOR2_X1 U511 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U512 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U513 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U514 ( .A(n458), .B(n457), .ZN(n460) );
  XOR2_X1 U515 ( .A(n460), .B(n459), .Z(n541) );
  NAND2_X1 U516 ( .A1(n571), .A2(n586), .ZN(n463) );
  AND2_X1 U517 ( .A1(n577), .A2(n565), .ZN(n519) );
  XOR2_X1 U518 ( .A(KEYINPUT28), .B(KEYINPUT68), .Z(n464) );
  XOR2_X1 U519 ( .A(n472), .B(n464), .Z(n540) );
  XNOR2_X1 U520 ( .A(n530), .B(KEYINPUT102), .ZN(n465) );
  XOR2_X1 U521 ( .A(KEYINPUT27), .B(n465), .Z(n538) );
  AND2_X1 U522 ( .A1(n540), .A2(n538), .ZN(n466) );
  INV_X1 U523 ( .A(n541), .ZN(n533) );
  NAND2_X1 U524 ( .A1(n466), .A2(n533), .ZN(n467) );
  NOR2_X1 U525 ( .A1(n535), .A2(n467), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n468), .B(KEYINPUT103), .ZN(n480) );
  NOR2_X1 U527 ( .A1(n541), .A2(n472), .ZN(n470) );
  XNOR2_X1 U528 ( .A(KEYINPUT26), .B(KEYINPUT104), .ZN(n469) );
  XNOR2_X1 U529 ( .A(n470), .B(n469), .ZN(n575) );
  NAND2_X1 U530 ( .A1(n575), .A2(n538), .ZN(n471) );
  XOR2_X1 U531 ( .A(KEYINPUT105), .B(n471), .Z(n477) );
  OR2_X1 U532 ( .A1(n530), .A2(n533), .ZN(n473) );
  NAND2_X1 U533 ( .A1(n473), .A2(n472), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n474), .B(KEYINPUT106), .ZN(n475) );
  XOR2_X1 U535 ( .A(KEYINPUT25), .B(n475), .Z(n476) );
  NAND2_X1 U536 ( .A1(n477), .A2(n476), .ZN(n478) );
  NAND2_X1 U537 ( .A1(n478), .A2(n535), .ZN(n479) );
  NAND2_X1 U538 ( .A1(n480), .A2(n479), .ZN(n495) );
  NAND2_X1 U539 ( .A1(n588), .A2(n495), .ZN(n481) );
  XOR2_X1 U540 ( .A(KEYINPUT37), .B(n482), .Z(n505) );
  NAND2_X1 U541 ( .A1(n519), .A2(n505), .ZN(n483) );
  XOR2_X1 U542 ( .A(KEYINPUT115), .B(n483), .Z(n532) );
  NOR2_X1 U543 ( .A1(n535), .A2(n532), .ZN(n486) );
  INV_X1 U544 ( .A(G85GAT), .ZN(n484) );
  NOR2_X1 U545 ( .A1(n540), .A2(n532), .ZN(n489) );
  XNOR2_X1 U546 ( .A(n489), .B(n488), .ZN(G1339GAT) );
  NAND2_X1 U547 ( .A1(n581), .A2(n563), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n490), .B(KEYINPUT79), .ZN(n506) );
  XOR2_X1 U549 ( .A(KEYINPUT88), .B(KEYINPUT16), .Z(n493) );
  NAND2_X1 U550 ( .A1(n586), .A2(n491), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n493), .B(n492), .ZN(n494) );
  NAND2_X1 U552 ( .A1(n495), .A2(n494), .ZN(n496) );
  XNOR2_X1 U553 ( .A(n496), .B(KEYINPUT107), .ZN(n518) );
  NAND2_X1 U554 ( .A1(n506), .A2(n518), .ZN(n503) );
  NOR2_X1 U555 ( .A1(n535), .A2(n503), .ZN(n498) );
  XNOR2_X1 U556 ( .A(KEYINPUT34), .B(KEYINPUT108), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U558 ( .A(G1GAT), .B(n499), .Z(G1324GAT) );
  NOR2_X1 U559 ( .A1(n530), .A2(n503), .ZN(n500) );
  XOR2_X1 U560 ( .A(G8GAT), .B(n500), .Z(G1325GAT) );
  NOR2_X1 U561 ( .A1(n533), .A2(n503), .ZN(n502) );
  XNOR2_X1 U562 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(G1326GAT) );
  NOR2_X1 U564 ( .A1(n540), .A2(n503), .ZN(n504) );
  XOR2_X1 U565 ( .A(G22GAT), .B(n504), .Z(G1327GAT) );
  NAND2_X1 U566 ( .A1(n506), .A2(n505), .ZN(n507) );
  XNOR2_X1 U567 ( .A(n507), .B(KEYINPUT38), .ZN(n514) );
  NOR2_X1 U568 ( .A1(n535), .A2(n514), .ZN(n508) );
  XNOR2_X1 U569 ( .A(n508), .B(KEYINPUT39), .ZN(n509) );
  XNOR2_X1 U570 ( .A(G29GAT), .B(n509), .ZN(G1328GAT) );
  NOR2_X1 U571 ( .A1(n514), .A2(n530), .ZN(n510) );
  XOR2_X1 U572 ( .A(G36GAT), .B(n510), .Z(G1329GAT) );
  NOR2_X1 U573 ( .A1(n514), .A2(n533), .ZN(n512) );
  XNOR2_X1 U574 ( .A(KEYINPUT40), .B(KEYINPUT109), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U576 ( .A(G43GAT), .B(n513), .ZN(G1330GAT) );
  NOR2_X1 U577 ( .A1(n514), .A2(n540), .ZN(n515) );
  XOR2_X1 U578 ( .A(G50GAT), .B(n515), .Z(G1331GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n517) );
  XNOR2_X1 U580 ( .A(G57GAT), .B(KEYINPUT110), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(n521) );
  NAND2_X1 U582 ( .A1(n519), .A2(n518), .ZN(n527) );
  NOR2_X1 U583 ( .A1(n535), .A2(n527), .ZN(n520) );
  XOR2_X1 U584 ( .A(n521), .B(n520), .Z(G1332GAT) );
  NOR2_X1 U585 ( .A1(n530), .A2(n527), .ZN(n522) );
  XOR2_X1 U586 ( .A(KEYINPUT112), .B(n522), .Z(n523) );
  XNOR2_X1 U587 ( .A(G64GAT), .B(n523), .ZN(G1333GAT) );
  NOR2_X1 U588 ( .A1(n533), .A2(n527), .ZN(n525) );
  XNOR2_X1 U589 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G71GAT), .B(n526), .ZN(G1334GAT) );
  NOR2_X1 U592 ( .A1(n540), .A2(n527), .ZN(n529) );
  XNOR2_X1 U593 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n529), .B(n528), .ZN(G1335GAT) );
  NOR2_X1 U595 ( .A1(n530), .A2(n532), .ZN(n531) );
  XOR2_X1 U596 ( .A(G92GAT), .B(n531), .Z(G1337GAT) );
  NOR2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U598 ( .A(G99GAT), .B(n534), .Z(G1338GAT) );
  XOR2_X1 U599 ( .A(G113GAT), .B(KEYINPUT119), .Z(n544) );
  NOR2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U601 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U602 ( .A(KEYINPUT118), .B(n539), .ZN(n554) );
  NAND2_X1 U603 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U604 ( .A1(n554), .A2(n542), .ZN(n550) );
  NAND2_X1 U605 ( .A1(n550), .A2(n563), .ZN(n543) );
  XNOR2_X1 U606 ( .A(n544), .B(n543), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT49), .B(KEYINPUT120), .Z(n546) );
  NAND2_X1 U608 ( .A1(n550), .A2(n565), .ZN(n545) );
  XNOR2_X1 U609 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U610 ( .A(G120GAT), .B(n547), .ZN(G1341GAT) );
  NAND2_X1 U611 ( .A1(n550), .A2(n586), .ZN(n548) );
  XNOR2_X1 U612 ( .A(n548), .B(KEYINPUT50), .ZN(n549) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n549), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT51), .Z(n552) );
  NAND2_X1 U615 ( .A1(n550), .A2(n570), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(G1343GAT) );
  INV_X1 U617 ( .A(n575), .ZN(n553) );
  NOR2_X1 U618 ( .A1(n554), .A2(n553), .ZN(n560) );
  NAND2_X1 U619 ( .A1(n563), .A2(n560), .ZN(n555) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n555), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n557) );
  NAND2_X1 U622 ( .A1(n560), .A2(n565), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n560), .A2(n586), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U627 ( .A(G162GAT), .B(KEYINPUT121), .Z(n562) );
  NAND2_X1 U628 ( .A1(n560), .A2(n570), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1347GAT) );
  NAND2_X1 U630 ( .A1(n571), .A2(n563), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U632 ( .A1(n571), .A2(n565), .ZN(n567) );
  XOR2_X1 U633 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n569) );
  XOR2_X1 U635 ( .A(G176GAT), .B(KEYINPUT56), .Z(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n573) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(G190GAT), .B(n574), .ZN(G1351GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n585) );
  NOR2_X1 U642 ( .A1(n577), .A2(n585), .ZN(n579) );
  XNOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(n580), .ZN(G1352GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n585), .ZN(n583) );
  XNOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(G204GAT), .B(n584), .ZN(G1353GAT) );
  INV_X1 U650 ( .A(n585), .ZN(n589) );
  AND2_X1 U651 ( .A1(n586), .A2(n589), .ZN(n587) );
  XOR2_X1 U652 ( .A(G211GAT), .B(n587), .Z(G1354GAT) );
  XOR2_X1 U653 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n591) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

