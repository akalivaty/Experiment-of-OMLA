//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT64), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AND2_X1   g0014(.A1(new_n212), .A2(new_n213), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n214), .B(new_n215), .C1(G77), .C2(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G116), .ZN(new_n219));
  INV_X1    g0019(.A(G270), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G50), .ZN(new_n222));
  INV_X1    g0022(.A(G226), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n203), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(G58), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(new_n217), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n206), .B(new_n226), .C1(new_n229), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G264), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n220), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(KEYINPUT65), .B(G107), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n219), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  NAND3_X1  g0050(.A1(new_n222), .A2(new_n230), .A3(new_n217), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  AOI22_X1  g0052(.A1(new_n251), .A2(G20), .B1(G150), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n230), .A2(KEYINPUT68), .A3(KEYINPUT8), .ZN(new_n254));
  XOR2_X1   g0054(.A(KEYINPUT8), .B(G58), .Z(new_n255));
  OAI21_X1  g0055(.A(new_n254), .B1(new_n255), .B2(KEYINPUT68), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n228), .A2(G33), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n253), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n227), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n258), .A2(new_n260), .B1(new_n222), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n260), .B1(new_n261), .B2(G20), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n264), .B1(new_n222), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n268));
  AND2_X1   g0068(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n269));
  OR3_X1    g0069(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n267), .A2(KEYINPUT76), .A3(KEYINPUT9), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G222), .ZN(new_n279));
  INV_X1    g0079(.A(G223), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n277), .B(new_n279), .C1(new_n280), .C2(new_n278), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(G77), .B2(new_n277), .ZN(new_n282));
  XOR2_X1   g0082(.A(new_n282), .B(KEYINPUT67), .Z(new_n283));
  AND2_X1   g0083(.A1(G33), .A2(G41), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(new_n227), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  INV_X1    g0087(.A(G45), .ZN(new_n288));
  AOI21_X1  g0088(.A(G1), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT66), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n290), .B1(new_n284), .B2(new_n227), .ZN(new_n291));
  AND2_X1   g0091(.A1(G1), .A2(G13), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(KEYINPUT66), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n289), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G274), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(new_n291), .B2(new_n294), .ZN(new_n297));
  AOI22_X1  g0097(.A1(G226), .A2(new_n295), .B1(new_n297), .B2(new_n289), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n286), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(KEYINPUT74), .B(G200), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n286), .A2(G190), .A3(new_n298), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n272), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT77), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n272), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n270), .A2(KEYINPUT77), .A3(new_n271), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  XOR2_X1   g0108(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n309));
  NAND3_X1  g0109(.A1(new_n301), .A2(new_n302), .A3(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n304), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NOR3_X1   g0111(.A1(new_n284), .A2(new_n290), .A3(new_n227), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT66), .B1(new_n292), .B2(new_n293), .ZN(new_n313));
  OAI211_X1 g0113(.A(G274), .B(new_n289), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n295), .ZN(new_n315));
  INV_X1    g0115(.A(G244), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT70), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AND2_X1   g0119(.A1(KEYINPUT3), .A2(G33), .ZN(new_n320));
  NOR2_X1   g0120(.A1(KEYINPUT3), .A2(G33), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n322), .B1(G238), .B2(G1698), .ZN(new_n323));
  INV_X1    g0123(.A(G232), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(G1698), .ZN(new_n325));
  OR2_X1    g0125(.A1(KEYINPUT71), .A2(G107), .ZN(new_n326));
  NAND2_X1  g0126(.A1(KEYINPUT71), .A2(G107), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n325), .B(new_n285), .C1(new_n277), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n317), .A2(new_n318), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n319), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  XOR2_X1   g0133(.A(KEYINPUT69), .B(G179), .Z(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G169), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G77), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n263), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n265), .A2(G77), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G20), .A2(G77), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT72), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n252), .B(new_n343), .ZN(new_n344));
  XNOR2_X1  g0144(.A(KEYINPUT8), .B(G58), .ZN(new_n345));
  XOR2_X1   g0145(.A(KEYINPUT15), .B(G87), .Z(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n342), .B1(new_n344), .B2(new_n345), .C1(new_n257), .C2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT73), .ZN(new_n349));
  AND3_X1   g0149(.A1(new_n348), .A2(new_n349), .A3(new_n260), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n349), .B1(new_n348), .B2(new_n260), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n340), .B(new_n341), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n336), .A2(new_n338), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n352), .B1(new_n332), .B2(new_n300), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT75), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n355), .A2(new_n356), .B1(G190), .B2(new_n333), .ZN(new_n357));
  INV_X1    g0157(.A(new_n352), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n332), .A2(new_n300), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT75), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n354), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n299), .A2(new_n337), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n363), .B(new_n267), .C1(new_n334), .C2(new_n299), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n311), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT82), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT16), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT7), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n277), .B2(G20), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n322), .A2(KEYINPUT7), .A3(new_n228), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n217), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(G58), .A2(G68), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT81), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT81), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n374), .A2(G58), .A3(G68), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n375), .A3(new_n231), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G20), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n252), .A2(G159), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n367), .B1(new_n371), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT7), .B1(new_n322), .B2(new_n228), .ZN(new_n381));
  NOR4_X1   g0181(.A1(new_n320), .A2(new_n321), .A3(new_n368), .A4(G20), .ZN(new_n382));
  OAI21_X1  g0182(.A(G68), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n376), .A2(G20), .B1(G159), .B2(new_n252), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(KEYINPUT16), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n380), .A2(new_n260), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n256), .A2(new_n263), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n266), .B2(new_n256), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n285), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n280), .A2(new_n278), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n277), .B(new_n391), .C1(G226), .C2(new_n278), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G87), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n390), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n295), .A2(G232), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n395), .A2(G190), .A3(new_n314), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n314), .ZN(new_n398));
  OAI21_X1  g0198(.A(G200), .B1(new_n398), .B2(new_n394), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n386), .A2(new_n389), .A3(new_n397), .A4(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT17), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n400), .A2(new_n401), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n366), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n260), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n383), .A2(new_n384), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n405), .B1(new_n406), .B2(new_n367), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n388), .B1(new_n407), .B2(new_n385), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n408), .A2(KEYINPUT17), .A3(new_n399), .A4(new_n397), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n400), .A2(new_n401), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT82), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n404), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n252), .ZN(new_n413));
  OAI22_X1  g0213(.A1(new_n413), .A2(new_n222), .B1(new_n228), .B2(G68), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n257), .A2(new_n339), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n260), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT11), .ZN(new_n417));
  OR3_X1    g0217(.A1(new_n262), .A2(KEYINPUT12), .A3(G68), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT12), .B1(new_n262), .B2(G68), .ZN(new_n419));
  AOI22_X1  g0219(.A1(G68), .A2(new_n265), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n289), .ZN(new_n423));
  OAI211_X1 g0223(.A(G238), .B(new_n423), .C1(new_n312), .C2(new_n313), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n314), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n223), .A2(new_n278), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n324), .A2(G1698), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n426), .B(new_n427), .C1(new_n320), .C2(new_n321), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n274), .A2(new_n210), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n390), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT13), .B1(new_n425), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n428), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n285), .B1(new_n433), .B2(new_n429), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT13), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n434), .A2(new_n435), .A3(new_n314), .A4(new_n424), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(G200), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n422), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G190), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n432), .A2(KEYINPUT79), .A3(new_n436), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n425), .A2(new_n431), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT79), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(new_n443), .A3(new_n435), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n440), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n439), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n441), .A2(new_n444), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G179), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT80), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(KEYINPUT14), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n437), .B2(new_n337), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n449), .A2(KEYINPUT14), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n432), .A2(new_n436), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n454), .A2(G169), .A3(new_n450), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n448), .A2(new_n452), .A3(new_n453), .A4(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n446), .B1(new_n456), .B2(new_n421), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n395), .A2(new_n335), .A3(new_n314), .A4(new_n396), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n337), .B1(new_n398), .B2(new_n394), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n386), .A2(new_n389), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT18), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT18), .B1(new_n460), .B2(new_n461), .ZN(new_n463));
  OR2_X1    g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n412), .A2(new_n457), .A3(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n365), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n261), .A2(G33), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n262), .A2(new_n468), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n469), .A2(new_n219), .A3(new_n260), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT20), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n228), .B1(new_n210), .B2(G33), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT84), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(G33), .A3(G283), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT84), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n472), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n260), .B1(new_n228), .B2(G116), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n471), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n476), .A2(new_n474), .ZN(new_n480));
  INV_X1    g0280(.A(new_n472), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n259), .A2(new_n227), .B1(G20), .B2(new_n219), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(KEYINPUT20), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n470), .B1(new_n479), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n262), .A2(G116), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n337), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G264), .A2(G1698), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n277), .B(new_n489), .C1(new_n211), .C2(G1698), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n490), .B(new_n285), .C1(G303), .C2(new_n277), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n261), .A2(G45), .ZN(new_n492));
  OR2_X1    g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  NAND2_X1  g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n495), .B1(new_n291), .B2(new_n294), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G270), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n495), .B(G274), .C1(new_n312), .C2(new_n313), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT85), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT85), .B1(new_n297), .B2(new_n495), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n491), .B(new_n497), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n488), .A2(KEYINPUT21), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT21), .B1(new_n488), .B2(new_n502), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n498), .A2(new_n499), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n297), .A2(KEYINPUT85), .A3(new_n495), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n507), .A2(G179), .A3(new_n491), .A4(new_n497), .ZN(new_n508));
  AOI211_X1 g0308(.A(new_n486), .B(new_n470), .C1(new_n479), .C2(new_n484), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n503), .A2(new_n504), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n346), .A2(new_n262), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n328), .A2(new_n208), .A3(new_n210), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n513), .B(KEYINPUT19), .C1(G20), .C2(new_n429), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n277), .A2(new_n228), .A3(G68), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT19), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n430), .B2(G20), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n512), .B1(new_n518), .B2(new_n260), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n469), .A2(new_n260), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n346), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n218), .A2(new_n278), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n277), .B(new_n522), .C1(G244), .C2(new_n278), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G116), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n285), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n291), .A2(new_n294), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n492), .A2(new_n209), .ZN(new_n528));
  INV_X1    g0328(.A(new_n492), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n296), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n519), .A2(new_n521), .B1(new_n337), .B2(new_n532), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n526), .A2(new_n531), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n335), .ZN(new_n535));
  INV_X1    g0335(.A(new_n300), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n536), .B1(new_n526), .B2(new_n531), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n537), .B1(G190), .B2(new_n534), .ZN(new_n538));
  INV_X1    g0338(.A(new_n520), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(new_n208), .ZN(new_n540));
  AOI211_X1 g0340(.A(new_n512), .B(new_n540), .C1(new_n518), .C2(new_n260), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n533), .A2(new_n535), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n502), .A2(G200), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n543), .B(new_n509), .C1(new_n440), .C2(new_n502), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n277), .A2(new_n228), .A3(G87), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT22), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT22), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n277), .A2(new_n547), .A3(new_n228), .A4(G87), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT23), .ZN(new_n549));
  INV_X1    g0349(.A(G107), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(G20), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n524), .A2(G20), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n228), .B1(new_n326), .B2(new_n327), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n551), .B(new_n553), .C1(new_n554), .C2(new_n549), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT88), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g0357(.A1(KEYINPUT71), .A2(G107), .ZN(new_n558));
  NOR2_X1   g0358(.A1(KEYINPUT71), .A2(G107), .ZN(new_n559));
  OAI21_X1  g0359(.A(G20), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n552), .B1(new_n560), .B2(KEYINPUT23), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n561), .A2(KEYINPUT88), .A3(new_n551), .ZN(new_n562));
  AOI221_X4 g0362(.A(KEYINPUT24), .B1(new_n546), .B2(new_n548), .C1(new_n557), .C2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT24), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n557), .A2(new_n562), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n546), .A2(new_n548), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n260), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n209), .A2(new_n278), .ZN(new_n569));
  OAI221_X1 g0369(.A(new_n569), .B1(G257), .B2(new_n278), .C1(new_n320), .C2(new_n321), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G33), .A2(G294), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n496), .A2(G264), .B1(new_n572), .B2(new_n285), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n507), .A2(new_n573), .A3(new_n440), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n493), .A2(new_n494), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n529), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n527), .A2(G264), .A3(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n275), .A2(new_n276), .B1(new_n211), .B2(G1698), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n578), .A2(new_n569), .B1(G33), .B2(G294), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n577), .B1(new_n579), .B2(new_n390), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n505), .B2(new_n506), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n574), .B1(new_n581), .B2(G200), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT25), .B1(new_n263), .B2(new_n550), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n263), .A2(KEYINPUT25), .A3(new_n550), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n584), .A2(new_n585), .B1(G107), .B2(new_n520), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n568), .A2(new_n582), .A3(new_n586), .ZN(new_n587));
  AND4_X1   g0387(.A1(new_n511), .A2(new_n542), .A3(new_n544), .A4(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(G169), .B1(new_n507), .B2(new_n573), .ZN(new_n589));
  INV_X1    g0389(.A(G179), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n589), .B1(new_n590), .B2(new_n581), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n555), .A2(new_n556), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT88), .B1(new_n561), .B2(new_n551), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n566), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT24), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n565), .A2(new_n564), .A3(new_n566), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n405), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n586), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n591), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n316), .A2(G1698), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n320), .B2(new_n321), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT4), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n277), .A2(G250), .A3(G1698), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n600), .B(KEYINPUT4), .C1(new_n321), .C2(new_n320), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n480), .A4(new_n605), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n606), .A2(new_n285), .B1(new_n496), .B2(G257), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n607), .A2(new_n335), .A3(new_n507), .ZN(new_n608));
  AOI21_X1  g0408(.A(G169), .B1(new_n607), .B2(new_n507), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n329), .B1(new_n381), .B2(new_n382), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT6), .ZN(new_n611));
  AND2_X1   g0411(.A1(G97), .A2(G107), .ZN(new_n612));
  NOR2_X1   g0412(.A1(G97), .A2(G107), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n550), .A2(KEYINPUT6), .A3(G97), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n616), .A2(G20), .B1(G77), .B2(new_n252), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n405), .B1(new_n610), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n262), .A2(G97), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(new_n520), .B2(G97), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n608), .A2(new_n609), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n607), .A2(new_n507), .ZN(new_n624));
  AOI21_X1  g0424(.A(KEYINPUT86), .B1(new_n624), .B2(G200), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT86), .ZN(new_n626));
  AOI211_X1 g0426(.A(new_n626), .B(new_n438), .C1(new_n607), .C2(new_n507), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT83), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n618), .B2(new_n621), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n614), .A2(new_n615), .ZN(new_n631));
  OAI22_X1  g0431(.A1(new_n631), .A2(new_n228), .B1(new_n339), .B2(new_n413), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n328), .B1(new_n369), .B2(new_n370), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n260), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(KEYINPUT83), .A3(new_n620), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n607), .A2(new_n507), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n630), .A2(new_n635), .B1(new_n636), .B2(G190), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n623), .B1(new_n628), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n638), .A2(KEYINPUT87), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n626), .B1(new_n636), .B2(new_n438), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n636), .A2(G190), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n635), .A2(new_n630), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n624), .A2(KEYINPUT86), .A3(G200), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n640), .A2(new_n641), .A3(new_n642), .A4(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n623), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n644), .A2(new_n645), .A3(KEYINPUT87), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n588), .B(new_n599), .C1(new_n639), .C2(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n467), .A2(new_n647), .ZN(G372));
  AOI22_X1  g0448(.A1(new_n447), .A2(G179), .B1(new_n449), .B2(KEYINPUT14), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n450), .B1(new_n454), .B2(G169), .ZN(new_n650));
  AOI211_X1 g0450(.A(new_n337), .B(new_n451), .C1(new_n432), .C2(new_n436), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n422), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n446), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n653), .B1(new_n354), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n412), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n464), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n311), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n658), .A2(new_n364), .ZN(new_n659));
  INV_X1    g0459(.A(new_n542), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n511), .A2(new_n599), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n661), .A2(new_n587), .A3(new_n638), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n608), .A2(new_n609), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n663), .A2(KEYINPUT90), .A3(new_n630), .A4(new_n635), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n624), .A2(new_n337), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n607), .A2(new_n335), .A3(new_n507), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n665), .A2(new_n666), .A3(new_n635), .A4(new_n630), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT90), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT26), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n664), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n660), .B1(new_n662), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n519), .A2(new_n521), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n532), .A2(new_n337), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(new_n535), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT89), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n533), .A2(KEYINPUT89), .A3(new_n535), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n542), .A2(new_n623), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n679), .B1(new_n681), .B2(new_n670), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n672), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n659), .B1(new_n467), .B2(new_n683), .ZN(G369));
  INV_X1    g0484(.A(G13), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n685), .A2(G1), .A3(G20), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT91), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT27), .ZN(new_n688));
  OR3_X1    g0488(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G213), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n690), .B1(new_n686), .B2(new_n688), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n687), .B1(new_n686), .B2(new_n688), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G343), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n509), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n511), .A2(new_n544), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n511), .B2(new_n698), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT92), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G330), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n507), .A2(new_n573), .A3(new_n590), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n581), .B2(G169), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n568), .B2(new_n586), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n695), .B1(new_n597), .B2(new_n598), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n706), .B1(new_n587), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n599), .A2(new_n695), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n703), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n511), .A2(new_n695), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n599), .B2(new_n695), .ZN(new_n715));
  OR2_X1    g0515(.A1(new_n712), .A2(new_n715), .ZN(G399));
  INV_X1    g0516(.A(new_n204), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(G41), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G1), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n513), .A2(G116), .ZN(new_n721));
  OAI22_X1  g0521(.A1(new_n720), .A2(new_n721), .B1(new_n232), .B2(new_n719), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT28), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n644), .A2(new_n645), .A3(new_n587), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n479), .A2(new_n484), .ZN(new_n725));
  INV_X1    g0525(.A(new_n470), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(new_n487), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n502), .A2(G169), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT21), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n507), .A2(new_n497), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(G179), .A3(new_n491), .A4(new_n727), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n488), .A2(KEYINPUT21), .A3(new_n502), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n730), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n706), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n671), .B1(new_n724), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n542), .ZN(new_n737));
  INV_X1    g0537(.A(new_n679), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n738), .B1(new_n680), .B2(KEYINPUT26), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n695), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT29), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n542), .A2(new_n670), .A3(new_n623), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n679), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n664), .A2(new_n669), .A3(new_n542), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n744), .B1(KEYINPUT26), .B2(new_n745), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n661), .A2(new_n542), .A3(new_n638), .A4(new_n587), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n695), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n742), .B1(new_n741), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT93), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n502), .A2(new_n335), .ZN(new_n751));
  INV_X1    g0551(.A(new_n581), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n751), .A2(new_n532), .A3(new_n752), .A4(new_n624), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n624), .A2(new_n532), .ZN(new_n754));
  INV_X1    g0554(.A(new_n508), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n754), .A2(new_n755), .A3(KEYINPUT30), .A4(new_n573), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT30), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n534), .A2(new_n607), .A3(new_n507), .A4(new_n573), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n757), .B1(new_n758), .B2(new_n508), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n753), .A2(new_n756), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n760), .A2(KEYINPUT31), .A3(new_n695), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(KEYINPUT31), .B1(new_n760), .B2(new_n695), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n750), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n763), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(KEYINPUT93), .A3(new_n761), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n764), .B(new_n766), .C1(new_n647), .C2(new_n695), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n767), .A2(G330), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n749), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n723), .B1(new_n769), .B2(G1), .ZN(G364));
  INV_X1    g0570(.A(KEYINPUT95), .ZN(new_n771));
  OAI21_X1  g0571(.A(G20), .B1(new_n771), .B2(G169), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n337), .A2(KEYINPUT95), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n292), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT96), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G190), .A2(G200), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n776), .A2(G20), .A3(new_n590), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G329), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n335), .A2(new_n228), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G190), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(KEYINPUT33), .B(G317), .Z(new_n784));
  NAND2_X1  g0584(.A1(new_n300), .A2(new_n590), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT99), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n228), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G190), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT101), .ZN(new_n789));
  INV_X1    g0589(.A(G303), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n779), .B1(new_n783), .B2(new_n784), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n787), .A2(new_n440), .ZN(new_n792));
  INV_X1    g0592(.A(G283), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n322), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n781), .A2(new_n440), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n440), .A2(G200), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n590), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n795), .A2(G326), .B1(G294), .B2(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT100), .Z(new_n800));
  NOR3_X1   g0600(.A1(new_n791), .A2(new_n794), .A3(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n780), .A2(new_n776), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n780), .A2(new_n796), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n804), .B1(G322), .B2(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT102), .Z(new_n808));
  INV_X1    g0608(.A(new_n795), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n792), .A2(new_n550), .B1(new_n809), .B2(new_n222), .ZN(new_n810));
  INV_X1    g0610(.A(new_n803), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n811), .A2(KEYINPUT98), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(KEYINPUT98), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n277), .B1(new_n208), .B2(new_n788), .C1(new_n814), .C2(new_n339), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n805), .B(KEYINPUT97), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n810), .B(new_n815), .C1(G58), .C2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G159), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n777), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT32), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n798), .A2(G97), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n817), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G68), .B2(new_n782), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n775), .B1(new_n808), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n249), .A2(G45), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n717), .A2(new_n277), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n825), .B(new_n826), .C1(G45), .C2(new_n232), .ZN(new_n827));
  INV_X1    g0627(.A(G355), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n277), .A2(new_n204), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n827), .B1(G116), .B2(new_n204), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT94), .ZN(new_n831));
  NOR2_X1   g0631(.A1(G13), .A2(G33), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(G20), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n775), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n685), .A2(G20), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n720), .B1(G45), .B2(new_n837), .ZN(new_n838));
  OR3_X1    g0638(.A1(new_n701), .A2(G20), .A3(new_n833), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n824), .A2(new_n836), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n701), .A2(G330), .ZN(new_n841));
  INV_X1    g0641(.A(new_n838), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n841), .A2(new_n702), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n840), .A2(new_n843), .ZN(G396));
  INV_X1    g0644(.A(G132), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n277), .B1(new_n777), .B2(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT104), .ZN(new_n847));
  INV_X1    g0647(.A(new_n814), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(G159), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n795), .A2(G137), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n816), .A2(G143), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n782), .A2(G150), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n849), .A2(new_n850), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n854), .A2(KEYINPUT34), .B1(new_n222), .B2(new_n789), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n847), .B(new_n855), .C1(KEYINPUT34), .C2(new_n854), .ZN(new_n856));
  INV_X1    g0656(.A(new_n798), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n856), .B1(new_n230), .B2(new_n857), .C1(new_n217), .C2(new_n792), .ZN(new_n858));
  INV_X1    g0658(.A(new_n789), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n859), .A2(G107), .B1(G311), .B2(new_n778), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n782), .A2(G283), .ZN(new_n861));
  INV_X1    g0661(.A(new_n792), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(G87), .ZN(new_n863));
  INV_X1    g0663(.A(G294), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n322), .B(new_n821), .C1(new_n805), .C2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(G303), .B2(new_n795), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n860), .A2(new_n861), .A3(new_n863), .A4(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n814), .A2(new_n219), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n858), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n360), .A2(KEYINPUT75), .B1(new_n440), .B2(new_n332), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n355), .A2(new_n356), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n870), .A2(new_n871), .B1(new_n358), .B2(new_n696), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n353), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n353), .A2(new_n695), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n869), .A2(new_n775), .B1(new_n832), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n775), .A2(new_n832), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n842), .B1(new_n878), .B2(new_n339), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT103), .Z(new_n880));
  NAND2_X1  g0680(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n362), .B(new_n696), .C1(new_n672), .C2(new_n682), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n874), .B1(new_n872), .B2(new_n353), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n882), .B1(new_n740), .B2(new_n883), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n768), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n842), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n881), .A2(new_n886), .ZN(G384));
  INV_X1    g0687(.A(new_n411), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT82), .B1(new_n409), .B2(new_n410), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n464), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT106), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n891), .B(new_n367), .C1(new_n371), .C2(new_n379), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n383), .B(new_n384), .C1(KEYINPUT106), .C2(KEYINPUT16), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n892), .A2(new_n893), .A3(new_n260), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n389), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT107), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n693), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n894), .A2(KEYINPUT107), .A3(new_n389), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n890), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n897), .A2(new_n460), .A3(new_n899), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n900), .A2(new_n903), .A3(new_n400), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n460), .A2(new_n461), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n906), .A2(new_n400), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT37), .ZN(new_n908));
  AOI211_X1 g0708(.A(KEYINPUT108), .B(new_n693), .C1(new_n386), .C2(new_n389), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT108), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n461), .B2(new_n898), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n907), .B(new_n908), .C1(new_n909), .C2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n905), .A2(new_n912), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n902), .A2(new_n913), .A3(KEYINPUT38), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n906), .B(new_n400), .C1(new_n911), .C2(new_n909), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n915), .A2(KEYINPUT37), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n911), .A2(new_n909), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n410), .B(new_n409), .C1(new_n462), .C2(new_n463), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n916), .A2(KEYINPUT109), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n915), .A2(KEYINPUT37), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT109), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n912), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT38), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT40), .B1(new_n914), .B2(new_n923), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n765), .B(new_n761), .C1(new_n647), .C2(new_n695), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT105), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n421), .A2(new_n695), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n926), .B1(new_n457), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n927), .ZN(new_n929));
  NOR4_X1   g0729(.A1(new_n653), .A2(new_n446), .A3(KEYINPUT105), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n456), .A2(new_n421), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n928), .A2(new_n930), .B1(new_n931), .B2(new_n696), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n925), .A2(new_n932), .A3(new_n883), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n924), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT110), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT40), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT38), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n916), .B1(KEYINPUT37), .B2(new_n904), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n900), .B1(new_n412), .B2(new_n464), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n902), .A2(new_n913), .A3(KEYINPUT38), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n936), .B(new_n937), .C1(new_n943), .C2(new_n933), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n931), .A2(new_n696), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n931), .A2(new_n654), .A3(new_n927), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT105), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n457), .A2(new_n926), .A3(new_n927), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n876), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n941), .A2(new_n942), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n951), .A2(new_n952), .A3(new_n925), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n936), .B1(new_n953), .B2(new_n937), .ZN(new_n954));
  OAI211_X1 g0754(.A(G330), .B(new_n935), .C1(new_n945), .C2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n925), .A2(G330), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n466), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n937), .B1(new_n943), .B2(new_n933), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT110), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n934), .B1(new_n961), .B2(new_n944), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n962), .A2(new_n466), .A3(new_n925), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n749), .A2(new_n466), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n659), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n464), .A2(new_n898), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n950), .B1(new_n882), .B2(new_n875), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n967), .B1(new_n968), .B2(new_n952), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT39), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n914), .B2(new_n923), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n931), .A2(new_n695), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n941), .A2(KEYINPUT39), .A3(new_n942), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n969), .A2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n966), .B(new_n975), .Z(new_n976));
  XNOR2_X1  g0776(.A(new_n964), .B(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n261), .B2(new_n837), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n219), .B1(new_n616), .B2(KEYINPUT35), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n979), .B(new_n229), .C1(KEYINPUT35), .C2(new_n616), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT36), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n233), .A2(G77), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n373), .A2(new_n375), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n982), .A2(new_n983), .B1(G50), .B2(new_n217), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n984), .A2(G1), .A3(new_n685), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n978), .A2(new_n981), .A3(new_n985), .ZN(G367));
  OAI22_X1  g0786(.A1(new_n814), .A2(new_n222), .B1(new_n788), .B2(new_n230), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n857), .A2(new_n217), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(new_n806), .B2(G150), .ZN(new_n989));
  INV_X1    g0789(.A(G137), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n989), .B1(new_n990), .B2(new_n777), .C1(new_n792), .C2(new_n339), .ZN(new_n991));
  NOR3_X1   g0791(.A1(new_n987), .A2(new_n991), .A3(new_n322), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n795), .A2(G143), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(new_n818), .C2(new_n783), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n322), .B1(new_n783), .B2(new_n864), .ZN(new_n995));
  OAI21_X1  g0795(.A(KEYINPUT46), .B1(new_n789), .B2(new_n219), .ZN(new_n996));
  OR3_X1    g0796(.A1(new_n788), .A2(KEYINPUT46), .A3(new_n219), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n210), .B2(new_n792), .C1(new_n328), .C2(new_n857), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n995), .B(new_n999), .C1(G283), .C2(new_n848), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(KEYINPUT113), .B(G317), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n778), .A2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1000), .B(new_n1002), .C1(new_n802), .C2(new_n809), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n816), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1004), .A2(new_n790), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n994), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT47), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n775), .ZN(new_n1008));
  OR3_X1    g0808(.A1(new_n679), .A2(new_n541), .A3(new_n696), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n542), .B1(new_n541), .B2(new_n696), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n834), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n826), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n835), .B1(new_n204), .B2(new_n347), .C1(new_n241), .C2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1008), .A2(new_n838), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n261), .B1(new_n837), .B2(G45), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n667), .A2(new_n696), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n635), .A2(new_n630), .A3(new_n695), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1019), .B1(new_n638), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n715), .A2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT44), .Z(new_n1023));
  NOR2_X1   g0823(.A1(new_n715), .A2(new_n1021), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT45), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(new_n712), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n702), .A2(KEYINPUT112), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n710), .B(new_n713), .Z(new_n1029));
  XNOR2_X1  g0829(.A(new_n1028), .B(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n769), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1027), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n769), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n718), .B(KEYINPUT41), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1018), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n714), .A2(new_n1021), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT42), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n645), .B1(new_n1021), .B2(new_n599), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n696), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1011), .B(KEYINPUT111), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT43), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1041), .B(new_n1044), .C1(new_n1043), .C2(new_n1012), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n1044), .B2(new_n1041), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n711), .A2(new_n1021), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1046), .B(new_n1047), .Z(new_n1048));
  OAI21_X1  g0848(.A(new_n1016), .B1(new_n1036), .B2(new_n1048), .ZN(G387));
  INV_X1    g0849(.A(new_n788), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(G77), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n217), .B2(new_n803), .C1(new_n818), .C2(new_n809), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G50), .B2(new_n806), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n798), .A2(new_n346), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n778), .A2(G150), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(new_n783), .C2(new_n256), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n862), .B2(G97), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1053), .A2(new_n277), .A3(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n848), .A2(G303), .B1(G322), .B2(new_n795), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n802), .B2(new_n783), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n816), .B2(new_n1001), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT48), .Z(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n793), .B2(new_n857), .C1(new_n864), .C2(new_n788), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT49), .Z(new_n1064));
  AOI21_X1  g0864(.A(new_n277), .B1(new_n778), .B2(G326), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n792), .B2(new_n219), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1058), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n775), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n834), .B1(new_n708), .B2(new_n709), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n721), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1070), .B(new_n288), .C1(new_n217), .C2(new_n339), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT115), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n255), .A2(new_n222), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT50), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n826), .B1(new_n288), .B2(new_n238), .C1(new_n1072), .C2(new_n1074), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(G107), .B2(new_n204), .C1(new_n1070), .C2(new_n829), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n835), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1068), .A2(new_n838), .A3(new_n1069), .A4(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1030), .A2(new_n1017), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT114), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1032), .A2(new_n718), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1078), .B(new_n1080), .C1(new_n1081), .C2(new_n1082), .ZN(G393));
  AOI21_X1  g0883(.A(new_n719), .B1(new_n1027), .B2(new_n1032), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1033), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n277), .B1(new_n778), .B2(G322), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1086), .B1(new_n788), .B2(new_n793), .C1(new_n550), .C2(new_n792), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT116), .Z(new_n1088));
  AOI22_X1  g0888(.A1(new_n795), .A2(G317), .B1(new_n806), .B2(G311), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT52), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G116), .B2(new_n798), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1088), .B(new_n1091), .C1(new_n864), .C2(new_n803), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G303), .B2(new_n782), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n795), .A2(G150), .B1(new_n806), .B2(G159), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT51), .Z(new_n1095));
  OAI211_X1 g0895(.A(new_n1095), .B(new_n863), .C1(new_n217), .C2(new_n788), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n857), .A2(new_n339), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n778), .A2(G143), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n277), .B1(new_n222), .B2(new_n783), .C1(new_n814), .C2(new_n345), .ZN(new_n1099));
  NOR4_X1   g0899(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n775), .B1(new_n1093), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1021), .A2(new_n834), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n835), .B1(new_n210), .B2(new_n204), .C1(new_n246), .C2(new_n1014), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1101), .A2(new_n838), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n1027), .B2(new_n1017), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1085), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(G390));
  NAND2_X1  g0907(.A1(new_n1050), .A2(G150), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT53), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n277), .B1(new_n792), .B2(new_n222), .ZN(new_n1110));
  XOR2_X1   g0910(.A(KEYINPUT54), .B(G143), .Z(new_n1111));
  NAND2_X1  g0911(.A1(new_n848), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(G128), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1112), .B1(new_n1113), .B2(new_n809), .C1(new_n990), .C2(new_n783), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1110), .B(new_n1114), .C1(G159), .C2(new_n798), .ZN(new_n1115));
  INV_X1    g0915(.A(G125), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n777), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1109), .B(new_n1117), .C1(G132), .C2(new_n806), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n862), .A2(G68), .B1(G294), .B2(new_n778), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1119), .A2(new_n1120), .B1(G283), .B2(new_n795), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1121), .B1(new_n210), .B2(new_n814), .C1(new_n219), .C2(new_n805), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n783), .A2(new_n328), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n322), .B1(new_n339), .B2(new_n857), .C1(new_n789), .C2(new_n208), .ZN(new_n1125));
  NOR4_X1   g0925(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n775), .B1(new_n1118), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n971), .A2(new_n973), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n832), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1127), .A2(new_n838), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n256), .B2(new_n878), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n941), .A2(KEYINPUT39), .A3(new_n942), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n912), .A2(new_n920), .A3(new_n921), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n918), .A2(new_n917), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n912), .B2(new_n921), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n938), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT39), .B1(new_n1136), .B2(new_n942), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1132), .A2(new_n1137), .B1(new_n968), .B2(new_n972), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n768), .A2(new_n883), .A3(new_n932), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n353), .B1(new_n870), .B2(new_n871), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n695), .B(new_n1140), .C1(new_n746), .C2(new_n747), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n932), .B1(new_n1141), .B2(new_n874), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n972), .B1(new_n1136), .B2(new_n942), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AND4_X1   g0944(.A1(KEYINPUT117), .A2(new_n1138), .A3(new_n1139), .A4(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n972), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n874), .B1(new_n740), .B2(new_n362), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1146), .B1(new_n1147), .B2(new_n950), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1148), .A2(new_n1128), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n957), .A2(new_n951), .ZN(new_n1150));
  OAI21_X1  g0950(.A(KEYINPUT117), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1138), .A2(new_n1139), .A3(new_n1144), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1145), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1131), .B1(new_n1153), .B2(new_n1018), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT120), .Z(new_n1155));
  AOI21_X1  g0955(.A(new_n1150), .B1(new_n1138), .B2(new_n1144), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT117), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1152), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n965), .A2(new_n958), .A3(new_n659), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1147), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n932), .B1(new_n768), .B2(new_n883), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n956), .A2(new_n876), .A3(new_n950), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1141), .A2(new_n874), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n950), .B1(new_n956), .B2(new_n876), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1139), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1159), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1149), .A2(KEYINPUT117), .A3(new_n1139), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1158), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT118), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1153), .A2(KEYINPUT118), .A3(new_n1167), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1173), .B(new_n718), .C1(new_n1167), .C2(new_n1153), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1155), .A2(new_n1174), .ZN(G378));
  XNOR2_X1  g0975(.A(new_n1159), .B(KEYINPUT122), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT118), .B1(new_n1153), .B2(new_n1167), .ZN(new_n1177));
  AND4_X1   g0977(.A1(KEYINPUT118), .A2(new_n1158), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1176), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n975), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n311), .A2(new_n364), .ZN(new_n1181));
  XOR2_X1   g0981(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1182));
  XOR2_X1   g0982(.A(new_n1181), .B(new_n1182), .Z(new_n1183));
  NAND2_X1  g0983(.A1(new_n267), .A2(new_n898), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1183), .B(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n955), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1184), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1183), .B(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n962), .B2(G330), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1180), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n955), .A2(new_n1185), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n962), .A2(G330), .A3(new_n1188), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1191), .A2(new_n1192), .A3(new_n975), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1190), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1179), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT57), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n719), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT123), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1198), .B(new_n1180), .C1(new_n1186), .C2(new_n1189), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1190), .A2(KEYINPUT123), .A3(new_n1193), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1179), .A2(KEYINPUT57), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(KEYINPUT124), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1196), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT124), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1203), .A2(new_n1204), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1197), .A2(new_n1202), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1194), .A2(new_n1018), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n862), .A2(G58), .B1(G107), .B2(new_n806), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n219), .B2(new_n809), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n988), .B(new_n1209), .C1(G283), .C2(new_n778), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n811), .A2(new_n346), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G41), .B(new_n277), .C1(new_n782), .C2(G97), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1210), .A2(new_n1051), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT58), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1050), .A2(new_n1111), .B1(G150), .B2(new_n798), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n782), .A2(G132), .B1(new_n811), .B2(G137), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n1116), .B2(new_n809), .C1(new_n1113), .C2(new_n805), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1219));
  AOI21_X1  g1019(.A(G41), .B1(new_n1218), .B2(KEYINPUT59), .ZN(new_n1220));
  AOI21_X1  g1020(.A(G33), .B1(new_n778), .B2(G124), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(new_n818), .C2(new_n792), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1214), .B1(new_n1219), .B2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(G50), .B1(new_n276), .B2(new_n287), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT121), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n775), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n842), .B1(new_n878), .B2(new_n222), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1226), .B(new_n1227), .C1(new_n1185), .C2(new_n833), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1207), .A2(new_n1228), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1206), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(G375));
  OAI221_X1 g1031(.A(new_n1054), .B1(new_n328), .B2(new_n814), .C1(new_n789), .C2(new_n210), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n322), .B1(new_n792), .B2(new_n339), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT125), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n783), .A2(new_n219), .B1(new_n790), .B2(new_n777), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1232), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n793), .B2(new_n805), .C1(new_n864), .C2(new_n809), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1004), .A2(new_n990), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n859), .A2(G159), .B1(G58), .B2(new_n862), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n811), .A2(G150), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n798), .A2(G50), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n277), .B1(new_n1113), .B2(new_n777), .C1(new_n809), .C2(new_n845), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n782), .B2(new_n1111), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .A4(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1237), .B1(new_n1238), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n775), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1246), .B(new_n838), .C1(new_n833), .C2(new_n932), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n217), .B2(new_n878), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1248), .B1(new_n1250), .B2(new_n1018), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1159), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1035), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1251), .B1(new_n1253), .B2(new_n1167), .ZN(G381));
  AND2_X1   g1054(.A1(new_n1174), .A2(new_n1154), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1230), .A2(new_n1255), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1257));
  XOR2_X1   g1057(.A(new_n1257), .B(KEYINPUT126), .Z(new_n1258));
  OAI211_X1 g1058(.A(new_n1106), .B(new_n1016), .C1(new_n1036), .C2(new_n1048), .ZN(new_n1259));
  OR4_X1    g1059(.A1(G381), .A2(new_n1256), .A3(new_n1258), .A4(new_n1259), .ZN(G407));
  OAI211_X1 g1060(.A(G407), .B(G213), .C1(G343), .C2(new_n1256), .ZN(G409));
  NOR2_X1   g1061(.A1(new_n690), .A2(G343), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1206), .A2(G378), .A3(new_n1229), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1179), .A2(new_n1035), .A3(new_n1194), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1200), .A2(new_n1018), .A3(new_n1199), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1228), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1255), .B1(new_n1264), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1262), .B1(new_n1263), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT60), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n719), .B(new_n1167), .C1(new_n1252), .C2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1249), .A2(KEYINPUT60), .A3(new_n1159), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1251), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(new_n886), .B2(new_n881), .ZN(new_n1274));
  AOI21_X1  g1074(.A(G384), .B1(new_n1272), .B2(new_n1251), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1262), .A2(G2897), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G2897), .B(new_n1262), .C1(new_n1274), .C2(new_n1275), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(KEYINPUT63), .B1(new_n1268), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1268), .A2(new_n1276), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G387), .A2(G390), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1259), .ZN(new_n1285));
  XOR2_X1   g1085(.A(G393), .B(G396), .Z(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(G393), .B(G396), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(new_n1259), .A3(new_n1284), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  XOR2_X1   g1090(.A(new_n1273), .B(G384), .Z(new_n1291));
  AOI211_X1 g1091(.A(new_n1262), .B(new_n1291), .C1(new_n1263), .C2(new_n1267), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1290), .B1(new_n1292), .B2(KEYINPUT63), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT61), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1283), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  XOR2_X1   g1095(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1296));
  AND3_X1   g1096(.A1(new_n1268), .A2(new_n1276), .A3(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1294), .B1(new_n1268), .B2(new_n1280), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1299), .B1(new_n1268), .B2(new_n1276), .ZN(new_n1300));
  NOR3_X1   g1100(.A1(new_n1297), .A2(new_n1298), .A3(new_n1300), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1295), .B1(new_n1301), .B2(new_n1302), .ZN(G405));
  INV_X1    g1103(.A(new_n1263), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1255), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1230), .A2(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1302), .B1(new_n1304), .B2(new_n1306), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1290), .B(new_n1263), .C1(new_n1230), .C2(new_n1305), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1291), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1307), .A2(new_n1308), .A3(new_n1276), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(G402));
endmodule


