//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1255,
    new_n1256, new_n1257, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AND3_X1   g0005(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n206));
  AOI21_X1  g0006(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT65), .ZN(new_n211));
  INV_X1    g0011(.A(new_n201), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G50), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G1), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT0), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G97), .ZN(new_n224));
  INV_X1    g0024(.A(G257), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n217), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n220), .B1(KEYINPUT1), .B2(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n214), .B(new_n231), .C1(KEYINPUT1), .C2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT66), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT67), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G58), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G1), .A3(G13), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G274), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n215), .B1(G41), .B2(G45), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT68), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n215), .B(KEYINPUT68), .C1(G41), .C2(G45), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(new_n251), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n254), .B1(new_n259), .B2(G238), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G33), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n262), .A2(new_n264), .A3(G232), .A4(G1698), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n262), .A2(new_n264), .A3(G226), .A4(new_n266), .ZN(new_n267));
  AND3_X1   g0067(.A1(KEYINPUT73), .A2(G33), .A3(G97), .ZN(new_n268));
  AOI21_X1  g0068(.A(KEYINPUT73), .B1(G33), .B2(G97), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n265), .A2(new_n267), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G1), .A2(G13), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT64), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n276), .A2(new_n250), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT74), .ZN(new_n278));
  AND3_X1   g0078(.A1(new_n271), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n278), .B1(new_n271), .B2(new_n277), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n260), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT13), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT13), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n283), .B(new_n260), .C1(new_n279), .C2(new_n280), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G200), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(G68), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n287), .A2(G50), .B1(G20), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G77), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n209), .A2(G33), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n208), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n295), .A2(KEYINPUT11), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n215), .A2(G13), .A3(G20), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n274), .A2(new_n297), .A3(new_n275), .A4(new_n293), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n215), .A2(G20), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(G68), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n297), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n288), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT12), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n295), .A2(KEYINPUT11), .ZN(new_n305));
  AND4_X1   g0105(.A1(new_n296), .A2(new_n301), .A3(new_n304), .A4(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n282), .A2(G190), .A3(new_n284), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n286), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(KEYINPUT75), .A2(G169), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n285), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT14), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n310), .B1(new_n282), .B2(new_n284), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT14), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n282), .A2(G179), .A3(new_n284), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n313), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n306), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n309), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n294), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT3), .B(G33), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT7), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n322), .A2(new_n323), .A3(G20), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n262), .A2(new_n264), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT7), .B1(new_n325), .B2(new_n209), .ZN(new_n326));
  OAI21_X1  g0126(.A(G68), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n222), .A2(new_n288), .ZN(new_n328));
  OAI21_X1  g0128(.A(G20), .B1(new_n328), .B2(new_n201), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n287), .A2(G159), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT16), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n321), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n327), .A2(KEYINPUT16), .A3(new_n332), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT8), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G58), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n222), .A2(KEYINPUT8), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT69), .ZN(new_n340));
  OR3_X1    g0140(.A1(new_n222), .A2(KEYINPUT69), .A3(KEYINPUT8), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n302), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n298), .B(KEYINPUT70), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n340), .A2(new_n341), .A3(new_n300), .ZN(new_n345));
  OAI211_X1 g0145(.A(KEYINPUT76), .B(new_n343), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT76), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n208), .A2(KEYINPUT70), .A3(new_n293), .A4(new_n297), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT70), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n298), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n345), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n343), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n347), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n335), .A2(new_n336), .B1(new_n346), .B2(new_n353), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n262), .A2(new_n264), .A3(G226), .A4(G1698), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n262), .A2(new_n264), .A3(G223), .A4(new_n266), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G33), .A2(G87), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT77), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT77), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n355), .A2(new_n356), .A3(new_n360), .A4(new_n357), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n277), .A3(new_n361), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n258), .A2(new_n223), .B1(new_n252), .B2(new_n253), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n362), .A2(G190), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G200), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(new_n362), .B2(new_n364), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT79), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n354), .A2(new_n368), .A3(new_n369), .A4(KEYINPUT17), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n369), .A2(KEYINPUT17), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(KEYINPUT17), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n346), .A2(new_n353), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n323), .B1(new_n322), .B2(G20), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n325), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n288), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n334), .B1(new_n376), .B2(new_n331), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n336), .A2(new_n377), .A3(new_n294), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n362), .A2(G190), .A3(new_n364), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n361), .A2(new_n277), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n363), .B1(new_n381), .B2(new_n359), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n380), .B1(new_n382), .B2(new_n366), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n371), .B(new_n372), .C1(new_n379), .C2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n370), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n362), .A2(G179), .A3(new_n364), .ZN(new_n386));
  INV_X1    g0186(.A(G169), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n386), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n379), .A2(KEYINPUT18), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT78), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n379), .A2(new_n388), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT18), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n392), .A2(new_n390), .A3(new_n393), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n385), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT72), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT10), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n398), .A2(KEYINPUT10), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n322), .A2(G222), .A3(new_n266), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n322), .A2(G1698), .ZN(new_n402));
  INV_X1    g0202(.A(G223), .ZN(new_n403));
  OAI221_X1 g0203(.A(new_n401), .B1(new_n290), .B2(new_n322), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n277), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n254), .B1(new_n259), .B2(G226), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G200), .ZN(new_n408));
  INV_X1    g0208(.A(G190), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n408), .B1(new_n409), .B2(new_n407), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n287), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n342), .B2(new_n291), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n412), .A2(new_n294), .B1(new_n202), .B2(new_n302), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n348), .A2(new_n350), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n414), .A2(G50), .A3(new_n300), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT9), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n416), .B1(new_n413), .B2(new_n415), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n399), .B(new_n400), .C1(new_n410), .C2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n287), .ZN(new_n422));
  XNOR2_X1  g0222(.A(KEYINPUT8), .B(G58), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT71), .ZN(new_n424));
  OR2_X1    g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n424), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n422), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g0227(.A(KEYINPUT15), .B(G87), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n428), .A2(new_n291), .B1(new_n209), .B2(new_n290), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n294), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n290), .B1(new_n215), .B2(G20), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n299), .A2(new_n431), .B1(new_n290), .B2(new_n302), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G238), .ZN(new_n434));
  INV_X1    g0234(.A(G107), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n402), .A2(new_n434), .B1(new_n435), .B2(new_n322), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n325), .A2(new_n223), .A3(G1698), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n277), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n254), .B1(new_n259), .B2(G244), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n433), .B1(G190), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n439), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G200), .ZN(new_n443));
  INV_X1    g0243(.A(G179), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n442), .A2(new_n387), .B1(new_n430), .B2(new_n432), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n441), .A2(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n419), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n417), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n366), .B1(new_n405), .B2(new_n406), .ZN(new_n450));
  INV_X1    g0250(.A(new_n407), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(G190), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n449), .A2(new_n452), .A3(new_n398), .A4(KEYINPUT10), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n407), .A2(new_n387), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n413), .A2(new_n415), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n454), .B(new_n455), .C1(G179), .C2(new_n407), .ZN(new_n456));
  AND4_X1   g0256(.A1(new_n421), .A2(new_n447), .A3(new_n453), .A4(new_n456), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n320), .A2(new_n397), .A3(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n262), .A2(new_n264), .A3(G257), .A4(new_n266), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT84), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT84), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n322), .A2(new_n461), .A3(G257), .A4(new_n266), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n325), .A2(G303), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n322), .A2(G264), .A3(G1698), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n460), .A2(new_n462), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n277), .ZN(new_n466));
  INV_X1    g0266(.A(G45), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(G1), .ZN(new_n468));
  AND2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  NOR2_X1   g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(G270), .A3(new_n251), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT5), .B(G41), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n473), .A2(G274), .A3(new_n468), .A4(new_n251), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n466), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT85), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT85), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n466), .A2(new_n479), .A3(new_n476), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(G200), .A3(new_n480), .ZN(new_n481));
  AOI211_X1 g0281(.A(KEYINPUT85), .B(new_n475), .C1(new_n465), .C2(new_n277), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n479), .B1(new_n466), .B2(new_n476), .ZN(new_n483));
  OAI21_X1  g0283(.A(G190), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(G20), .B1(G33), .B2(G283), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n261), .A2(G97), .ZN(new_n486));
  INV_X1    g0286(.A(G116), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n485), .A2(new_n486), .B1(G20), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n294), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT20), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n294), .A2(KEYINPUT20), .A3(new_n488), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n491), .A2(new_n492), .B1(new_n487), .B2(new_n302), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n261), .A2(G1), .ZN(new_n494));
  XNOR2_X1  g0294(.A(new_n494), .B(KEYINPUT81), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n299), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G116), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n481), .A2(new_n484), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT86), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n481), .A2(new_n484), .A3(new_n500), .A4(KEYINPUT86), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n482), .A2(new_n483), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n387), .B1(new_n493), .B2(new_n498), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n506), .A2(KEYINPUT21), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n466), .A2(G179), .A3(new_n476), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n499), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT21), .B1(new_n506), .B2(new_n507), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n505), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n471), .A2(new_n251), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n474), .B1(new_n516), .B2(new_n225), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n262), .A2(new_n264), .A3(G250), .A4(G1698), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT82), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n322), .A2(KEYINPUT82), .A3(G250), .A4(G1698), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n322), .A2(KEYINPUT4), .A3(G244), .A4(new_n266), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n262), .A2(new_n264), .A3(G244), .A4(new_n266), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT4), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n524), .A2(new_n525), .B1(G33), .B2(G283), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n522), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n517), .B1(new_n527), .B2(new_n277), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT83), .B1(new_n528), .B2(new_n366), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT83), .ZN(new_n530));
  INV_X1    g0330(.A(new_n277), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n524), .A2(new_n525), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G283), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n532), .A2(new_n523), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n531), .B1(new_n534), .B2(new_n522), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n530), .B(G200), .C1(new_n535), .C2(new_n517), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n495), .A2(new_n299), .A3(G97), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n297), .A2(G97), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT80), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT6), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n224), .A2(new_n435), .ZN(new_n543));
  NOR2_X1   g0343(.A1(G97), .A2(G107), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n435), .A2(KEYINPUT6), .A3(G97), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n209), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n422), .A2(new_n290), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n541), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(G107), .B1(new_n324), .B2(new_n326), .ZN(new_n550));
  INV_X1    g0350(.A(new_n548), .ZN(new_n551));
  INV_X1    g0351(.A(new_n546), .ZN(new_n552));
  XNOR2_X1  g0352(.A(G97), .B(G107), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n552), .B1(new_n542), .B2(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(KEYINPUT80), .B(new_n551), .C1(new_n554), .C2(new_n209), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n549), .A2(new_n550), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n540), .B1(new_n556), .B2(new_n294), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n528), .A2(G190), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n529), .A2(new_n536), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n556), .A2(new_n294), .ZN(new_n560));
  INV_X1    g0360(.A(new_n540), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n528), .A2(new_n444), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n527), .A2(new_n277), .ZN(new_n564));
  INV_X1    g0364(.A(new_n517), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n387), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n562), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n322), .A2(new_n209), .A3(G68), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n291), .A2(new_n224), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n569), .B1(KEYINPUT19), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT19), .B1(new_n268), .B2(new_n269), .ZN(new_n572));
  INV_X1    g0372(.A(G87), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n572), .A2(new_n209), .B1(new_n573), .B2(new_n544), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n294), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n428), .A2(new_n302), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n575), .B(new_n576), .C1(new_n496), .C2(new_n428), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n251), .A2(G274), .A3(new_n468), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n215), .A2(G45), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n251), .A2(G250), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n262), .A2(new_n264), .A3(G238), .A4(new_n266), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n262), .A2(new_n264), .A3(G244), .A4(G1698), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n582), .B(new_n583), .C1(new_n261), .C2(new_n487), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n581), .B1(new_n584), .B2(new_n277), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n585), .A2(G169), .ZN(new_n586));
  AOI211_X1 g0386(.A(G179), .B(new_n581), .C1(new_n277), .C2(new_n584), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI211_X1 g0388(.A(new_n409), .B(new_n581), .C1(new_n277), .C2(new_n584), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n584), .A2(new_n277), .ZN(new_n590));
  INV_X1    g0390(.A(new_n581), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n366), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n495), .A2(new_n299), .A3(G87), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n575), .A2(new_n594), .A3(new_n576), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n577), .A2(new_n588), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n559), .A2(new_n568), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n322), .A2(G250), .A3(new_n266), .ZN(new_n598));
  NAND2_X1  g0398(.A1(G33), .A2(G294), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n598), .B(new_n599), .C1(new_n402), .C2(new_n225), .ZN(new_n600));
  INV_X1    g0400(.A(new_n516), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n600), .A2(new_n277), .B1(G264), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n474), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n387), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(new_n444), .A3(new_n474), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n322), .A2(new_n209), .A3(G87), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT22), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT22), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n322), .A2(new_n608), .A3(new_n209), .A4(G87), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT23), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n611), .A2(new_n435), .A3(G20), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT87), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n611), .B2(new_n435), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n615));
  OAI22_X1  g0415(.A1(new_n612), .A2(KEYINPUT87), .B1(new_n615), .B2(G20), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n610), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT24), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT24), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n610), .A2(new_n620), .A3(new_n617), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n321), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT25), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n297), .B2(G107), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n302), .A2(KEYINPUT25), .A3(new_n435), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n497), .A2(G107), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n604), .B(new_n605), .C1(new_n622), .C2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n621), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n620), .B1(new_n610), .B2(new_n617), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n294), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n603), .A2(G200), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n602), .A2(G190), .A3(new_n474), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n631), .A2(new_n632), .A3(new_n626), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n628), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n597), .A2(new_n635), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n458), .A2(new_n515), .A3(new_n636), .ZN(G372));
  AND2_X1   g0437(.A1(new_n421), .A2(new_n453), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n317), .B1(new_n314), .B2(new_n315), .ZN(new_n639));
  AOI211_X1 g0439(.A(KEYINPUT14), .B(new_n310), .C1(new_n282), .C2(new_n284), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n319), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n446), .A2(new_n445), .ZN(new_n642));
  AOI211_X1 g0442(.A(new_n385), .B(new_n309), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n394), .A2(new_n389), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n638), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n645), .A2(new_n456), .ZN(new_n646));
  INV_X1    g0446(.A(new_n458), .ZN(new_n647));
  INV_X1    g0447(.A(new_n634), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n597), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n513), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n650), .A2(new_n511), .A3(new_n508), .A4(new_n628), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n562), .A2(new_n563), .A3(new_n567), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n653), .A2(KEYINPUT26), .A3(new_n596), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n593), .A2(new_n595), .ZN(new_n656));
  INV_X1    g0456(.A(new_n587), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n585), .A2(G169), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n577), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n655), .B1(new_n568), .B2(new_n660), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n654), .A2(new_n661), .B1(new_n577), .B2(new_n588), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n652), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n646), .B1(new_n647), .B2(new_n663), .ZN(G369));
  INV_X1    g0464(.A(new_n514), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n215), .A2(new_n209), .A3(G13), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n500), .A2(new_n672), .ZN(new_n673));
  MUX2_X1   g0473(.A(new_n515), .B(new_n665), .S(new_n673), .Z(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n628), .A2(new_n671), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n671), .B1(new_n622), .B2(new_n627), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n634), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n677), .B1(new_n628), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n514), .A2(new_n671), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n677), .B1(new_n682), .B2(new_n680), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(G399));
  INV_X1    g0484(.A(new_n218), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G41), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n544), .A2(new_n573), .A3(new_n487), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT88), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n686), .A2(new_n215), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n213), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n689), .B1(new_n690), .B2(new_n686), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT28), .Z(new_n692));
  AOI211_X1 g0492(.A(KEYINPUT29), .B(new_n671), .C1(new_n652), .C2(new_n662), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT91), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n652), .B1(new_n662), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(KEYINPUT26), .B1(new_n653), .B2(new_n596), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n568), .A2(new_n660), .A3(new_n655), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n659), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(KEYINPUT91), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n672), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n693), .B1(new_n700), .B2(KEYINPUT29), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT31), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n564), .A2(new_n565), .A3(new_n602), .A4(new_n585), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n703), .B1(new_n704), .B2(new_n509), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n602), .A2(new_n585), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n510), .A2(new_n706), .A3(KEYINPUT30), .A4(new_n528), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n566), .A2(new_n603), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n585), .A2(G179), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n478), .A2(new_n480), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n709), .B1(new_n711), .B2(KEYINPUT89), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT89), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n506), .A2(new_n713), .A3(new_n710), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n708), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n702), .B1(new_n715), .B2(new_n672), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT90), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n712), .A2(new_n714), .ZN(new_n719));
  OAI211_X1 g0519(.A(KEYINPUT31), .B(new_n671), .C1(new_n719), .C2(new_n708), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n636), .A2(new_n505), .A3(new_n514), .A4(new_n672), .ZN(new_n721));
  OAI211_X1 g0521(.A(KEYINPUT90), .B(new_n702), .C1(new_n715), .C2(new_n672), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n718), .A2(new_n720), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G330), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n701), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n692), .B1(new_n725), .B2(G1), .ZN(G364));
  INV_X1    g0526(.A(G13), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n727), .A2(new_n467), .A3(G20), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n728), .A2(KEYINPUT92), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(KEYINPUT92), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n729), .A2(G1), .A3(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n686), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g0532(.A(new_n732), .B(KEYINPUT93), .Z(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n208), .B1(G20), .B2(new_n387), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n209), .A2(G190), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G179), .A2(G200), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G159), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT32), .ZN(new_n742));
  NAND3_X1  g0542(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G190), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n743), .A2(new_n409), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n745), .A2(new_n288), .B1(new_n747), .B2(new_n202), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n209), .B1(new_n738), .B2(G190), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n224), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n366), .A2(G179), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n737), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n209), .A2(new_n409), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n751), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n322), .B1(new_n752), .B2(new_n435), .C1(new_n573), .C2(new_n754), .ZN(new_n755));
  NOR4_X1   g0555(.A1(new_n742), .A2(new_n748), .A3(new_n750), .A4(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n444), .A2(G200), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT96), .ZN(new_n758));
  AND3_X1   g0558(.A1(new_n757), .A2(new_n737), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n758), .B1(new_n757), .B2(new_n737), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n753), .A2(new_n757), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n761), .A2(new_n290), .B1(new_n222), .B2(new_n762), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n763), .A2(KEYINPUT97), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(KEYINPUT97), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n756), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G283), .ZN(new_n767));
  INV_X1    g0567(.A(G329), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n752), .A2(new_n767), .B1(new_n739), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G294), .ZN(new_n770));
  INV_X1    g0570(.A(G303), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n325), .B1(new_n749), .B2(new_n770), .C1(new_n771), .C2(new_n754), .ZN(new_n772));
  INV_X1    g0572(.A(new_n762), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n769), .B(new_n772), .C1(G322), .C2(new_n773), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n746), .B(KEYINPUT98), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G326), .ZN(new_n777));
  INV_X1    g0577(.A(new_n761), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G311), .ZN(new_n779));
  XNOR2_X1  g0579(.A(KEYINPUT33), .B(G317), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT99), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n745), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(new_n781), .B2(new_n780), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n774), .A2(new_n777), .A3(new_n779), .A4(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n736), .B1(new_n766), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G13), .A2(G33), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(G20), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n736), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT94), .Z(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT95), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n218), .A2(G355), .A3(new_n322), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n685), .A2(new_n322), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(G45), .B2(new_n213), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n248), .A2(new_n467), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n793), .B1(G116), .B2(new_n218), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n734), .B(new_n785), .C1(new_n792), .C2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT100), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n674), .B2(new_n789), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n675), .B1(new_n686), .B2(new_n731), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n674), .A2(G330), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT101), .Z(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  AOI21_X1  g0605(.A(new_n671), .B1(new_n652), .B2(new_n662), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n642), .B(KEYINPUT103), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n441), .A2(new_n443), .B1(new_n433), .B2(new_n671), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT104), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n642), .B2(new_n672), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n446), .A2(new_n445), .A3(KEYINPUT104), .A4(new_n671), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n807), .A2(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n806), .B(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n732), .B1(new_n814), .B2(new_n724), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n724), .B2(new_n814), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n736), .A2(new_n787), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n733), .B1(G77), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n745), .A2(KEYINPUT102), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n745), .A2(KEYINPUT102), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(G283), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n325), .B1(new_n754), .B2(new_n435), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n750), .B(new_n824), .C1(G303), .C2(new_n746), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n778), .A2(G116), .ZN(new_n826));
  INV_X1    g0626(.A(G311), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n762), .A2(new_n770), .B1(new_n739), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n752), .A2(new_n573), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n823), .A2(new_n825), .A3(new_n826), .A4(new_n830), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n773), .A2(G143), .B1(G137), .B2(new_n746), .ZN(new_n832));
  INV_X1    g0632(.A(G150), .ZN(new_n833));
  INV_X1    g0633(.A(G159), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n832), .B1(new_n833), .B2(new_n745), .C1(new_n834), .C2(new_n761), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT34), .Z(new_n836));
  INV_X1    g0636(.A(new_n752), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n837), .A2(G68), .B1(new_n740), .B2(G132), .ZN(new_n838));
  INV_X1    g0638(.A(new_n754), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n325), .B1(new_n839), .B2(G50), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n838), .B(new_n840), .C1(new_n222), .C2(new_n749), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n831), .B1(new_n836), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n818), .B1(new_n842), .B2(new_n735), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n813), .B2(new_n787), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n816), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(G384));
  INV_X1    g0646(.A(KEYINPUT35), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n487), .B1(new_n554), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n847), .B2(new_n554), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n849), .A2(new_n211), .ZN(new_n850));
  XNOR2_X1  g0650(.A(KEYINPUT105), .B(KEYINPUT36), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n850), .B(new_n851), .ZN(new_n852));
  OR3_X1    g0652(.A1(new_n213), .A2(new_n290), .A3(new_n328), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n202), .A2(G68), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n215), .B(G13), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(G330), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n354), .A2(new_n368), .ZN(new_n858));
  INV_X1    g0658(.A(new_n669), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n379), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT107), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n858), .B(new_n860), .C1(new_n392), .C2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n362), .A2(new_n364), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(G169), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n865), .A2(new_n386), .B1(new_n373), .B2(new_n378), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n863), .B1(new_n866), .B2(KEYINPUT107), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n351), .A2(new_n352), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n378), .A2(new_n870), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n354), .A2(new_n368), .B1(new_n859), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n388), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n863), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n869), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT106), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n871), .A2(new_n859), .ZN(new_n878));
  NOR3_X1   g0678(.A1(new_n397), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n370), .A2(new_n384), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT18), .B1(new_n379), .B2(new_n388), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(new_n390), .B2(new_n389), .ZN(new_n882));
  INV_X1    g0682(.A(new_n396), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n878), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT106), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n876), .B1(new_n879), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT38), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n877), .B1(new_n397), .B2(new_n878), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n884), .A2(KEYINPUT106), .A3(new_n885), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT38), .B1(new_n868), .B2(new_n874), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT108), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT108), .ZN(new_n896));
  AOI211_X1 g0696(.A(new_n896), .B(new_n893), .C1(new_n890), .C2(new_n891), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n889), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n319), .B(new_n671), .C1(new_n318), .C2(new_n309), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n306), .A2(new_n672), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n641), .A2(new_n308), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n812), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n721), .A2(new_n720), .A3(new_n716), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT40), .B1(new_n898), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT109), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n379), .B(new_n859), .C1(new_n644), .C2(new_n385), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n858), .A2(new_n392), .A3(new_n860), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n910), .A2(new_n863), .B1(new_n862), .B2(new_n867), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n892), .B2(new_n894), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n903), .A2(new_n904), .A3(KEYINPUT40), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n908), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n903), .A2(new_n904), .A3(KEYINPUT40), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n893), .B1(new_n890), .B2(new_n891), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n916), .B(KEYINPUT109), .C1(new_n917), .C2(new_n912), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n907), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n458), .A2(new_n904), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n857), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n919), .B2(new_n920), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n807), .A2(new_n671), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n806), .B2(new_n813), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n899), .A2(new_n902), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n898), .A2(new_n927), .B1(new_n644), .B2(new_n669), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n917), .A2(KEYINPUT39), .A3(new_n912), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n898), .B2(KEYINPUT39), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n318), .A2(new_n319), .A3(new_n672), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n646), .B1(new_n701), .B2(new_n647), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n932), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n922), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(G1), .B1(new_n727), .B2(G20), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n922), .A2(new_n934), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n856), .B1(new_n937), .B2(new_n938), .ZN(G367));
  INV_X1    g0739(.A(new_n791), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n218), .B2(new_n428), .ZN(new_n941));
  INV_X1    g0741(.A(new_n794), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n236), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n733), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(G137), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n752), .A2(new_n290), .B1(new_n739), .B2(new_n945), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n322), .B1(new_n749), .B2(new_n288), .C1(new_n762), .C2(new_n833), .ZN(new_n947));
  AOI211_X1 g0747(.A(new_n946), .B(new_n947), .C1(G58), .C2(new_n839), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n202), .B2(new_n761), .ZN(new_n949));
  INV_X1    g0749(.A(G143), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n821), .A2(new_n834), .B1(new_n950), .B2(new_n775), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n839), .A2(G116), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT46), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n952), .A2(new_n953), .B1(new_n435), .B2(new_n749), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n953), .B2(new_n952), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n778), .A2(G283), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n322), .B1(new_n773), .B2(G303), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n837), .A2(G97), .B1(new_n740), .B2(G317), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n955), .A2(new_n956), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n821), .A2(new_n770), .B1(new_n827), .B2(new_n775), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n949), .A2(new_n951), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT47), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n944), .B1(new_n962), .B2(new_n735), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n595), .A2(new_n672), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n964), .A2(new_n577), .A3(new_n588), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n660), .B2(new_n964), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n963), .B1(new_n789), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n653), .A2(new_n671), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT110), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n559), .B(new_n568), .C1(new_n557), .C2(new_n672), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(new_n680), .A3(new_n682), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT42), .Z(new_n974));
  NOR2_X1   g0774(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n568), .B1(new_n971), .B2(new_n628), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n672), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n974), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n978), .A2(KEYINPUT111), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n974), .A2(new_n977), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n966), .B(KEYINPUT43), .Z(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n978), .A2(KEYINPUT111), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n979), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n681), .A2(new_n971), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n984), .B(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n683), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n971), .A2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT44), .Z(new_n990));
  NOR2_X1   g0790(.A1(new_n971), .A2(new_n988), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n993), .A2(new_n676), .A3(new_n680), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n990), .A2(new_n681), .A3(new_n992), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n682), .B(new_n680), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n675), .B(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n725), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n725), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n686), .B(KEYINPUT41), .Z(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n731), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n967), .B1(new_n987), .B2(new_n1007), .ZN(G387));
  NOR2_X1   g0808(.A1(new_n680), .A2(new_n789), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n688), .ZN(new_n1010));
  AOI21_X1  g0810(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n425), .A2(new_n426), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n202), .ZN(new_n1013));
  XOR2_X1   g0813(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n1014));
  OAI211_X1 g0814(.A(new_n1010), .B(new_n1011), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n794), .B1(new_n240), .B2(new_n467), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n688), .A2(new_n218), .A3(new_n322), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(G107), .C2(new_n218), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n792), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n733), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n749), .A2(new_n428), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n322), .B1(new_n752), .B2(new_n224), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(G159), .C2(new_n746), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n342), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n744), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n778), .A2(G68), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n202), .A2(new_n762), .B1(new_n754), .B2(new_n290), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G150), .B2(new_n740), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n322), .B1(new_n740), .B2(G326), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n754), .A2(new_n770), .B1(new_n749), .B2(new_n767), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n778), .A2(G303), .B1(G317), .B2(new_n773), .ZN(new_n1033));
  INV_X1    g0833(.A(G322), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1033), .B1(new_n1034), .B2(new_n775), .C1(new_n821), .C2(new_n827), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT48), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1032), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n1036), .B2(new_n1035), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT49), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1031), .B1(new_n487), .B2(new_n752), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1030), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1009), .B(new_n1021), .C1(new_n1042), .C2(new_n735), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n1000), .B2(new_n731), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1001), .A2(new_n686), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1000), .A2(new_n725), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(G393));
  INV_X1    g0847(.A(new_n686), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n997), .B2(new_n1002), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n996), .A2(new_n1001), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n940), .B1(new_n224), .B2(new_n218), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n245), .A2(new_n942), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n733), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n749), .A2(new_n487), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G283), .A2(new_n839), .B1(new_n740), .B2(G322), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1056), .B(new_n325), .C1(new_n435), .C2(new_n752), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1055), .B(new_n1057), .C1(G294), .C2(new_n778), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n773), .A2(G311), .B1(G317), .B2(new_n746), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT52), .Z(new_n1060));
  OAI211_X1 g0860(.A(new_n1058), .B(new_n1060), .C1(new_n771), .C2(new_n821), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1061), .A2(KEYINPUT113), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n822), .A2(G50), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n747), .A2(new_n833), .B1(new_n762), .B2(new_n834), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT51), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n778), .A2(new_n1012), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n754), .A2(new_n288), .B1(new_n739), .B2(new_n950), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n749), .A2(new_n290), .ZN(new_n1068));
  NOR4_X1   g0868(.A1(new_n1067), .A2(new_n829), .A3(new_n1068), .A4(new_n325), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1063), .A2(new_n1065), .A3(new_n1066), .A4(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1061), .A2(KEYINPUT113), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1062), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1054), .B1(new_n1072), .B2(new_n735), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n972), .B2(new_n789), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n731), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1074), .B1(new_n996), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1051), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(G390));
  INV_X1    g0878(.A(new_n929), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n931), .B1(new_n924), .B2(new_n926), .ZN(new_n1080));
  AOI21_X1  g0880(.A(KEYINPUT38), .B1(new_n892), .B2(new_n876), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n894), .B1(new_n879), .B2(new_n886), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n896), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n917), .A2(KEYINPUT108), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1081), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT39), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1079), .B(new_n1080), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n723), .A2(G330), .A3(new_n813), .A4(new_n925), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n912), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1082), .A2(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n931), .B(KEYINPUT114), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n698), .A2(KEYINPUT91), .B1(new_n649), .B2(new_n651), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n662), .A2(new_n694), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n671), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n923), .B1(new_n1094), .B2(new_n813), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1090), .B(new_n1091), .C1(new_n1095), .C2(new_n926), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1087), .A2(new_n1088), .A3(new_n1096), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n1087), .A2(new_n1096), .ZN(new_n1098));
  AND4_X1   g0898(.A1(G330), .A2(new_n904), .A3(new_n813), .A4(new_n925), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n731), .B(new_n1097), .C1(new_n1098), .C2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n733), .B1(new_n1025), .B2(new_n817), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n749), .A2(new_n834), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n839), .A2(G150), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT53), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1103), .B(new_n1105), .C1(G128), .C2(new_n746), .ZN(new_n1106));
  INV_X1    g0906(.A(G132), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n762), .A2(new_n1107), .B1(new_n752), .B2(new_n202), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n325), .B(new_n1108), .C1(G125), .C2(new_n740), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(KEYINPUT54), .B(G143), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1106), .B(new_n1109), .C1(new_n761), .C2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n821), .A2(new_n945), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n821), .A2(new_n435), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n325), .B1(new_n754), .B2(new_n573), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1068), .B(new_n1114), .C1(G283), .C2(new_n746), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n762), .A2(new_n487), .B1(new_n752), .B2(new_n288), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(G294), .B2(new_n740), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1115), .B(new_n1117), .C1(new_n224), .C2(new_n761), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1111), .A2(new_n1112), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1102), .B1(new_n1119), .B2(new_n735), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1079), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1120), .B1(new_n1121), .B2(new_n787), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1101), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT117), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1101), .A2(KEYINPUT117), .A3(new_n1122), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1097), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n458), .A2(new_n904), .A3(G330), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT115), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1129), .B(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(KEYINPUT116), .B1(new_n933), .B2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1129), .B(KEYINPUT115), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n693), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT29), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1134), .B1(new_n1094), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n458), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT116), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1133), .A2(new_n1137), .A3(new_n1138), .A4(new_n646), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n904), .A2(G330), .A3(new_n813), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n926), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1095), .A2(new_n1088), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n723), .A2(G330), .A3(new_n813), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1099), .B1(new_n926), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1142), .B1(new_n1144), .B2(new_n924), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1132), .A2(new_n1139), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1048), .B1(new_n1128), .B2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1146), .B(new_n1097), .C1(new_n1098), .C2(new_n1100), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1127), .A2(new_n1150), .ZN(G378));
  INV_X1    g0951(.A(KEYINPUT40), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n1085), .B2(new_n905), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n857), .B1(new_n915), .B2(new_n918), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n638), .A2(new_n456), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n455), .A2(new_n859), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1155), .B(new_n1156), .Z(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1157), .B(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1153), .A2(new_n1154), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1160), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(new_n1161), .A2(new_n1162), .A3(new_n932), .ZN(new_n1163));
  AOI21_X1  g0963(.A(KEYINPUT109), .B1(new_n1090), .B2(new_n916), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n913), .A2(new_n908), .A3(new_n914), .ZN(new_n1165));
  OAI21_X1  g0965(.A(G330), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1159), .B1(new_n1166), .B2(new_n907), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1153), .A2(new_n1154), .A3(new_n1160), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n931), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1121), .A2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1167), .A2(new_n1168), .B1(new_n1170), .B2(new_n928), .ZN(new_n1171));
  OAI21_X1  g0971(.A(KEYINPUT57), .B1(new_n1163), .B2(new_n1171), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1132), .A2(new_n1139), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1087), .A2(new_n1088), .A3(new_n1096), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1100), .B1(new_n1087), .B2(new_n1096), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1174), .B1(new_n1177), .B2(new_n1146), .ZN(new_n1178));
  OAI21_X1  g0978(.A(KEYINPUT121), .B1(new_n1172), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1149), .A2(new_n1173), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT121), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n932), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1167), .A2(new_n1170), .A3(new_n928), .A4(new_n1168), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1180), .A2(new_n1181), .A3(new_n1184), .A4(KEYINPUT57), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1179), .A2(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1149), .A2(new_n1173), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n686), .B1(new_n1187), .B2(KEYINPUT57), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n322), .A2(G41), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G77), .B2(new_n839), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(new_n222), .B2(new_n752), .C1(new_n767), .C2(new_n739), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT118), .Z(new_n1193));
  OAI22_X1  g0993(.A1(new_n745), .A2(new_n224), .B1(new_n747), .B2(new_n487), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n762), .A2(new_n435), .B1(new_n749), .B2(new_n288), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1193), .B(new_n1196), .C1(new_n428), .C2(new_n761), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT119), .Z(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT120), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1199), .A2(KEYINPUT58), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(KEYINPUT58), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1190), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1202));
  AOI211_X1 g1002(.A(G33), .B(G41), .C1(new_n740), .C2(G124), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n746), .A2(G125), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n833), .B2(new_n749), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n773), .A2(G128), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n754), .B2(new_n1110), .C1(new_n745), .C2(new_n1107), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1205), .B(new_n1207), .C1(G137), .C2(new_n778), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT59), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1203), .B1(new_n834), .B2(new_n752), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1202), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1200), .A2(new_n1201), .A3(new_n1212), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n732), .B1(G50), .B2(new_n817), .C1(new_n1213), .C2(new_n736), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n786), .B2(new_n1159), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n1184), .B2(new_n731), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1189), .A2(new_n1216), .ZN(G375));
  INV_X1    g1017(.A(new_n1145), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1174), .A2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1219), .A2(new_n1006), .A3(new_n1147), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT122), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1145), .A2(new_n1221), .A3(new_n731), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n821), .A2(new_n487), .B1(new_n435), .B2(new_n761), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT124), .Z(new_n1225));
  OAI22_X1  g1025(.A1(new_n224), .A2(new_n754), .B1(new_n762), .B2(new_n767), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G303), .B2(new_n740), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1022), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n746), .A2(G294), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n322), .B1(new_n837), .B2(G77), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1225), .A2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n325), .B1(new_n837), .B2(G58), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n202), .B2(new_n749), .C1(new_n747), .C2(new_n1107), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n821), .A2(new_n1110), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G137), .A2(new_n773), .B1(new_n740), .B2(G128), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n834), .B2(new_n754), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n761), .A2(new_n833), .ZN(new_n1238));
  NOR4_X1   g1038(.A1(new_n1234), .A2(new_n1235), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n735), .B1(new_n1232), .B2(new_n1239), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1240), .B(new_n733), .C1(G68), .C2(new_n817), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(KEYINPUT125), .Z(new_n1242));
  NAND2_X1  g1042(.A1(new_n926), .A2(new_n786), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1242), .B1(new_n1243), .B2(KEYINPUT123), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(KEYINPUT123), .B2(new_n1243), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1221), .B1(new_n1145), .B2(new_n731), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1223), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1220), .A2(new_n1247), .ZN(G381));
  OAI211_X1 g1048(.A(new_n1077), .B(new_n967), .C1(new_n1007), .C2(new_n987), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT126), .Z(new_n1251));
  NOR3_X1   g1051(.A1(new_n1249), .A2(G381), .A3(new_n1251), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1125), .A2(new_n1126), .B1(new_n1149), .B2(new_n1148), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1252), .A2(new_n1253), .A3(new_n1216), .A4(new_n1189), .ZN(G407));
  NAND2_X1  g1054(.A1(new_n670), .A2(G213), .ZN(new_n1255));
  XOR2_X1   g1055(.A(new_n1255), .B(KEYINPUT127), .Z(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  OAI211_X1 g1057(.A(G407), .B(G213), .C1(G375), .C2(new_n1257), .ZN(G409));
  OAI211_X1 g1058(.A(G378), .B(new_n1216), .C1(new_n1186), .C2(new_n1188), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1187), .A2(new_n1006), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1216), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1253), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1259), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1256), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1256), .A2(G2897), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1147), .A2(KEYINPUT60), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1219), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1174), .A2(KEYINPUT60), .A3(new_n1218), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1269), .A2(new_n686), .A3(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1271), .A2(G384), .A3(new_n1247), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(G384), .B1(new_n1271), .B2(new_n1247), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1267), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1271), .A2(new_n1247), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n845), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(new_n1272), .A3(new_n1266), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT61), .B1(new_n1265), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1281), .B1(new_n1265), .B2(new_n1283), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(G393), .B(new_n804), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(G387), .A2(G390), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1285), .B1(new_n1286), .B2(new_n1249), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1286), .A2(new_n1249), .A3(new_n1285), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1256), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1291), .A2(KEYINPUT63), .A3(new_n1282), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1280), .A2(new_n1284), .A3(new_n1290), .A4(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT62), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1291), .A2(new_n1294), .A3(new_n1282), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT61), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1296), .B1(new_n1291), .B2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1294), .B1(new_n1291), .B2(new_n1282), .ZN(new_n1299));
  NOR3_X1   g1099(.A1(new_n1295), .A2(new_n1298), .A3(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1293), .B1(new_n1300), .B2(new_n1290), .ZN(G405));
  INV_X1    g1101(.A(new_n1289), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1302), .A2(new_n1287), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(G375), .A2(new_n1253), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1304), .A2(new_n1283), .A3(new_n1259), .ZN(new_n1305));
  AOI21_X1  g1105(.A(G378), .B1(new_n1189), .B2(new_n1216), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1259), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1282), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1303), .A2(new_n1305), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1303), .B1(new_n1308), .B2(new_n1305), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(G402));
endmodule


