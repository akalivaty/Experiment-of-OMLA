//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n824, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950;
  INV_X1    g000(.A(G8gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n203), .A2(G1gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n205), .B2(G1gat), .ZN(new_n206));
  AND2_X1   g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n202), .B1(new_n207), .B2(KEYINPUT94), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(KEYINPUT94), .B2(new_n206), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(KEYINPUT95), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n202), .B(new_n210), .C1(new_n207), .C2(KEYINPUT95), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT21), .ZN(new_n212));
  NAND2_X1  g011(.A1(G71gat), .A2(G78gat), .ZN(new_n213));
  OR2_X1    g012(.A1(G71gat), .A2(G78gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(G57gat), .B(G64gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(KEYINPUT99), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT9), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n213), .B(new_n214), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n215), .B(KEYINPUT100), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n213), .B1(new_n214), .B2(new_n217), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n209), .B(new_n211), .C1(new_n212), .C2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(G183gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n222), .A2(new_n212), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n227), .B(G211gat), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n226), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G127gat), .B(G155gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(G231gat), .A2(G233gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n229), .B(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G232gat), .A2(G233gat), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n235), .B(KEYINPUT101), .Z(new_n236));
  INV_X1    g035(.A(KEYINPUT41), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XOR2_X1   g037(.A(G134gat), .B(G162gat), .Z(new_n239));
  XOR2_X1   g038(.A(new_n238), .B(new_n239), .Z(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT17), .ZN(new_n242));
  INV_X1    g041(.A(G43gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G50gat), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n244), .A2(KEYINPUT90), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(KEYINPUT15), .ZN(new_n246));
  INV_X1    g045(.A(G50gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G43gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n244), .A2(new_n248), .A3(KEYINPUT90), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n246), .A2(new_n249), .B1(G29gat), .B2(G36gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n244), .A2(new_n248), .A3(KEYINPUT15), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT89), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT88), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT14), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(KEYINPUT88), .A2(KEYINPUT14), .ZN(new_n257));
  OAI22_X1  g056(.A1(new_n256), .A2(new_n257), .B1(G29gat), .B2(G36gat), .ZN(new_n258));
  INV_X1    g057(.A(G29gat), .ZN(new_n259));
  INV_X1    g058(.A(G36gat), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n259), .B(new_n260), .C1(new_n254), .C2(new_n255), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n262), .A2(KEYINPUT91), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT91), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n264), .B1(new_n258), .B2(new_n261), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n250), .B(new_n253), .C1(new_n263), .C2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n262), .B1(new_n259), .B2(new_n260), .ZN(new_n267));
  INV_X1    g066(.A(new_n251), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n266), .A2(KEYINPUT92), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT92), .B1(new_n266), .B2(new_n269), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n242), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT93), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g073(.A(KEYINPUT93), .B(new_n242), .C1(new_n270), .C2(new_n271), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n266), .A2(new_n269), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT96), .B1(new_n277), .B2(new_n242), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT96), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n266), .A2(new_n279), .A3(KEYINPUT17), .A4(new_n269), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G85gat), .ZN(new_n282));
  INV_X1    g081(.A(G92gat), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT102), .ZN(new_n284));
  OR2_X1    g083(.A1(new_n284), .A2(KEYINPUT7), .ZN(new_n285));
  NAND2_X1  g084(.A1(G99gat), .A2(G106gat), .ZN(new_n286));
  AOI22_X1  g085(.A1(KEYINPUT8), .A2(new_n286), .B1(new_n282), .B2(new_n283), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n284), .A2(KEYINPUT7), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G99gat), .B(G106gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n281), .A3(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n236), .A2(new_n237), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT92), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n277), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n266), .A2(KEYINPUT92), .A3(new_n269), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n294), .B1(new_n298), .B2(new_n291), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n293), .A2(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(G190gat), .B(G218gat), .Z(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n293), .A2(new_n301), .A3(new_n299), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n241), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT103), .ZN(new_n306));
  OR2_X1    g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n306), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n303), .A2(KEYINPUT104), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT104), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n300), .A2(new_n310), .A3(new_n302), .ZN(new_n311));
  AND3_X1   g110(.A1(new_n309), .A2(new_n304), .A3(new_n311), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n307), .A2(new_n308), .B1(new_n312), .B2(new_n241), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n291), .B(new_n222), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT10), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n291), .A2(KEYINPUT10), .A3(new_n221), .A4(new_n218), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G230gat), .ZN(new_n319));
  INV_X1    g118(.A(G233gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n314), .A2(new_n322), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G120gat), .B(G148gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(G176gat), .B(G204gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n328), .B1(new_n324), .B2(KEYINPUT105), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n330), .B(new_n323), .C1(KEYINPUT105), .C2(new_n324), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n234), .A2(new_n313), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT98), .ZN(new_n335));
  XNOR2_X1  g134(.A(G141gat), .B(G148gat), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT77), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  XOR2_X1   g137(.A(G155gat), .B(G162gat), .Z(new_n339));
  XOR2_X1   g138(.A(KEYINPUT78), .B(KEYINPUT2), .Z(new_n340));
  NAND2_X1  g139(.A1(new_n336), .A2(new_n337), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .A4(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT80), .B(G162gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G155gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT79), .B(G141gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G148gat), .ZN(new_n346));
  INV_X1    g145(.A(G148gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G141gat), .ZN(new_n348));
  AOI22_X1  g147(.A1(KEYINPUT2), .A2(new_n344), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n342), .B1(new_n349), .B2(new_n339), .ZN(new_n350));
  NAND2_X1  g149(.A1(G211gat), .A2(G218gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(G197gat), .A2(G204gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(G197gat), .A2(G204gat), .ZN(new_n354));
  OAI22_X1  g153(.A1(new_n352), .A2(KEYINPUT22), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n355), .A2(KEYINPUT74), .ZN(new_n356));
  XNOR2_X1  g155(.A(G211gat), .B(G218gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n356), .B(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT3), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n350), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n350), .A2(new_n362), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n359), .B1(new_n364), .B2(new_n360), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  AND2_X1   g165(.A1(G228gat), .A2(G233gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n350), .ZN(new_n369));
  OR2_X1    g168(.A1(new_n355), .A2(new_n357), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n357), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(new_n360), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT83), .ZN(new_n373));
  OR2_X1    g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n373), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(new_n362), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n365), .B1(new_n369), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n368), .B1(new_n367), .B2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G78gat), .B(G106gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT31), .B(G50gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  OR3_X1    g180(.A1(new_n378), .A2(G22gat), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT84), .B1(new_n378), .B2(new_n381), .ZN(new_n383));
  OAI21_X1  g182(.A(G22gat), .B1(new_n378), .B2(new_n381), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n383), .B1(new_n382), .B2(new_n384), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AND2_X1   g186(.A1(G169gat), .A2(G176gat), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NOR3_X1   g190(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n389), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT64), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AND3_X1   g194(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(G183gat), .A2(G190gat), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT23), .ZN(new_n401));
  INV_X1    g200(.A(G169gat), .ZN(new_n402));
  INV_X1    g201(.A(G176gat), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n390), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(KEYINPUT64), .A3(new_n389), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n395), .A2(new_n400), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT65), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT25), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n408), .B1(new_n407), .B2(new_n409), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT66), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n404), .A2(new_n390), .B1(new_n412), .B2(new_n389), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n388), .A2(KEYINPUT66), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n413), .A2(new_n400), .A3(KEYINPUT25), .A4(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n410), .A2(new_n411), .A3(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT27), .B(G183gat), .ZN(new_n418));
  INV_X1    g217(.A(G190gat), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT67), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n420), .B(KEYINPUT28), .Z(new_n421));
  OR3_X1    g220(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(new_n389), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G183gat), .A2(G190gat), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n421), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  AND2_X1   g226(.A1(G226gat), .A2(G233gat), .ZN(new_n428));
  OAI22_X1  g227(.A1(new_n417), .A2(new_n427), .B1(KEYINPUT29), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT64), .B1(new_n405), .B2(new_n389), .ZN(new_n430));
  AOI211_X1 g229(.A(new_n394), .B(new_n388), .C1(new_n404), .C2(new_n390), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n430), .A2(new_n431), .A3(new_n399), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT65), .B1(new_n432), .B2(KEYINPUT25), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n434), .A3(new_n415), .ZN(new_n435));
  INV_X1    g234(.A(new_n428), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n436), .A3(new_n426), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n429), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n359), .ZN(new_n439));
  INV_X1    g238(.A(new_n359), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n429), .A2(new_n440), .A3(new_n437), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT75), .B(G8gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(G36gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(G64gat), .B(G92gat), .ZN(new_n445));
  XOR2_X1   g244(.A(new_n444), .B(new_n445), .Z(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT30), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(KEYINPUT76), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT76), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n446), .B1(new_n439), .B2(new_n441), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n451), .B1(new_n452), .B2(KEYINPUT30), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(KEYINPUT30), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n439), .A2(new_n446), .A3(new_n441), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n450), .A2(new_n453), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(G1gat), .B(G29gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n457), .B(new_n282), .ZN(new_n458));
  XNOR2_X1  g257(.A(KEYINPUT0), .B(G57gat), .ZN(new_n459));
  XOR2_X1   g258(.A(new_n458), .B(new_n459), .Z(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT82), .ZN(new_n462));
  NAND2_X1  g261(.A1(G225gat), .A2(G233gat), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT1), .ZN(new_n464));
  XOR2_X1   g263(.A(G127gat), .B(G134gat), .Z(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  XOR2_X1   g265(.A(KEYINPUT70), .B(G120gat), .Z(new_n467));
  INV_X1    g266(.A(G113gat), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(G120gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(KEYINPUT71), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n464), .B(new_n466), .C1(new_n469), .C2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(G113gat), .B(G120gat), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT68), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT1), .B1(new_n473), .B2(new_n474), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n466), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT69), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(G120gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(G113gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n470), .A2(new_n481), .A3(new_n474), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n464), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n473), .A2(new_n474), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n465), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n485), .A2(KEYINPUT69), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n472), .B1(new_n479), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(new_n369), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n350), .B(new_n472), .C1(new_n479), .C2(new_n486), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n463), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT5), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n462), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n463), .ZN(new_n493));
  INV_X1    g292(.A(new_n489), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n478), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n485), .A2(KEYINPUT69), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n350), .B1(new_n497), .B2(new_n472), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n493), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT81), .B1(new_n492), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n489), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n369), .A2(KEYINPUT3), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n505), .A2(new_n364), .A3(new_n487), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n502), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n507), .A2(new_n493), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n501), .A2(new_n508), .A3(new_n491), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n507), .A2(new_n493), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n492), .A2(new_n500), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(KEYINPUT81), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n461), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT81), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n515), .A2(KEYINPUT5), .A3(new_n510), .ZN(new_n516));
  INV_X1    g315(.A(new_n512), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(new_n460), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT6), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n513), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT6), .A4(new_n460), .ZN(new_n521));
  AOI211_X1 g320(.A(KEYINPUT35), .B(new_n456), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n487), .B1(new_n417), .B2(new_n427), .ZN(new_n523));
  INV_X1    g322(.A(new_n472), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n524), .B1(new_n496), .B2(new_n495), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n435), .A2(new_n426), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G227gat), .A2(G233gat), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT34), .B1(new_n529), .B2(KEYINPUT73), .ZN(new_n532));
  XNOR2_X1  g331(.A(G15gat), .B(G43gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(G71gat), .B(G99gat), .ZN(new_n534));
  XOR2_X1   g333(.A(new_n533), .B(new_n534), .Z(new_n535));
  AOI21_X1  g334(.A(new_n528), .B1(new_n523), .B2(new_n526), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT32), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT33), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n535), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT72), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n435), .A2(new_n426), .A3(new_n525), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n525), .B1(new_n435), .B2(new_n426), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n529), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n538), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n546), .A2(KEYINPUT72), .A3(new_n535), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n535), .A2(KEYINPUT33), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n545), .A2(KEYINPUT32), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n532), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n532), .ZN(new_n553));
  AOI211_X1 g352(.A(new_n553), .B(new_n550), .C1(new_n542), .C2(new_n547), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n531), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT72), .B1(new_n546), .B2(new_n535), .ZN(new_n556));
  INV_X1    g355(.A(new_n535), .ZN(new_n557));
  AOI211_X1 g356(.A(new_n541), .B(new_n557), .C1(new_n545), .C2(new_n538), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n551), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n553), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n548), .A2(new_n532), .A3(new_n551), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(new_n530), .A3(new_n561), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n555), .A2(KEYINPUT86), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT86), .B1(new_n555), .B2(new_n562), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n387), .B(new_n522), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT87), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n520), .A2(new_n521), .ZN(new_n568));
  INV_X1    g367(.A(new_n456), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n555), .A2(new_n387), .A3(new_n562), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT35), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT86), .ZN(new_n573));
  NOR3_X1   g372(.A1(new_n552), .A2(new_n554), .A3(new_n531), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n530), .B1(new_n560), .B2(new_n561), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n555), .A2(KEYINPUT86), .A3(new_n562), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n578), .A2(KEYINPUT87), .A3(new_n387), .A4(new_n522), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n567), .A2(new_n572), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n568), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n442), .B(KEYINPUT37), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(new_n446), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n583), .B1(KEYINPUT38), .B2(new_n452), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n581), .B(new_n584), .C1(KEYINPUT38), .C2(new_n583), .ZN(new_n585));
  NOR3_X1   g384(.A1(new_n494), .A2(new_n498), .A3(new_n493), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT85), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n507), .A2(new_n493), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT85), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g389(.A(KEYINPUT39), .B(new_n587), .C1(new_n590), .C2(new_n586), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n507), .A2(new_n493), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n591), .B(new_n461), .C1(KEYINPUT39), .C2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT40), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(new_n518), .A3(new_n456), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n585), .A2(new_n595), .A3(new_n387), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n597));
  NOR3_X1   g396(.A1(new_n574), .A2(new_n575), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT36), .B1(new_n555), .B2(new_n562), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n387), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n570), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n596), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n580), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n209), .A2(new_n211), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n606), .B1(new_n278), .B2(new_n280), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT93), .B1(new_n298), .B2(new_n242), .ZN(new_n608));
  INV_X1    g407(.A(new_n275), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n298), .ZN(new_n611));
  INV_X1    g410(.A(new_n606), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G229gat), .A2(G233gat), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n610), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT18), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n611), .A2(new_n612), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n615), .B(KEYINPUT13), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n613), .B1(new_n276), .B2(new_n607), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(KEYINPUT18), .A3(new_n615), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n618), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G113gat), .B(G141gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(G197gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT11), .B(G169gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n628), .B(new_n629), .Z(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  NAND2_X1  g430(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n631), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n618), .A2(new_n625), .A3(new_n623), .A4(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n634), .A2(KEYINPUT97), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(KEYINPUT97), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n335), .B1(new_n605), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT18), .B1(new_n624), .B2(new_n615), .ZN(new_n640));
  AND4_X1   g439(.A1(KEYINPUT18), .A2(new_n610), .A3(new_n614), .A4(new_n615), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT97), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n642), .A2(new_n643), .A3(new_n623), .A4(new_n633), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n634), .A2(KEYINPUT97), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n644), .A2(new_n645), .B1(new_n626), .B2(new_n631), .ZN(new_n646));
  AOI211_X1 g445(.A(KEYINPUT98), .B(new_n646), .C1(new_n580), .C2(new_n604), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n334), .B1(new_n639), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n568), .B(KEYINPUT106), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(G1gat), .ZN(G1324gat));
  INV_X1    g451(.A(KEYINPUT42), .ZN(new_n653));
  INV_X1    g452(.A(new_n334), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n456), .B(new_n654), .C1(new_n638), .C2(new_n647), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT16), .B(G8gat), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT107), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OR3_X1    g458(.A1(new_n655), .A2(new_n653), .A3(new_n656), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n655), .A2(G8gat), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n657), .A2(new_n658), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n659), .A2(new_n660), .A3(new_n661), .A4(new_n662), .ZN(G1325gat));
  AOI21_X1  g462(.A(G15gat), .B1(new_n649), .B2(new_n578), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n600), .A2(G15gat), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n664), .B1(new_n649), .B2(new_n665), .ZN(G1326gat));
  NAND2_X1  g465(.A1(new_n649), .A2(new_n602), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT43), .B(G22gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  NOR2_X1   g468(.A1(new_n234), .A2(new_n332), .ZN(new_n670));
  INV_X1    g469(.A(new_n313), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n673), .B1(new_n638), .B2(new_n647), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT108), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n675), .A2(new_n676), .A3(new_n259), .A4(new_n650), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n259), .B(new_n673), .C1(new_n638), .C2(new_n647), .ZN(new_n678));
  INV_X1    g477(.A(new_n650), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT108), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT45), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n684), .B1(new_n605), .B2(new_n671), .ZN(new_n685));
  AOI211_X1 g484(.A(KEYINPUT44), .B(new_n313), .C1(new_n580), .C2(new_n604), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n637), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT109), .Z(new_n689));
  NAND3_X1  g488(.A1(new_n687), .A2(new_n650), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(G29gat), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n677), .A2(new_n680), .A3(KEYINPUT45), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n683), .A2(new_n691), .A3(new_n692), .ZN(G1328gat));
  NAND2_X1  g492(.A1(new_n675), .A2(new_n260), .ZN(new_n694));
  OR3_X1    g493(.A1(new_n694), .A2(KEYINPUT46), .A3(new_n569), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n687), .A2(new_n456), .A3(new_n689), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(G36gat), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT46), .B1(new_n694), .B2(new_n569), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(G1329gat));
  NAND4_X1  g498(.A1(new_n687), .A2(G43gat), .A3(new_n600), .A4(new_n689), .ZN(new_n700));
  INV_X1    g499(.A(new_n578), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n243), .B1(new_n674), .B2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n700), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT111), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n700), .A2(new_n702), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(KEYINPUT47), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT111), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n700), .A2(new_n702), .A3(new_n708), .A4(new_n703), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n705), .A2(new_n707), .A3(new_n709), .ZN(G1330gat));
  NAND3_X1  g509(.A1(new_n687), .A2(new_n602), .A3(new_n689), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G50gat), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT48), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n675), .A2(new_n247), .A3(new_n602), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n713), .B1(new_n712), .B2(new_n714), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(G1331gat));
  AOI211_X1 g516(.A(new_n637), .B(new_n333), .C1(new_n580), .C2(new_n604), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n234), .A2(new_n313), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n650), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g522(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n721), .A2(new_n456), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT112), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT112), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n721), .A2(new_n727), .A3(new_n456), .A4(new_n724), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  OR2_X1    g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1333gat));
  NAND4_X1  g530(.A1(new_n718), .A2(G71gat), .A3(new_n600), .A4(new_n720), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT113), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n721), .A2(new_n578), .ZN(new_n734));
  INV_X1    g533(.A(G71gat), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT50), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT50), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n733), .A2(new_n739), .A3(new_n736), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(G1334gat));
  NAND2_X1  g540(.A1(new_n721), .A2(new_n602), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g542(.A1(new_n233), .A2(new_n646), .ZN(new_n744));
  XOR2_X1   g543(.A(new_n744), .B(KEYINPUT114), .Z(new_n745));
  OAI211_X1 g544(.A(new_n332), .B(new_n745), .C1(new_n685), .C2(new_n686), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n746), .A2(new_n282), .A3(new_n679), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n605), .A2(new_n671), .A3(new_n745), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n749), .A2(KEYINPUT115), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n313), .B1(new_n580), .B2(new_n604), .ZN(new_n752));
  INV_X1    g551(.A(new_n750), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n749), .A2(KEYINPUT115), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n752), .A2(new_n753), .A3(new_n745), .A4(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n751), .A2(new_n332), .A3(new_n755), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n756), .A2(new_n679), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n747), .B1(new_n757), .B2(new_n282), .ZN(G1336gat));
  INV_X1    g557(.A(KEYINPUT116), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n751), .A2(new_n755), .A3(new_n456), .A4(new_n332), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n760), .A2(new_n283), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n746), .A2(new_n283), .A3(new_n569), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT52), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n759), .B(new_n765), .C1(new_n761), .C2(new_n762), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(G1337gat));
  OAI21_X1  g566(.A(G99gat), .B1(new_n746), .B2(new_n601), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n756), .A2(G99gat), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n769), .B2(new_n701), .ZN(G1338gat));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n751), .A2(new_n755), .A3(new_n602), .A4(new_n332), .ZN(new_n772));
  INV_X1    g571(.A(G106gat), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n746), .A2(new_n773), .A3(new_n387), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n771), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT53), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n771), .B(new_n778), .C1(new_n774), .C2(new_n775), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1339gat));
  INV_X1    g579(.A(new_n630), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n624), .A2(new_n615), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n614), .A2(new_n619), .A3(new_n621), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n332), .B(new_n785), .C1(new_n635), .C2(new_n636), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT119), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n316), .A2(new_n317), .A3(new_n321), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n323), .A2(KEYINPUT54), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT118), .ZN(new_n790));
  INV_X1    g589(.A(new_n328), .ZN(new_n791));
  INV_X1    g590(.A(new_n323), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n323), .A2(new_n795), .A3(KEYINPUT54), .A4(new_n788), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n790), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n790), .A2(new_n794), .A3(KEYINPUT55), .A4(new_n796), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(new_n331), .A3(new_n800), .ZN(new_n801));
  OAI22_X1  g600(.A1(new_n786), .A2(new_n787), .B1(new_n646), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n784), .B1(new_n644), .B2(new_n645), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT119), .B1(new_n803), .B2(new_n332), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n313), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n799), .A2(new_n331), .A3(new_n800), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n671), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n234), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n334), .A2(new_n637), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n810), .A2(new_n650), .ZN(new_n811));
  INV_X1    g610(.A(new_n571), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n813), .A2(new_n569), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n814), .A2(new_n468), .A3(new_n637), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n701), .A2(new_n602), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n811), .A2(new_n569), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(G113gat), .B1(new_n817), .B2(new_n646), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(new_n818), .ZN(G1340gat));
  INV_X1    g618(.A(new_n467), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n814), .A2(new_n820), .A3(new_n332), .ZN(new_n821));
  OAI21_X1  g620(.A(G120gat), .B1(new_n817), .B2(new_n333), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(G1341gat));
  INV_X1    g622(.A(G127gat), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n817), .A2(new_n824), .A3(new_n233), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n814), .A2(new_n234), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n825), .B1(new_n826), .B2(new_n824), .ZN(G1342gat));
  INV_X1    g626(.A(G134gat), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n313), .A2(new_n456), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  OR2_X1    g629(.A1(new_n830), .A2(KEYINPUT56), .ZN(new_n831));
  OAI21_X1  g630(.A(G134gat), .B1(new_n817), .B2(new_n313), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(KEYINPUT56), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(G1343gat));
  NOR2_X1   g633(.A1(new_n679), .A2(new_n600), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n569), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n838), .B(new_n602), .C1(new_n808), .C2(new_n809), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n644), .A2(new_n645), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n801), .B1(new_n840), .B2(new_n632), .ZN(new_n841));
  AOI211_X1 g640(.A(new_n333), .B(new_n784), .C1(new_n644), .C2(new_n645), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT120), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n637), .A2(new_n806), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n845), .A3(new_n786), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n671), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n807), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n233), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n809), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n387), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n837), .B(new_n839), .C1(new_n851), .C2(new_n838), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(new_n646), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n602), .B1(new_n808), .B2(new_n809), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(new_n836), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n646), .A2(G141gat), .ZN(new_n857));
  OAI22_X1  g656(.A1(new_n853), .A2(new_n345), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT58), .ZN(G1344gat));
  NAND2_X1  g658(.A1(new_n854), .A2(KEYINPUT57), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n387), .A2(KEYINPUT57), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n841), .A2(new_n842), .A3(KEYINPUT120), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n845), .B1(new_n844), .B2(new_n786), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n313), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n671), .A2(KEYINPUT122), .A3(new_n806), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n866), .B1(new_n313), .B2(new_n801), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(new_n867), .A3(new_n803), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n234), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n861), .B1(new_n869), .B2(new_n809), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n860), .A2(new_n870), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n871), .A2(new_n333), .A3(new_n836), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT59), .B1(new_n872), .B2(new_n347), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n851), .A2(new_n838), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n875), .A2(new_n332), .A3(new_n837), .A4(new_n839), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n347), .A2(KEYINPUT59), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n874), .B(new_n877), .C1(new_n852), .C2(new_n333), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n873), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n855), .A2(new_n347), .A3(new_n332), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(G1345gat));
  AOI21_X1  g682(.A(G155gat), .B1(new_n855), .B2(new_n234), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n852), .A2(new_n233), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(G155gat), .ZN(G1346gat));
  OR3_X1    g685(.A1(new_n852), .A2(KEYINPUT123), .A3(new_n313), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT123), .B1(new_n852), .B2(new_n313), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n887), .A2(new_n343), .A3(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n854), .ZN(new_n890));
  INV_X1    g689(.A(new_n343), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n890), .A2(new_n891), .A3(new_n829), .A4(new_n835), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n889), .A2(new_n892), .ZN(G1347gat));
  AND3_X1   g692(.A1(new_n810), .A2(new_n456), .A3(new_n679), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n812), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n402), .A3(new_n637), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n810), .A2(new_n456), .A3(new_n816), .A4(new_n679), .ZN(new_n898));
  OAI21_X1  g697(.A(G169gat), .B1(new_n898), .B2(new_n646), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(G1348gat));
  NOR3_X1   g699(.A1(new_n898), .A2(new_n403), .A3(new_n333), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n896), .A2(new_n332), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n902), .B2(new_n403), .ZN(G1349gat));
  OAI21_X1  g702(.A(G183gat), .B1(new_n898), .B2(new_n233), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n234), .A2(new_n418), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n895), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g706(.A(G190gat), .B1(new_n898), .B2(new_n313), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n908), .A2(KEYINPUT124), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(KEYINPUT124), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(KEYINPUT61), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n419), .A3(new_n671), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT61), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n908), .A2(KEYINPUT124), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(G1351gat));
  NOR2_X1   g714(.A1(new_n600), .A2(new_n569), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n679), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n871), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n637), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(G197gat), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n854), .A2(new_n917), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n922), .A2(G197gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n920), .B1(new_n646), .B2(new_n923), .ZN(G1352gat));
  INV_X1    g723(.A(G204gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n921), .A2(new_n925), .A3(new_n332), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n926), .A2(KEYINPUT62), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(KEYINPUT62), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n871), .A2(new_n333), .ZN(new_n930));
  INV_X1    g729(.A(new_n917), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n925), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT125), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n930), .A2(new_n931), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G204gat), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n935), .A2(new_n936), .A3(new_n928), .A4(new_n927), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n933), .A2(new_n937), .ZN(G1353gat));
  NAND4_X1  g737(.A1(new_n860), .A2(new_n870), .A3(new_n234), .A4(new_n931), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n939), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT63), .B1(new_n939), .B2(G211gat), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n233), .A2(G211gat), .ZN(new_n942));
  OAI22_X1  g741(.A1(new_n940), .A2(new_n941), .B1(new_n922), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT126), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n945));
  OAI221_X1 g744(.A(new_n945), .B1(new_n922), .B2(new_n942), .C1(new_n940), .C2(new_n941), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(G1354gat));
  AOI21_X1  g746(.A(G218gat), .B1(new_n921), .B2(new_n671), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n671), .A2(G218gat), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT127), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n948), .B1(new_n918), .B2(new_n950), .ZN(G1355gat));
endmodule


