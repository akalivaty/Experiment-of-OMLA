

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U550 ( .A1(G2105), .A2(G2104), .ZN(n543) );
  OR2_X1 U551 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U552 ( .A1(G8), .A2(n729), .ZN(n802) );
  AND2_X1 U553 ( .A1(n706), .A2(G1996), .ZN(n707) );
  AND2_X1 U554 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U555 ( .A(n546), .B(KEYINPUT83), .Z(n514) );
  AND2_X1 U556 ( .A1(n705), .A2(n704), .ZN(n515) );
  XOR2_X1 U557 ( .A(n699), .B(KEYINPUT31), .Z(n516) );
  NOR2_X1 U558 ( .A1(n729), .A2(n713), .ZN(n715) );
  NOR2_X1 U559 ( .A1(n702), .A2(n701), .ZN(n709) );
  NOR2_X1 U560 ( .A1(n698), .A2(n697), .ZN(n699) );
  INV_X1 U561 ( .A(n989), .ZN(n753) );
  NOR2_X1 U562 ( .A1(n683), .A2(n682), .ZN(n685) );
  NOR2_X1 U563 ( .A1(G651), .A2(G543), .ZN(n645) );
  NOR2_X1 U564 ( .A1(G651), .A2(n624), .ZN(n653) );
  NAND2_X1 U565 ( .A1(n645), .A2(G91), .ZN(n520) );
  INV_X1 U566 ( .A(G651), .ZN(n522) );
  NOR2_X1 U567 ( .A1(G543), .A2(n522), .ZN(n517) );
  XOR2_X1 U568 ( .A(KEYINPUT1), .B(n517), .Z(n518) );
  XNOR2_X1 U569 ( .A(KEYINPUT66), .B(n518), .ZN(n649) );
  NAND2_X1 U570 ( .A1(G65), .A2(n649), .ZN(n519) );
  NAND2_X1 U571 ( .A1(n520), .A2(n519), .ZN(n526) );
  XNOR2_X1 U572 ( .A(G543), .B(KEYINPUT0), .ZN(n521) );
  XNOR2_X1 U573 ( .A(n521), .B(KEYINPUT65), .ZN(n624) );
  NOR2_X1 U574 ( .A1(n624), .A2(n522), .ZN(n646) );
  NAND2_X1 U575 ( .A1(G78), .A2(n646), .ZN(n524) );
  NAND2_X1 U576 ( .A1(G53), .A2(n653), .ZN(n523) );
  NAND2_X1 U577 ( .A1(n524), .A2(n523), .ZN(n525) );
  OR2_X1 U578 ( .A1(n526), .A2(n525), .ZN(G299) );
  XOR2_X1 U579 ( .A(G2438), .B(G2454), .Z(n528) );
  XNOR2_X1 U580 ( .A(G2435), .B(G2430), .ZN(n527) );
  XNOR2_X1 U581 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U582 ( .A(n529), .B(KEYINPUT104), .Z(n531) );
  XNOR2_X1 U583 ( .A(G1348), .B(G1341), .ZN(n530) );
  XNOR2_X1 U584 ( .A(n531), .B(n530), .ZN(n535) );
  XOR2_X1 U585 ( .A(G2446), .B(G2451), .Z(n533) );
  XNOR2_X1 U586 ( .A(G2443), .B(G2427), .ZN(n532) );
  XNOR2_X1 U587 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U588 ( .A(n535), .B(n534), .Z(n536) );
  AND2_X1 U589 ( .A1(G14), .A2(n536), .ZN(G401) );
  AND2_X1 U590 ( .A1(G2105), .A2(G2104), .ZN(n885) );
  NAND2_X1 U591 ( .A1(G114), .A2(n885), .ZN(n537) );
  XNOR2_X1 U592 ( .A(n537), .B(KEYINPUT82), .ZN(n541) );
  INV_X1 U593 ( .A(KEYINPUT81), .ZN(n539) );
  XOR2_X1 U594 ( .A(G2104), .B(KEYINPUT64), .Z(n542) );
  AND2_X2 U595 ( .A1(G2105), .A2(n542), .ZN(n886) );
  NAND2_X1 U596 ( .A1(G126), .A2(n886), .ZN(n538) );
  XNOR2_X1 U597 ( .A(n539), .B(n538), .ZN(n540) );
  NAND2_X1 U598 ( .A1(n541), .A2(n540), .ZN(n547) );
  NOR2_X4 U599 ( .A1(n542), .A2(G2105), .ZN(n881) );
  NAND2_X1 U600 ( .A1(G102), .A2(n881), .ZN(n545) );
  XOR2_X2 U601 ( .A(KEYINPUT17), .B(n543), .Z(n882) );
  NAND2_X1 U602 ( .A1(G138), .A2(n882), .ZN(n544) );
  NAND2_X1 U603 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U604 ( .A1(n547), .A2(n514), .ZN(n548) );
  XNOR2_X1 U605 ( .A(KEYINPUT84), .B(n548), .ZN(G164) );
  NAND2_X1 U606 ( .A1(n653), .A2(G52), .ZN(n550) );
  NAND2_X1 U607 ( .A1(G64), .A2(n649), .ZN(n549) );
  NAND2_X1 U608 ( .A1(n550), .A2(n549), .ZN(n555) );
  NAND2_X1 U609 ( .A1(G90), .A2(n645), .ZN(n552) );
  NAND2_X1 U610 ( .A1(G77), .A2(n646), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U612 ( .A(KEYINPUT9), .B(n553), .Z(n554) );
  NOR2_X1 U613 ( .A1(n555), .A2(n554), .ZN(G171) );
  INV_X1 U614 ( .A(G57), .ZN(G237) );
  INV_X1 U615 ( .A(G132), .ZN(G219) );
  INV_X1 U616 ( .A(G82), .ZN(G220) );
  NAND2_X1 U617 ( .A1(n645), .A2(G89), .ZN(n556) );
  XNOR2_X1 U618 ( .A(n556), .B(KEYINPUT4), .ZN(n558) );
  NAND2_X1 U619 ( .A1(G76), .A2(n646), .ZN(n557) );
  NAND2_X1 U620 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U621 ( .A(n559), .B(KEYINPUT5), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n653), .A2(G51), .ZN(n561) );
  NAND2_X1 U623 ( .A1(G63), .A2(n649), .ZN(n560) );
  NAND2_X1 U624 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U625 ( .A(KEYINPUT6), .B(n562), .Z(n563) );
  NAND2_X1 U626 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U627 ( .A(n565), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U628 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U629 ( .A1(G101), .A2(n881), .ZN(n566) );
  XNOR2_X1 U630 ( .A(n566), .B(KEYINPUT23), .ZN(n567) );
  INV_X1 U631 ( .A(n567), .ZN(n569) );
  NAND2_X1 U632 ( .A1(n885), .A2(G113), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n683) );
  NAND2_X1 U634 ( .A1(G137), .A2(n882), .ZN(n571) );
  NAND2_X1 U635 ( .A1(G125), .A2(n886), .ZN(n570) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n681) );
  NOR2_X1 U637 ( .A1(n683), .A2(n681), .ZN(G160) );
  NAND2_X1 U638 ( .A1(G94), .A2(G452), .ZN(n572) );
  XOR2_X1 U639 ( .A(KEYINPUT68), .B(n572), .Z(G173) );
  NAND2_X1 U640 ( .A1(G7), .A2(G661), .ZN(n573) );
  XOR2_X1 U641 ( .A(n573), .B(KEYINPUT10), .Z(n912) );
  NAND2_X1 U642 ( .A1(n912), .A2(G567), .ZN(n574) );
  XOR2_X1 U643 ( .A(KEYINPUT11), .B(n574), .Z(G234) );
  NAND2_X1 U644 ( .A1(n649), .A2(G56), .ZN(n575) );
  XOR2_X1 U645 ( .A(KEYINPUT14), .B(n575), .Z(n581) );
  NAND2_X1 U646 ( .A1(n645), .A2(G81), .ZN(n576) );
  XNOR2_X1 U647 ( .A(n576), .B(KEYINPUT12), .ZN(n578) );
  NAND2_X1 U648 ( .A1(G68), .A2(n646), .ZN(n577) );
  NAND2_X1 U649 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U650 ( .A(KEYINPUT13), .B(n579), .Z(n580) );
  NOR2_X1 U651 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U652 ( .A1(n653), .A2(G43), .ZN(n582) );
  NAND2_X1 U653 ( .A1(n583), .A2(n582), .ZN(n984) );
  INV_X1 U654 ( .A(G860), .ZN(n597) );
  OR2_X1 U655 ( .A1(n984), .A2(n597), .ZN(G153) );
  XNOR2_X1 U656 ( .A(G171), .B(KEYINPUT69), .ZN(G301) );
  NAND2_X1 U657 ( .A1(G868), .A2(G301), .ZN(n584) );
  XNOR2_X1 U658 ( .A(n584), .B(KEYINPUT70), .ZN(n593) );
  INV_X1 U659 ( .A(G868), .ZN(n594) );
  NAND2_X1 U660 ( .A1(n645), .A2(G92), .ZN(n586) );
  NAND2_X1 U661 ( .A1(G66), .A2(n649), .ZN(n585) );
  NAND2_X1 U662 ( .A1(n586), .A2(n585), .ZN(n590) );
  NAND2_X1 U663 ( .A1(G79), .A2(n646), .ZN(n588) );
  NAND2_X1 U664 ( .A1(G54), .A2(n653), .ZN(n587) );
  NAND2_X1 U665 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U666 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U667 ( .A(KEYINPUT15), .B(n591), .ZN(n988) );
  NAND2_X1 U668 ( .A1(n594), .A2(n988), .ZN(n592) );
  NAND2_X1 U669 ( .A1(n593), .A2(n592), .ZN(G284) );
  NOR2_X1 U670 ( .A1(G286), .A2(n594), .ZN(n596) );
  NOR2_X1 U671 ( .A1(G868), .A2(G299), .ZN(n595) );
  NOR2_X1 U672 ( .A1(n596), .A2(n595), .ZN(G297) );
  NAND2_X1 U673 ( .A1(n597), .A2(G559), .ZN(n598) );
  INV_X1 U674 ( .A(n988), .ZN(n613) );
  NAND2_X1 U675 ( .A1(n598), .A2(n613), .ZN(n599) );
  XNOR2_X1 U676 ( .A(n599), .B(KEYINPUT71), .ZN(n600) );
  XOR2_X1 U677 ( .A(KEYINPUT16), .B(n600), .Z(G148) );
  NOR2_X1 U678 ( .A1(G868), .A2(n984), .ZN(n603) );
  NAND2_X1 U679 ( .A1(G868), .A2(n613), .ZN(n601) );
  NOR2_X1 U680 ( .A1(G559), .A2(n601), .ZN(n602) );
  NOR2_X1 U681 ( .A1(n603), .A2(n602), .ZN(G282) );
  NAND2_X1 U682 ( .A1(G99), .A2(n881), .ZN(n605) );
  NAND2_X1 U683 ( .A1(G111), .A2(n885), .ZN(n604) );
  NAND2_X1 U684 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U685 ( .A(KEYINPUT72), .B(n606), .ZN(n611) );
  NAND2_X1 U686 ( .A1(G123), .A2(n886), .ZN(n607) );
  XNOR2_X1 U687 ( .A(n607), .B(KEYINPUT18), .ZN(n609) );
  NAND2_X1 U688 ( .A1(n882), .A2(G135), .ZN(n608) );
  NAND2_X1 U689 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U690 ( .A1(n611), .A2(n610), .ZN(n941) );
  XNOR2_X1 U691 ( .A(G2096), .B(n941), .ZN(n612) );
  INV_X1 U692 ( .A(G2100), .ZN(n851) );
  NAND2_X1 U693 ( .A1(n612), .A2(n851), .ZN(G156) );
  NAND2_X1 U694 ( .A1(G559), .A2(n613), .ZN(n614) );
  XNOR2_X1 U695 ( .A(n984), .B(n614), .ZN(n662) );
  NOR2_X1 U696 ( .A1(n662), .A2(G860), .ZN(n623) );
  NAND2_X1 U697 ( .A1(G93), .A2(n645), .ZN(n616) );
  NAND2_X1 U698 ( .A1(G80), .A2(n646), .ZN(n615) );
  NAND2_X1 U699 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U700 ( .A1(G67), .A2(n649), .ZN(n617) );
  XNOR2_X1 U701 ( .A(KEYINPUT73), .B(n617), .ZN(n618) );
  NOR2_X1 U702 ( .A1(n619), .A2(n618), .ZN(n621) );
  NAND2_X1 U703 ( .A1(n653), .A2(G55), .ZN(n620) );
  NAND2_X1 U704 ( .A1(n621), .A2(n620), .ZN(n901) );
  XOR2_X1 U705 ( .A(n901), .B(KEYINPUT74), .Z(n622) );
  XNOR2_X1 U706 ( .A(n623), .B(n622), .ZN(G145) );
  NAND2_X1 U707 ( .A1(n653), .A2(G49), .ZN(n629) );
  NAND2_X1 U708 ( .A1(G87), .A2(n624), .ZN(n626) );
  NAND2_X1 U709 ( .A1(G74), .A2(G651), .ZN(n625) );
  NAND2_X1 U710 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U711 ( .A1(n649), .A2(n627), .ZN(n628) );
  NAND2_X1 U712 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U713 ( .A(KEYINPUT75), .B(n630), .Z(G288) );
  NAND2_X1 U714 ( .A1(G88), .A2(n645), .ZN(n632) );
  NAND2_X1 U715 ( .A1(G75), .A2(n646), .ZN(n631) );
  NAND2_X1 U716 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n653), .A2(G50), .ZN(n634) );
  NAND2_X1 U718 ( .A1(G62), .A2(n649), .ZN(n633) );
  NAND2_X1 U719 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U720 ( .A1(n636), .A2(n635), .ZN(G166) );
  INV_X1 U721 ( .A(G166), .ZN(G303) );
  NAND2_X1 U722 ( .A1(G73), .A2(n646), .ZN(n637) );
  XNOR2_X1 U723 ( .A(n637), .B(KEYINPUT2), .ZN(n644) );
  NAND2_X1 U724 ( .A1(n653), .A2(G48), .ZN(n639) );
  NAND2_X1 U725 ( .A1(G61), .A2(n649), .ZN(n638) );
  NAND2_X1 U726 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U727 ( .A1(n645), .A2(G86), .ZN(n640) );
  XOR2_X1 U728 ( .A(KEYINPUT76), .B(n640), .Z(n641) );
  NOR2_X1 U729 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U730 ( .A1(n644), .A2(n643), .ZN(G305) );
  NAND2_X1 U731 ( .A1(G85), .A2(n645), .ZN(n648) );
  NAND2_X1 U732 ( .A1(G72), .A2(n646), .ZN(n647) );
  NAND2_X1 U733 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U734 ( .A1(G60), .A2(n649), .ZN(n650) );
  XNOR2_X1 U735 ( .A(KEYINPUT67), .B(n650), .ZN(n651) );
  NOR2_X1 U736 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U737 ( .A1(n653), .A2(G47), .ZN(n654) );
  NAND2_X1 U738 ( .A1(n655), .A2(n654), .ZN(G290) );
  XOR2_X1 U739 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n657) );
  XOR2_X1 U740 ( .A(G303), .B(KEYINPUT19), .Z(n656) );
  XNOR2_X1 U741 ( .A(n657), .B(n656), .ZN(n658) );
  XOR2_X1 U742 ( .A(n658), .B(G305), .Z(n659) );
  XNOR2_X1 U743 ( .A(G288), .B(n659), .ZN(n661) );
  XOR2_X1 U744 ( .A(G290), .B(G299), .Z(n660) );
  XNOR2_X1 U745 ( .A(n661), .B(n660), .ZN(n902) );
  XOR2_X1 U746 ( .A(n662), .B(n902), .Z(n663) );
  NAND2_X1 U747 ( .A1(n663), .A2(G868), .ZN(n664) );
  XNOR2_X1 U748 ( .A(n664), .B(n901), .ZN(G295) );
  NAND2_X1 U749 ( .A1(G2084), .A2(G2078), .ZN(n665) );
  XOR2_X1 U750 ( .A(KEYINPUT20), .B(n665), .Z(n666) );
  NAND2_X1 U751 ( .A1(G2090), .A2(n666), .ZN(n667) );
  XNOR2_X1 U752 ( .A(KEYINPUT21), .B(n667), .ZN(n668) );
  NAND2_X1 U753 ( .A1(n668), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U755 ( .A1(G220), .A2(G219), .ZN(n669) );
  XOR2_X1 U756 ( .A(KEYINPUT22), .B(n669), .Z(n670) );
  NOR2_X1 U757 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U758 ( .A1(G96), .A2(n671), .ZN(n830) );
  NAND2_X1 U759 ( .A1(n830), .A2(G2106), .ZN(n677) );
  NAND2_X1 U760 ( .A1(G120), .A2(G69), .ZN(n672) );
  XNOR2_X1 U761 ( .A(KEYINPUT79), .B(n672), .ZN(n673) );
  NAND2_X1 U762 ( .A1(n673), .A2(G108), .ZN(n674) );
  NOR2_X1 U763 ( .A1(G237), .A2(n674), .ZN(n675) );
  XOR2_X1 U764 ( .A(KEYINPUT80), .B(n675), .Z(n831) );
  NAND2_X1 U765 ( .A1(n831), .A2(G567), .ZN(n676) );
  NAND2_X1 U766 ( .A1(n677), .A2(n676), .ZN(n832) );
  NAND2_X1 U767 ( .A1(G661), .A2(G483), .ZN(n678) );
  NOR2_X1 U768 ( .A1(n832), .A2(n678), .ZN(n829) );
  NAND2_X1 U769 ( .A1(n829), .A2(G36), .ZN(G176) );
  XOR2_X1 U770 ( .A(KEYINPUT25), .B(G2078), .Z(n915) );
  NOR2_X1 U771 ( .A1(G1384), .A2(G164), .ZN(n773) );
  INV_X1 U772 ( .A(G40), .ZN(n680) );
  OR2_X1 U773 ( .A1(n681), .A2(n680), .ZN(n682) );
  INV_X1 U774 ( .A(KEYINPUT86), .ZN(n684) );
  XNOR2_X1 U775 ( .A(n685), .B(n684), .ZN(n774) );
  XOR2_X1 U776 ( .A(n774), .B(KEYINPUT92), .Z(n686) );
  NAND2_X2 U777 ( .A1(n773), .A2(n686), .ZN(n729) );
  OR2_X1 U778 ( .A1(n915), .A2(n729), .ZN(n690) );
  INV_X1 U779 ( .A(G1961), .ZN(n687) );
  AND2_X1 U780 ( .A1(n729), .A2(n687), .ZN(n688) );
  XNOR2_X1 U781 ( .A(KEYINPUT93), .B(n688), .ZN(n689) );
  AND2_X1 U782 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U783 ( .A(KEYINPUT94), .B(n691), .Z(n700) );
  NOR2_X1 U784 ( .A1(G171), .A2(n700), .ZN(n698) );
  NOR2_X1 U785 ( .A1(G1966), .A2(n802), .ZN(n746) );
  NOR2_X1 U786 ( .A1(G2084), .A2(n729), .ZN(n742) );
  NOR2_X1 U787 ( .A1(n746), .A2(n742), .ZN(n693) );
  INV_X1 U788 ( .A(KEYINPUT99), .ZN(n692) );
  XNOR2_X1 U789 ( .A(n693), .B(n692), .ZN(n694) );
  NAND2_X1 U790 ( .A1(n694), .A2(G8), .ZN(n695) );
  XNOR2_X1 U791 ( .A(KEYINPUT30), .B(n695), .ZN(n696) );
  NOR2_X1 U792 ( .A1(n696), .A2(G168), .ZN(n697) );
  XNOR2_X1 U793 ( .A(n516), .B(KEYINPUT100), .ZN(n743) );
  NAND2_X1 U794 ( .A1(n700), .A2(G171), .ZN(n728) );
  INV_X1 U795 ( .A(n729), .ZN(n706) );
  NOR2_X1 U796 ( .A1(n706), .A2(G1348), .ZN(n702) );
  NOR2_X1 U797 ( .A1(G2067), .A2(n729), .ZN(n701) );
  NAND2_X1 U798 ( .A1(n988), .A2(n709), .ZN(n705) );
  AND2_X1 U799 ( .A1(n729), .A2(G1341), .ZN(n703) );
  NOR2_X1 U800 ( .A1(n703), .A2(n984), .ZN(n704) );
  XOR2_X1 U801 ( .A(n707), .B(KEYINPUT26), .Z(n708) );
  NAND2_X1 U802 ( .A1(n515), .A2(n708), .ZN(n711) );
  OR2_X1 U803 ( .A1(n709), .A2(n988), .ZN(n710) );
  NAND2_X1 U804 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U805 ( .A(KEYINPUT97), .B(n712), .Z(n721) );
  INV_X1 U806 ( .A(G2072), .ZN(n713) );
  XOR2_X1 U807 ( .A(KEYINPUT95), .B(KEYINPUT27), .Z(n714) );
  XNOR2_X1 U808 ( .A(n715), .B(n714), .ZN(n717) );
  NAND2_X1 U809 ( .A1(n729), .A2(G1956), .ZN(n716) );
  NAND2_X1 U810 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U811 ( .A(KEYINPUT96), .B(n718), .ZN(n722) );
  NOR2_X1 U812 ( .A1(n722), .A2(G299), .ZN(n719) );
  XNOR2_X1 U813 ( .A(KEYINPUT98), .B(n719), .ZN(n720) );
  NOR2_X1 U814 ( .A1(n721), .A2(n720), .ZN(n725) );
  NAND2_X1 U815 ( .A1(n722), .A2(G299), .ZN(n723) );
  XOR2_X1 U816 ( .A(KEYINPUT28), .B(n723), .Z(n724) );
  NOR2_X1 U817 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U818 ( .A(n726), .B(KEYINPUT29), .ZN(n727) );
  NAND2_X1 U819 ( .A1(n728), .A2(n727), .ZN(n744) );
  INV_X1 U820 ( .A(G8), .ZN(n734) );
  NOR2_X1 U821 ( .A1(G1971), .A2(n802), .ZN(n731) );
  NOR2_X1 U822 ( .A1(G2090), .A2(n729), .ZN(n730) );
  NOR2_X1 U823 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U824 ( .A1(n732), .A2(G303), .ZN(n733) );
  OR2_X1 U825 ( .A1(n734), .A2(n733), .ZN(n736) );
  AND2_X1 U826 ( .A1(n744), .A2(n736), .ZN(n735) );
  NAND2_X1 U827 ( .A1(n743), .A2(n735), .ZN(n739) );
  INV_X1 U828 ( .A(n736), .ZN(n737) );
  OR2_X1 U829 ( .A1(n737), .A2(G286), .ZN(n738) );
  NAND2_X1 U830 ( .A1(n739), .A2(n738), .ZN(n741) );
  XOR2_X1 U831 ( .A(KEYINPUT32), .B(KEYINPUT101), .Z(n740) );
  XNOR2_X1 U832 ( .A(n741), .B(n740), .ZN(n750) );
  NAND2_X1 U833 ( .A1(G8), .A2(n742), .ZN(n748) );
  AND2_X1 U834 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U835 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U837 ( .A1(n750), .A2(n749), .ZN(n798) );
  NOR2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n757) );
  NOR2_X1 U839 ( .A1(G1971), .A2(G303), .ZN(n751) );
  NOR2_X1 U840 ( .A1(n757), .A2(n751), .ZN(n1002) );
  NAND2_X1 U841 ( .A1(n798), .A2(n1002), .ZN(n755) );
  NAND2_X1 U842 ( .A1(G288), .A2(G1976), .ZN(n752) );
  XNOR2_X1 U843 ( .A(n752), .B(KEYINPUT102), .ZN(n989) );
  NOR2_X1 U844 ( .A1(n802), .A2(n753), .ZN(n754) );
  NOR2_X1 U845 ( .A1(KEYINPUT33), .A2(n756), .ZN(n760) );
  NAND2_X1 U846 ( .A1(n757), .A2(KEYINPUT33), .ZN(n758) );
  NOR2_X1 U847 ( .A1(n758), .A2(n802), .ZN(n759) );
  NOR2_X1 U848 ( .A1(n760), .A2(n759), .ZN(n795) );
  XOR2_X1 U849 ( .A(G1981), .B(G305), .Z(n991) );
  XNOR2_X1 U850 ( .A(G2067), .B(KEYINPUT37), .ZN(n820) );
  XNOR2_X1 U851 ( .A(KEYINPUT89), .B(KEYINPUT36), .ZN(n772) );
  NAND2_X1 U852 ( .A1(n885), .A2(G116), .ZN(n761) );
  XNOR2_X1 U853 ( .A(n761), .B(KEYINPUT88), .ZN(n763) );
  NAND2_X1 U854 ( .A1(G128), .A2(n886), .ZN(n762) );
  NAND2_X1 U855 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U856 ( .A(KEYINPUT35), .B(n764), .ZN(n770) );
  NAND2_X1 U857 ( .A1(n881), .A2(G104), .ZN(n765) );
  XOR2_X1 U858 ( .A(KEYINPUT87), .B(n765), .Z(n767) );
  NAND2_X1 U859 ( .A1(n882), .A2(G140), .ZN(n766) );
  NAND2_X1 U860 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U861 ( .A(KEYINPUT34), .B(n768), .Z(n769) );
  NAND2_X1 U862 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U863 ( .A(n772), .B(n771), .ZN(n896) );
  NOR2_X1 U864 ( .A1(n820), .A2(n896), .ZN(n954) );
  NOR2_X1 U865 ( .A1(n774), .A2(n773), .ZN(n822) );
  NAND2_X1 U866 ( .A1(n954), .A2(n822), .ZN(n775) );
  XNOR2_X1 U867 ( .A(n775), .B(KEYINPUT90), .ZN(n818) );
  NAND2_X1 U868 ( .A1(G95), .A2(n881), .ZN(n777) );
  NAND2_X1 U869 ( .A1(G107), .A2(n885), .ZN(n776) );
  NAND2_X1 U870 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U871 ( .A1(G131), .A2(n882), .ZN(n778) );
  XNOR2_X1 U872 ( .A(KEYINPUT91), .B(n778), .ZN(n779) );
  NOR2_X1 U873 ( .A1(n780), .A2(n779), .ZN(n782) );
  NAND2_X1 U874 ( .A1(n886), .A2(G119), .ZN(n781) );
  NAND2_X1 U875 ( .A1(n782), .A2(n781), .ZN(n875) );
  AND2_X1 U876 ( .A1(n875), .A2(G1991), .ZN(n791) );
  NAND2_X1 U877 ( .A1(G117), .A2(n885), .ZN(n784) );
  NAND2_X1 U878 ( .A1(G129), .A2(n886), .ZN(n783) );
  NAND2_X1 U879 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U880 ( .A1(n881), .A2(G105), .ZN(n785) );
  XOR2_X1 U881 ( .A(KEYINPUT38), .B(n785), .Z(n786) );
  NOR2_X1 U882 ( .A1(n787), .A2(n786), .ZN(n789) );
  NAND2_X1 U883 ( .A1(n882), .A2(G141), .ZN(n788) );
  NAND2_X1 U884 ( .A1(n789), .A2(n788), .ZN(n877) );
  AND2_X1 U885 ( .A1(n877), .A2(G1996), .ZN(n790) );
  NOR2_X1 U886 ( .A1(n791), .A2(n790), .ZN(n948) );
  INV_X1 U887 ( .A(n822), .ZN(n792) );
  NOR2_X1 U888 ( .A1(n948), .A2(n792), .ZN(n814) );
  INV_X1 U889 ( .A(n814), .ZN(n793) );
  AND2_X1 U890 ( .A1(n818), .A2(n793), .ZN(n806) );
  AND2_X1 U891 ( .A1(n991), .A2(n806), .ZN(n794) );
  NAND2_X1 U892 ( .A1(n795), .A2(n794), .ZN(n808) );
  NOR2_X1 U893 ( .A1(G2090), .A2(G303), .ZN(n796) );
  NAND2_X1 U894 ( .A1(G8), .A2(n796), .ZN(n797) );
  NAND2_X1 U895 ( .A1(n798), .A2(n797), .ZN(n799) );
  AND2_X1 U896 ( .A1(n799), .A2(n802), .ZN(n804) );
  NOR2_X1 U897 ( .A1(G1981), .A2(G305), .ZN(n800) );
  XOR2_X1 U898 ( .A(n800), .B(KEYINPUT24), .Z(n801) );
  NOR2_X1 U899 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U901 ( .A1(n808), .A2(n807), .ZN(n811) );
  XOR2_X1 U902 ( .A(G1986), .B(KEYINPUT85), .Z(n809) );
  XNOR2_X1 U903 ( .A(G290), .B(n809), .ZN(n1001) );
  NAND2_X1 U904 ( .A1(n1001), .A2(n822), .ZN(n810) );
  NAND2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n825) );
  NOR2_X1 U906 ( .A1(G1996), .A2(n877), .ZN(n939) );
  NOR2_X1 U907 ( .A1(G1991), .A2(n875), .ZN(n942) );
  NOR2_X1 U908 ( .A1(G1986), .A2(G290), .ZN(n812) );
  NOR2_X1 U909 ( .A1(n942), .A2(n812), .ZN(n813) );
  NOR2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U911 ( .A1(n939), .A2(n815), .ZN(n817) );
  XOR2_X1 U912 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n816) );
  XNOR2_X1 U913 ( .A(n817), .B(n816), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n820), .A2(n896), .ZN(n951) );
  NAND2_X1 U916 ( .A1(n821), .A2(n951), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U918 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U919 ( .A(n826), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n912), .ZN(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U922 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U924 ( .A1(n829), .A2(n828), .ZN(G188) );
  XNOR2_X1 U925 ( .A(G69), .B(KEYINPUT105), .ZN(G235) );
  NOR2_X1 U926 ( .A1(n831), .A2(n830), .ZN(G325) );
  XOR2_X1 U927 ( .A(KEYINPUT106), .B(G325), .Z(G261) );
  XNOR2_X1 U928 ( .A(G108), .B(KEYINPUT117), .ZN(G238) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  INV_X1 U932 ( .A(n832), .ZN(G319) );
  XOR2_X1 U933 ( .A(KEYINPUT110), .B(G1976), .Z(n834) );
  XNOR2_X1 U934 ( .A(G1956), .B(G1981), .ZN(n833) );
  XNOR2_X1 U935 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U936 ( .A(n835), .B(KEYINPUT41), .Z(n837) );
  XNOR2_X1 U937 ( .A(G1996), .B(G1991), .ZN(n836) );
  XNOR2_X1 U938 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U939 ( .A(G1971), .B(G1961), .Z(n839) );
  XNOR2_X1 U940 ( .A(G1986), .B(G1966), .ZN(n838) );
  XNOR2_X1 U941 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U942 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U943 ( .A(KEYINPUT111), .B(G2474), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(G229) );
  XNOR2_X1 U945 ( .A(G2067), .B(G2072), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n844), .B(KEYINPUT109), .ZN(n855) );
  XOR2_X1 U947 ( .A(G2678), .B(KEYINPUT108), .Z(n846) );
  XNOR2_X1 U948 ( .A(G2096), .B(KEYINPUT43), .ZN(n845) );
  XNOR2_X1 U949 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U950 ( .A(KEYINPUT107), .B(G2090), .Z(n848) );
  XNOR2_X1 U951 ( .A(G2084), .B(G2078), .ZN(n847) );
  XNOR2_X1 U952 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U953 ( .A(n850), .B(n849), .Z(n853) );
  XOR2_X1 U954 ( .A(KEYINPUT42), .B(n851), .Z(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(G227) );
  NAND2_X1 U957 ( .A1(G112), .A2(n885), .ZN(n857) );
  NAND2_X1 U958 ( .A1(G136), .A2(n882), .ZN(n856) );
  NAND2_X1 U959 ( .A1(n857), .A2(n856), .ZN(n863) );
  NAND2_X1 U960 ( .A1(G124), .A2(n886), .ZN(n858) );
  XNOR2_X1 U961 ( .A(n858), .B(KEYINPUT44), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n859), .B(KEYINPUT112), .ZN(n861) );
  NAND2_X1 U963 ( .A1(G100), .A2(n881), .ZN(n860) );
  NAND2_X1 U964 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U965 ( .A1(n863), .A2(n862), .ZN(G162) );
  NAND2_X1 U966 ( .A1(G106), .A2(n881), .ZN(n865) );
  NAND2_X1 U967 ( .A1(G142), .A2(n882), .ZN(n864) );
  NAND2_X1 U968 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U969 ( .A(n866), .B(KEYINPUT45), .ZN(n868) );
  NAND2_X1 U970 ( .A1(G118), .A2(n885), .ZN(n867) );
  NAND2_X1 U971 ( .A1(n868), .A2(n867), .ZN(n871) );
  NAND2_X1 U972 ( .A1(G130), .A2(n886), .ZN(n869) );
  XNOR2_X1 U973 ( .A(KEYINPUT113), .B(n869), .ZN(n870) );
  NOR2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U975 ( .A(n941), .B(n872), .ZN(n895) );
  XOR2_X1 U976 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n874) );
  XNOR2_X1 U977 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n873) );
  XNOR2_X1 U978 ( .A(n874), .B(n873), .ZN(n876) );
  XNOR2_X1 U979 ( .A(n876), .B(n875), .ZN(n879) );
  XOR2_X1 U980 ( .A(G160), .B(n877), .Z(n878) );
  XNOR2_X1 U981 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U982 ( .A(G162), .B(n880), .ZN(n893) );
  NAND2_X1 U983 ( .A1(G103), .A2(n881), .ZN(n884) );
  NAND2_X1 U984 ( .A1(G139), .A2(n882), .ZN(n883) );
  NAND2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n891) );
  NAND2_X1 U986 ( .A1(G115), .A2(n885), .ZN(n888) );
  NAND2_X1 U987 ( .A1(G127), .A2(n886), .ZN(n887) );
  NAND2_X1 U988 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  NOR2_X1 U990 ( .A1(n891), .A2(n890), .ZN(n933) );
  XNOR2_X1 U991 ( .A(G164), .B(n933), .ZN(n892) );
  XNOR2_X1 U992 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U993 ( .A(n895), .B(n894), .ZN(n897) );
  XOR2_X1 U994 ( .A(n897), .B(n896), .Z(n898) );
  NOR2_X1 U995 ( .A1(G37), .A2(n898), .ZN(G395) );
  XNOR2_X1 U996 ( .A(n984), .B(G286), .ZN(n900) );
  XOR2_X1 U997 ( .A(G171), .B(n988), .Z(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U999 ( .A(n902), .B(n901), .Z(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n905), .ZN(G397) );
  NOR2_X1 U1002 ( .A1(G229), .A2(G227), .ZN(n906) );
  XOR2_X1 U1003 ( .A(KEYINPUT49), .B(n906), .Z(n907) );
  NAND2_X1 U1004 ( .A1(G319), .A2(n907), .ZN(n908) );
  NOR2_X1 U1005 ( .A1(G401), .A2(n908), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(KEYINPUT116), .B(n909), .ZN(n911) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n910) );
  NAND2_X1 U1008 ( .A1(n911), .A2(n910), .ZN(G225) );
  INV_X1 U1009 ( .A(G225), .ZN(G308) );
  INV_X1 U1010 ( .A(n912), .ZN(G223) );
  XNOR2_X1 U1011 ( .A(G32), .B(G1996), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(n913), .B(KEYINPUT121), .ZN(n924) );
  XOR2_X1 U1013 ( .A(G25), .B(G1991), .Z(n914) );
  NAND2_X1 U1014 ( .A1(n914), .A2(G28), .ZN(n922) );
  XOR2_X1 U1015 ( .A(n915), .B(G27), .Z(n920) );
  XNOR2_X1 U1016 ( .A(G2067), .B(G26), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(G2072), .B(G33), .ZN(n916) );
  NOR2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(n918), .B(KEYINPUT120), .ZN(n919) );
  NAND2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(n925), .B(KEYINPUT53), .ZN(n928) );
  XOR2_X1 U1024 ( .A(G2084), .B(G34), .Z(n926) );
  XNOR2_X1 U1025 ( .A(KEYINPUT54), .B(n926), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n931) );
  XOR2_X1 U1027 ( .A(KEYINPUT119), .B(G2090), .Z(n929) );
  XNOR2_X1 U1028 ( .A(G35), .B(n929), .ZN(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n1015) );
  NAND2_X1 U1030 ( .A1(KEYINPUT55), .A2(n1015), .ZN(n932) );
  NAND2_X1 U1031 ( .A1(G11), .A2(n932), .ZN(n1014) );
  XNOR2_X1 U1032 ( .A(G164), .B(G2078), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(G2072), .B(n933), .ZN(n934) );
  XNOR2_X1 U1034 ( .A(n934), .B(KEYINPUT118), .ZN(n935) );
  NAND2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1036 ( .A(n937), .B(KEYINPUT50), .ZN(n950) );
  XOR2_X1 U1037 ( .A(G2090), .B(G162), .Z(n938) );
  NOR2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1039 ( .A(KEYINPUT51), .B(n940), .Z(n944) );
  NOR2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n946) );
  XOR2_X1 U1042 ( .A(G160), .B(G2084), .Z(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n952) );
  NAND2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(KEYINPUT52), .B(n955), .ZN(n957) );
  INV_X1 U1049 ( .A(KEYINPUT55), .ZN(n956) );
  NAND2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1051 ( .A1(n958), .A2(G29), .ZN(n1012) );
  XOR2_X1 U1052 ( .A(G1976), .B(G23), .Z(n961) );
  XOR2_X1 U1053 ( .A(G22), .B(KEYINPUT124), .Z(n959) );
  XNOR2_X1 U1054 ( .A(n959), .B(G1971), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n964) );
  XOR2_X1 U1056 ( .A(KEYINPUT125), .B(G1986), .Z(n962) );
  XNOR2_X1 U1057 ( .A(G24), .B(n962), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(KEYINPUT58), .B(n965), .ZN(n969) );
  XNOR2_X1 U1060 ( .A(G1966), .B(G21), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(G5), .B(G1961), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n980) );
  XNOR2_X1 U1064 ( .A(G1956), .B(G20), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(G1341), .B(G19), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(G1981), .B(G6), .ZN(n970) );
  NOR2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1068 ( .A(KEYINPUT123), .B(n972), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(G1348), .B(KEYINPUT59), .ZN(n975) );
  XNOR2_X1 U1071 ( .A(n975), .B(G4), .ZN(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(KEYINPUT60), .B(n978), .ZN(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1075 ( .A(n981), .B(KEYINPUT61), .Z(n982) );
  XNOR2_X1 U1076 ( .A(KEYINPUT126), .B(n982), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(G16), .A2(n983), .ZN(n1009) );
  XOR2_X1 U1078 ( .A(G16), .B(KEYINPUT56), .Z(n1007) );
  XNOR2_X1 U1079 ( .A(G1341), .B(KEYINPUT122), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(n985), .B(n984), .ZN(n987) );
  XOR2_X1 U1081 ( .A(G171), .B(G1961), .Z(n986) );
  NOR2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n997) );
  XOR2_X1 U1083 ( .A(G1348), .B(n988), .Z(n990) );
  NAND2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(G1966), .B(G168), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1087 ( .A(KEYINPUT57), .B(n993), .Z(n994) );
  NOR2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n1005) );
  NAND2_X1 U1090 ( .A1(G1971), .A2(G303), .ZN(n999) );
  XOR2_X1 U1091 ( .A(G1956), .B(G299), .Z(n998) );
  NAND2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1098 ( .A(KEYINPUT127), .B(n1010), .Z(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1019) );
  INV_X1 U1101 ( .A(n1015), .ZN(n1017) );
  NOR2_X1 U1102 ( .A1(G29), .A2(KEYINPUT55), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1020), .ZN(G150) );
  INV_X1 U1106 ( .A(G150), .ZN(G311) );
endmodule

