//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 0 0 1 1 1 0 1 0 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n597, new_n598, new_n599, new_n600, new_n601, new_n603,
    new_n604, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n783, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898;
  XOR2_X1   g000(.A(G15gat), .B(G22gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT90), .ZN(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n204), .A2(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n206), .B2(new_n203), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(G8gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT17), .ZN(new_n209));
  INV_X1    g008(.A(G29gat), .ZN(new_n210));
  AND3_X1   g009(.A1(new_n210), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT14), .B(G29gat), .ZN(new_n212));
  INV_X1    g011(.A(G36gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT15), .ZN(new_n215));
  INV_X1    g014(.A(G43gat), .ZN(new_n216));
  INV_X1    g015(.A(G50gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G43gat), .A2(G50gat), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n215), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(new_n221), .B(KEYINPUT88), .Z(new_n222));
  NOR2_X1   g021(.A1(new_n214), .A2(new_n220), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT89), .B(G50gat), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n215), .B(new_n219), .C1(new_n224), .C2(G43gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n208), .B1(new_n209), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n222), .A2(KEYINPUT17), .A3(new_n226), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n228), .A2(new_n229), .B1(new_n208), .B2(new_n227), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT18), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(KEYINPUT18), .A3(new_n231), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n208), .B(new_n227), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n231), .B(KEYINPUT13), .Z(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n234), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G113gat), .B(G141gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n240), .B(G197gat), .ZN(new_n241));
  XOR2_X1   g040(.A(KEYINPUT11), .B(G169gat), .Z(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g042(.A(new_n243), .B(KEYINPUT12), .Z(new_n244));
  NAND2_X1  g043(.A1(new_n239), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n244), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n234), .A2(new_n246), .A3(new_n235), .A4(new_n238), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G197gat), .B(G204gat), .ZN(new_n250));
  INV_X1    g049(.A(G211gat), .ZN(new_n251));
  INV_X1    g050(.A(G218gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n250), .B1(KEYINPUT22), .B2(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(G211gat), .B(G218gat), .Z(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT71), .ZN(new_n258));
  INV_X1    g057(.A(G183gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT27), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT27), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G183gat), .ZN(new_n262));
  INV_X1    g061(.A(G190gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n260), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  AND2_X1   g063(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G183gat), .A2(G190gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NOR3_X1   g067(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(G169gat), .A2(G176gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT26), .ZN(new_n271));
  NAND2_X1  g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n274));
  OAI22_X1  g073(.A1(new_n269), .A2(new_n273), .B1(new_n264), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n268), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT25), .ZN(new_n277));
  INV_X1    g076(.A(G169gat), .ZN(new_n278));
  INV_X1    g077(.A(G176gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n279), .A3(KEYINPUT23), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT23), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n281), .B1(G169gat), .B2(G176gat), .ZN(new_n282));
  AND3_X1   g081(.A1(new_n280), .A2(new_n282), .A3(new_n272), .ZN(new_n283));
  NOR2_X1   g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n267), .A2(KEYINPUT24), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT24), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n286), .A2(G183gat), .A3(G190gat), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n284), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n283), .B1(new_n288), .B2(KEYINPUT64), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT64), .ZN(new_n290));
  AOI211_X1 g089(.A(new_n290), .B(new_n284), .C1(new_n285), .C2(new_n287), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n277), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n280), .A2(new_n282), .A3(KEYINPUT25), .A4(new_n272), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT65), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n284), .B(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n285), .A2(new_n287), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n276), .B1(new_n292), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G226gat), .A2(G233gat), .ZN(new_n300));
  XOR2_X1   g099(.A(new_n300), .B(KEYINPUT69), .Z(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n258), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n285), .A2(new_n287), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n290), .B1(new_n304), .B2(new_n284), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n288), .A2(KEYINPUT64), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(new_n306), .A3(new_n283), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n297), .B1(new_n307), .B2(new_n277), .ZN(new_n308));
  OAI211_X1 g107(.A(KEYINPUT71), .B(new_n301), .C1(new_n308), .C2(new_n276), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n257), .B1(new_n303), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT70), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(new_n308), .B2(new_n276), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n312), .B1(new_n314), .B2(new_n300), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n312), .B(new_n300), .C1(new_n299), .C2(KEYINPUT29), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n310), .B(new_n311), .C1(new_n315), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n314), .A2(new_n302), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n319), .B1(new_n299), .B2(new_n300), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(new_n257), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n300), .B1(new_n299), .B2(KEYINPUT29), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT70), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n316), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n311), .B1(new_n325), .B2(new_n310), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n328));
  XNOR2_X1  g127(.A(G8gat), .B(G36gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(G64gat), .B(G92gat), .ZN(new_n330));
  XOR2_X1   g129(.A(new_n329), .B(new_n330), .Z(new_n331));
  NAND4_X1  g130(.A1(new_n327), .A2(new_n328), .A3(KEYINPUT30), .A4(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n331), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n333), .B1(new_n322), .B2(new_n326), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT73), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT30), .ZN(new_n336));
  NOR4_X1   g135(.A1(new_n322), .A2(new_n326), .A3(new_n336), .A4(new_n333), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n332), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n327), .A2(new_n331), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n336), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT85), .ZN(new_n342));
  INV_X1    g141(.A(G22gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(G228gat), .A2(G233gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(KEYINPUT84), .ZN(new_n345));
  NAND2_X1  g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346));
  INV_X1    g145(.A(G155gat), .ZN(new_n347));
  INV_X1    g146(.A(G162gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n346), .B1(new_n349), .B2(KEYINPUT2), .ZN(new_n350));
  INV_X1    g149(.A(G141gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT75), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G141gat), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n352), .A2(new_n354), .A3(G148gat), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT76), .B1(new_n351), .B2(G148gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n357));
  INV_X1    g156(.A(G148gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n358), .A3(G141gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n350), .B1(new_n355), .B2(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G141gat), .B(G148gat), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n346), .B(new_n349), .C1(new_n362), .C2(KEYINPUT2), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n256), .A2(new_n313), .ZN(new_n365));
  XOR2_X1   g164(.A(KEYINPUT77), .B(KEYINPUT3), .Z(new_n366));
  AOI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n361), .A2(new_n363), .A3(new_n366), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n256), .B1(new_n313), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n345), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT3), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n371), .B1(new_n361), .B2(new_n363), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n372), .A2(new_n344), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n368), .A2(new_n313), .ZN(new_n374));
  OAI221_X1 g173(.A(new_n373), .B1(new_n365), .B2(new_n364), .C1(new_n374), .C2(new_n256), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G78gat), .B(G106gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(new_n217), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT83), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n380), .B(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n342), .B(new_n343), .C1(new_n376), .C2(new_n383), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n376), .A2(new_n383), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n383), .B1(new_n370), .B2(new_n375), .ZN(new_n386));
  OAI21_X1  g185(.A(G22gat), .B1(new_n386), .B2(KEYINPUT85), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n385), .B1(new_n384), .B2(new_n387), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G113gat), .B(G120gat), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT1), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT67), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G127gat), .B(G134gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n395), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(new_n391), .B2(new_n393), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n299), .B(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(G227gat), .ZN(new_n401));
  INV_X1    g200(.A(G233gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(KEYINPUT34), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT32), .B1(new_n400), .B2(new_n404), .ZN(new_n408));
  XOR2_X1   g207(.A(G71gat), .B(G99gat), .Z(new_n409));
  XNOR2_X1  g208(.A(G15gat), .B(G43gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n400), .A2(new_n404), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n408), .B(new_n411), .C1(new_n412), .C2(KEYINPUT33), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT68), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT32), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n396), .A2(new_n398), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n299), .B(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n417), .B2(new_n403), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n411), .A2(KEYINPUT33), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n414), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n418), .A2(new_n414), .A3(new_n419), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n407), .B(new_n413), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n413), .B1(new_n421), .B2(new_n420), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n406), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n390), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G1gat), .B(G29gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT0), .ZN(new_n427));
  XNOR2_X1  g226(.A(G57gat), .B(G85gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  NAND3_X1  g228(.A1(new_n364), .A2(new_n416), .A3(KEYINPUT4), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n361), .A2(new_n396), .A3(new_n398), .A4(new_n363), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT4), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n368), .A2(new_n399), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT78), .B1(new_n435), .B2(new_n372), .ZN(new_n436));
  INV_X1    g235(.A(new_n372), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT78), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n437), .A2(new_n438), .A3(new_n368), .A4(new_n399), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n434), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(G225gat), .A2(G233gat), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(KEYINPUT5), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n361), .A2(new_n363), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n399), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n445), .A2(KEYINPUT79), .A3(new_n431), .ZN(new_n446));
  INV_X1    g245(.A(new_n441), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT79), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n444), .A2(new_n399), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n440), .A2(new_n441), .B1(KEYINPUT5), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n429), .B1(new_n443), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n440), .A2(new_n441), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(KEYINPUT5), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n429), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(new_n456), .A3(new_n442), .ZN(new_n457));
  XOR2_X1   g256(.A(KEYINPUT80), .B(KEYINPUT6), .Z(new_n458));
  NAND3_X1  g257(.A1(new_n452), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n457), .A2(new_n458), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n462), .A2(KEYINPUT35), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n341), .A2(new_n425), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT74), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n338), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n332), .B(KEYINPUT74), .C1(new_n335), .C2(new_n337), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT81), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n461), .B1(new_n459), .B2(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n452), .A2(new_n457), .A3(KEYINPUT81), .A4(new_n458), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n469), .A2(new_n470), .B1(new_n336), .B2(new_n339), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n466), .A2(new_n425), .A3(new_n467), .A4(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT87), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n472), .A2(new_n473), .A3(KEYINPUT35), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n473), .B1(new_n472), .B2(KEYINPUT35), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n464), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT37), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n331), .B1(new_n327), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n477), .B1(new_n320), .B2(new_n256), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n256), .B1(new_n303), .B2(new_n309), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n325), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT38), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n483), .A2(new_n462), .A3(new_n339), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT38), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT37), .B1(new_n322), .B2(new_n326), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n485), .B1(new_n478), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n440), .A2(new_n441), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT39), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n447), .B1(new_n446), .B2(new_n449), .ZN(new_n490));
  OR3_X1    g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n456), .B1(new_n488), .B2(new_n489), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n493), .A2(KEYINPUT40), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(KEYINPUT40), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n457), .A3(new_n495), .ZN(new_n496));
  OAI221_X1 g295(.A(new_n390), .B1(new_n484), .B2(new_n487), .C1(new_n341), .C2(new_n496), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n422), .A2(new_n424), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(KEYINPUT36), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n466), .A2(new_n467), .A3(new_n471), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n390), .B(KEYINPUT86), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n497), .B(new_n499), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n249), .B1(new_n476), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n469), .A2(new_n470), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n227), .A2(new_n209), .ZN(new_n506));
  NAND2_X1  g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507));
  INV_X1    g306(.A(G85gat), .ZN(new_n508));
  INV_X1    g307(.A(G92gat), .ZN(new_n509));
  AOI22_X1  g308(.A1(KEYINPUT8), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT96), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT7), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n512), .A2(KEYINPUT94), .ZN(new_n513));
  NAND2_X1  g312(.A1(G85gat), .A2(G92gat), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n512), .B1(new_n514), .B2(KEYINPUT94), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT95), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n516), .A2(G85gat), .A3(G92gat), .ZN(new_n517));
  MUX2_X1   g316(.A(new_n513), .B(new_n515), .S(new_n517), .Z(new_n518));
  NAND2_X1  g317(.A1(new_n511), .A2(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(G99gat), .B(G106gat), .Z(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n506), .A2(new_n229), .A3(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n522), .B(KEYINPUT97), .Z(new_n523));
  INV_X1    g322(.A(new_n521), .ZN(new_n524));
  AND2_X1   g323(.A1(G232gat), .A2(G233gat), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n524), .A2(new_n227), .B1(KEYINPUT41), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G190gat), .B(G218gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT98), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n527), .A2(new_n529), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n525), .A2(KEYINPUT41), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT93), .ZN(new_n534));
  XNOR2_X1  g333(.A(G134gat), .B(G162gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n530), .A2(new_n536), .A3(new_n531), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OR2_X1    g339(.A1(G57gat), .A2(G64gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(G57gat), .A2(G64gat), .ZN(new_n542));
  AND2_X1   g341(.A1(G71gat), .A2(G78gat), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n541), .B(new_n542), .C1(new_n543), .C2(KEYINPUT9), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT91), .B1(G71gat), .B2(G78gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G71gat), .B(G78gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT21), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G231gat), .A2(G233gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(G127gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n548), .B(KEYINPUT92), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n208), .B1(new_n555), .B2(KEYINPUT21), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n554), .B(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(new_n347), .ZN(new_n559));
  XOR2_X1   g358(.A(G183gat), .B(G211gat), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n557), .B(new_n561), .ZN(new_n562));
  OR3_X1    g361(.A1(new_n540), .A2(KEYINPUT99), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT99), .B1(new_n540), .B2(new_n562), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n519), .A2(new_n520), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT100), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n548), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(new_n521), .ZN(new_n568));
  NAND2_X1  g367(.A1(G230gat), .A2(G233gat), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n570), .B(KEYINPUT101), .Z(new_n571));
  INV_X1    g370(.A(KEYINPUT10), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n524), .A2(new_n555), .A3(KEYINPUT10), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n569), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G120gat), .B(G148gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(G176gat), .B(G204gat), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n578), .B(new_n579), .Z(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n577), .A2(new_n581), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n563), .A2(new_n564), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n503), .A2(new_n505), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(G1gat), .ZN(G1324gat));
  INV_X1    g388(.A(new_n341), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n503), .A2(new_n590), .A3(new_n587), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n591), .A2(G8gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT16), .B(G8gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT42), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n595), .B1(KEYINPUT42), .B2(new_n594), .ZN(G1325gat));
  NAND2_X1  g395(.A1(new_n503), .A2(new_n587), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n499), .B(KEYINPUT102), .Z(new_n598));
  OAI21_X1  g397(.A(G15gat), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n498), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n600), .A2(G15gat), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n599), .B1(new_n597), .B2(new_n601), .ZN(G1326gat));
  NOR2_X1   g401(.A1(new_n597), .A2(new_n501), .ZN(new_n603));
  XOR2_X1   g402(.A(KEYINPUT43), .B(G22gat), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(G1327gat));
  INV_X1    g404(.A(new_n540), .ZN(new_n606));
  INV_X1    g405(.A(new_n562), .ZN(new_n607));
  NOR3_X1   g406(.A1(new_n606), .A2(new_n607), .A3(new_n585), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n503), .A2(new_n608), .ZN(new_n609));
  NOR3_X1   g408(.A1(new_n609), .A2(G29gat), .A3(new_n504), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(KEYINPUT45), .Z(new_n611));
  INV_X1    g410(.A(new_n502), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT105), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n476), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g413(.A(KEYINPUT105), .B(new_n464), .C1(new_n474), .C2(new_n475), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(KEYINPUT106), .B1(new_n538), .B2(new_n539), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n538), .A2(KEYINPUT106), .A3(new_n539), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(KEYINPUT44), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT44), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n606), .B1(new_n476), .B2(new_n502), .ZN(new_n624));
  OAI22_X1  g423(.A1(new_n616), .A2(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n562), .B(KEYINPUT104), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n245), .A2(KEYINPUT103), .A3(new_n247), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT103), .B1(new_n245), .B2(new_n247), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n627), .A2(new_n631), .A3(new_n585), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n625), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(G29gat), .B1(new_n633), .B2(new_n504), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n611), .A2(new_n634), .ZN(G1328gat));
  NOR3_X1   g434(.A1(new_n609), .A2(G36gat), .A3(new_n341), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT46), .ZN(new_n637));
  OAI21_X1  g436(.A(G36gat), .B1(new_n633), .B2(new_n341), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(G1329gat));
  NOR3_X1   g438(.A1(new_n609), .A2(G43gat), .A3(new_n600), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT108), .ZN(new_n641));
  OAI21_X1  g440(.A(G43gat), .B1(new_n633), .B2(new_n499), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n641), .A2(new_n642), .A3(KEYINPUT47), .ZN(new_n643));
  INV_X1    g442(.A(new_n598), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n625), .A2(new_n644), .A3(new_n632), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(G43gat), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT107), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT107), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n645), .A2(new_n648), .A3(G43gat), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n647), .A2(new_n649), .A3(new_n641), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n643), .B1(new_n650), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g450(.A(new_n224), .B1(new_n633), .B2(new_n390), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n609), .A2(new_n501), .A3(new_n224), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n652), .A2(KEYINPUT48), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n501), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n625), .A2(new_n656), .A3(new_n632), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n653), .B1(new_n657), .B2(new_n224), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n659));
  OAI21_X1  g458(.A(new_n655), .B1(new_n658), .B2(new_n659), .ZN(G1331gat));
  NAND2_X1  g459(.A1(new_n563), .A2(new_n564), .ZN(new_n661));
  NOR4_X1   g460(.A1(new_n616), .A2(new_n661), .A3(new_n586), .A4(new_n630), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n505), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n590), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n665), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT49), .B(G64gat), .Z(new_n667));
  OAI21_X1  g466(.A(new_n666), .B1(new_n665), .B2(new_n667), .ZN(G1333gat));
  NAND2_X1  g467(.A1(new_n662), .A2(new_n644), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n600), .A2(G71gat), .ZN(new_n670));
  AOI22_X1  g469(.A1(new_n669), .A2(G71gat), .B1(new_n662), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g471(.A1(new_n662), .A2(new_n656), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT110), .B(G78gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1335gat));
  INV_X1    g474(.A(KEYINPUT112), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n476), .A2(new_n502), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n623), .B1(new_n677), .B2(new_n540), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n472), .A2(KEYINPUT35), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT87), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n472), .A2(new_n473), .A3(KEYINPUT35), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT105), .B1(new_n682), .B2(new_n464), .ZN(new_n683));
  INV_X1    g482(.A(new_n615), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n502), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n678), .B1(new_n685), .B2(new_n621), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n631), .A2(new_n562), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n586), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT111), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT111), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n625), .A2(new_n691), .A3(new_n688), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n676), .B1(new_n693), .B2(new_n504), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G85gat), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n693), .A2(new_n676), .A3(new_n504), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n631), .A2(new_n562), .A3(new_n540), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n616), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT51), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n585), .A2(new_n508), .A3(new_n505), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT113), .ZN(new_n702));
  OAI22_X1  g501(.A1(new_n695), .A2(new_n696), .B1(new_n700), .B2(new_n702), .ZN(G1336gat));
  NAND3_X1  g502(.A1(new_n690), .A2(new_n590), .A3(new_n692), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(G92gat), .ZN(new_n705));
  INV_X1    g504(.A(new_n697), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n685), .A2(KEYINPUT114), .A3(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT114), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n708), .B1(new_n616), .B2(new_n697), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n707), .A2(new_n709), .A3(new_n699), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT115), .B1(new_n698), .B2(KEYINPUT51), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n586), .A2(G92gat), .A3(new_n341), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n707), .A2(new_n709), .A3(KEYINPUT115), .A4(new_n699), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n705), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT52), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n698), .B(KEYINPUT51), .ZN(new_n718));
  AOI21_X1  g517(.A(KEYINPUT52), .B1(new_n718), .B2(new_n713), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n686), .A2(new_n341), .A3(new_n689), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n719), .B1(new_n509), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n717), .A2(new_n721), .ZN(G1337gat));
  OAI21_X1  g521(.A(G99gat), .B1(new_n693), .B2(new_n598), .ZN(new_n723));
  OR3_X1    g522(.A1(new_n586), .A2(G99gat), .A3(new_n600), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n723), .B1(new_n700), .B2(new_n724), .ZN(G1338gat));
  INV_X1    g524(.A(new_n390), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n625), .A2(new_n726), .A3(new_n688), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT116), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n625), .A2(KEYINPUT116), .A3(new_n726), .A4(new_n688), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n729), .A2(G106gat), .A3(new_n730), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n586), .A2(G106gat), .A3(new_n390), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n718), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT53), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n712), .A2(new_n714), .A3(new_n732), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n735), .A2(KEYINPUT53), .ZN(new_n736));
  OAI21_X1  g535(.A(G106gat), .B1(new_n693), .B2(new_n501), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(G1339gat));
  INV_X1    g537(.A(KEYINPUT118), .ZN(new_n739));
  OR2_X1    g538(.A1(new_n575), .A2(new_n569), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n740), .A2(KEYINPUT54), .A3(new_n576), .ZN(new_n741));
  OR2_X1    g540(.A1(new_n576), .A2(KEYINPUT54), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n741), .A2(new_n742), .A3(KEYINPUT55), .A4(new_n581), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT117), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n741), .A2(new_n581), .A3(new_n742), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT55), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n582), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n538), .A2(KEYINPUT106), .A3(new_n539), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(new_n617), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n230), .A2(new_n231), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n236), .A2(new_n237), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n243), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n247), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n749), .A2(new_n751), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n630), .A2(new_n745), .A3(new_n748), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n585), .A2(new_n755), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n739), .B(new_n756), .C1(new_n759), .C2(new_n751), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n751), .B1(new_n757), .B2(new_n758), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n748), .A3(new_n755), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n620), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT118), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n760), .A2(new_n764), .A3(new_n626), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n587), .A2(new_n631), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n504), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n425), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n590), .A2(new_n768), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(G113gat), .B1(new_n770), .B2(new_n630), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n656), .B1(new_n765), .B2(new_n766), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n590), .A2(new_n600), .A3(new_n504), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(G113gat), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n774), .A2(new_n775), .A3(new_n249), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n771), .A2(new_n776), .ZN(G1340gat));
  NOR2_X1   g576(.A1(new_n586), .A2(G120gat), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n778), .B(KEYINPUT119), .Z(new_n779));
  NAND2_X1  g578(.A1(new_n770), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(G120gat), .B1(new_n774), .B2(new_n586), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(G1341gat));
  NAND3_X1  g581(.A1(new_n770), .A2(new_n553), .A3(new_n607), .ZN(new_n783));
  OAI21_X1  g582(.A(G127gat), .B1(new_n774), .B2(new_n626), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1342gat));
  INV_X1    g584(.A(KEYINPUT56), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n606), .A2(G134gat), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n770), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT120), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n770), .A2(KEYINPUT120), .A3(new_n786), .A4(new_n787), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n786), .B1(new_n770), .B2(new_n787), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n772), .A2(new_n540), .A3(new_n773), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n793), .B1(G134gat), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n792), .A2(new_n795), .ZN(G1343gat));
  AOI21_X1  g595(.A(new_n390), .B1(new_n765), .B2(new_n766), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n499), .A2(new_n505), .A3(new_n341), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n745), .A2(new_n748), .A3(new_n248), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n540), .B1(new_n801), .B2(new_n758), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n562), .B1(new_n802), .B2(new_n763), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n766), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n656), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n800), .B1(new_n805), .B2(KEYINPUT57), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n799), .A2(new_n806), .ZN(new_n807));
  AOI22_X1  g606(.A1(new_n807), .A2(new_n248), .B1(new_n352), .B2(new_n354), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n598), .A2(new_n726), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT121), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n341), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n810), .B2(new_n809), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n767), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n249), .A2(G141gat), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT58), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n799), .A2(new_n630), .A3(new_n806), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n352), .A2(new_n354), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n818), .A2(new_n819), .B1(new_n813), .B2(new_n814), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n808), .A2(new_n817), .B1(new_n820), .B2(new_n816), .ZN(G1344gat));
  NAND3_X1  g620(.A1(new_n813), .A2(new_n358), .A3(new_n585), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT59), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G148gat), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n824), .B1(new_n807), .B2(new_n585), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n762), .A2(new_n606), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n562), .B1(new_n802), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n587), .A2(new_n249), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n829), .A2(new_n798), .A3(new_n656), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n800), .A2(new_n586), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n830), .B(new_n831), .C1(new_n797), .C2(new_n798), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n823), .B1(new_n832), .B2(G148gat), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n822), .B1(new_n825), .B2(new_n833), .ZN(G1345gat));
  NAND3_X1  g633(.A1(new_n813), .A2(new_n347), .A3(new_n607), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n807), .A2(new_n627), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(new_n347), .ZN(G1346gat));
  AOI21_X1  g636(.A(G162gat), .B1(new_n813), .B2(new_n540), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n620), .A2(new_n348), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n807), .B2(new_n839), .ZN(G1347gat));
  NAND2_X1  g639(.A1(new_n765), .A2(new_n766), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n341), .A2(new_n505), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n768), .ZN(new_n844));
  AOI21_X1  g643(.A(G169gat), .B1(new_n844), .B2(new_n630), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n842), .A2(new_n498), .ZN(new_n846));
  AOI211_X1 g645(.A(new_n656), .B(new_n846), .C1(new_n765), .C2(new_n766), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n249), .A2(new_n278), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(G1348gat));
  NAND3_X1  g648(.A1(new_n847), .A2(G176gat), .A3(new_n585), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT122), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  AOI21_X1  g652(.A(G176gat), .B1(new_n844), .B2(new_n585), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(G1349gat));
  NAND2_X1  g654(.A1(new_n260), .A2(new_n262), .ZN(new_n856));
  NOR4_X1   g655(.A1(new_n843), .A2(new_n856), .A3(new_n768), .A4(new_n562), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n259), .B1(new_n847), .B2(new_n627), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n859), .A2(KEYINPUT60), .ZN(new_n860));
  OR3_X1    g659(.A1(new_n857), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n860), .B1(new_n857), .B2(new_n858), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1350gat));
  NAND3_X1  g662(.A1(new_n844), .A2(new_n263), .A3(new_n751), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT61), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n847), .A2(new_n540), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n865), .B1(new_n866), .B2(G190gat), .ZN(new_n867));
  AOI211_X1 g666(.A(KEYINPUT61), .B(new_n263), .C1(new_n847), .C2(new_n540), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n864), .B1(new_n867), .B2(new_n868), .ZN(G1351gat));
  AND2_X1   g668(.A1(new_n598), .A2(new_n842), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n830), .B(new_n870), .C1(new_n797), .C2(new_n798), .ZN(new_n871));
  OAI21_X1  g670(.A(G197gat), .B1(new_n871), .B2(new_n249), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n843), .A2(new_n809), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n631), .A2(G197gat), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n873), .A2(KEYINPUT124), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT124), .B1(new_n873), .B2(new_n874), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n872), .B1(new_n875), .B2(new_n876), .ZN(G1352gat));
  INV_X1    g676(.A(new_n809), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n586), .A2(G204gat), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n841), .A2(new_n878), .A3(new_n842), .A4(new_n879), .ZN(new_n880));
  XOR2_X1   g679(.A(new_n880), .B(KEYINPUT62), .Z(new_n881));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n882), .B1(new_n871), .B2(new_n586), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(G204gat), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n871), .A2(new_n882), .A3(new_n586), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n881), .B1(new_n884), .B2(new_n885), .ZN(G1353gat));
  OAI21_X1  g685(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(new_n871), .B2(new_n562), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(KEYINPUT127), .A3(KEYINPUT63), .ZN(new_n890));
  NAND2_X1  g689(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n891), .B(new_n888), .C1(new_n871), .C2(new_n562), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n562), .A2(G211gat), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n841), .A2(new_n878), .A3(new_n842), .A4(new_n893), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT126), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n890), .A2(new_n892), .A3(new_n895), .ZN(G1354gat));
  OAI21_X1  g695(.A(G218gat), .B1(new_n871), .B2(new_n606), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n873), .A2(new_n252), .A3(new_n751), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1355gat));
endmodule


