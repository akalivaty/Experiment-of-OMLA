

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U548 ( .A1(G8), .A2(n677), .ZN(n717) );
  NAND2_X1 U549 ( .A1(n622), .A2(n621), .ZN(n677) );
  NOR2_X4 U550 ( .A1(n519), .A2(G2105), .ZN(n879) );
  NOR2_X1 U551 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U552 ( .A1(G1966), .A2(n717), .ZN(n693) );
  NOR2_X1 U553 ( .A1(n724), .A2(n723), .ZN(n726) );
  NAND2_X1 U554 ( .A1(n879), .A2(G101), .ZN(n514) );
  INV_X1 U555 ( .A(KEYINPUT29), .ZN(n673) );
  XNOR2_X1 U556 ( .A(n674), .B(n673), .ZN(n675) );
  AND2_X1 U557 ( .A1(n690), .A2(n685), .ZN(n684) );
  INV_X1 U558 ( .A(KEYINPUT101), .ZN(n725) );
  NOR2_X1 U559 ( .A1(G2105), .A2(G2104), .ZN(n516) );
  NOR2_X1 U560 ( .A1(G651), .A2(n570), .ZN(n784) );
  NOR2_X1 U561 ( .A1(n524), .A2(n523), .ZN(G160) );
  INV_X1 U562 ( .A(G2104), .ZN(n519) );
  XOR2_X1 U563 ( .A(KEYINPUT64), .B(n514), .Z(n515) );
  XNOR2_X1 U564 ( .A(n515), .B(KEYINPUT23), .ZN(n518) );
  XOR2_X1 U565 ( .A(KEYINPUT17), .B(n516), .Z(n880) );
  NAND2_X1 U566 ( .A1(G137), .A2(n880), .ZN(n517) );
  NAND2_X1 U567 ( .A1(n518), .A2(n517), .ZN(n524) );
  INV_X1 U568 ( .A(G2105), .ZN(n520) );
  NOR2_X1 U569 ( .A1(G2104), .A2(n520), .ZN(n875) );
  NAND2_X1 U570 ( .A1(G125), .A2(n875), .ZN(n522) );
  NOR2_X1 U571 ( .A1(n520), .A2(n519), .ZN(n876) );
  NAND2_X1 U572 ( .A1(G113), .A2(n876), .ZN(n521) );
  NAND2_X1 U573 ( .A1(n522), .A2(n521), .ZN(n523) );
  NAND2_X1 U574 ( .A1(n880), .A2(G138), .ZN(n527) );
  NAND2_X1 U575 ( .A1(G102), .A2(n879), .ZN(n525) );
  XOR2_X1 U576 ( .A(KEYINPUT91), .B(n525), .Z(n526) );
  NAND2_X1 U577 ( .A1(n527), .A2(n526), .ZN(n531) );
  NAND2_X1 U578 ( .A1(G126), .A2(n875), .ZN(n529) );
  NAND2_X1 U579 ( .A1(G114), .A2(n876), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U581 ( .A1(n531), .A2(n530), .ZN(G164) );
  XOR2_X1 U582 ( .A(KEYINPUT0), .B(G543), .Z(n570) );
  INV_X1 U583 ( .A(G651), .ZN(n537) );
  NOR2_X1 U584 ( .A1(n570), .A2(n537), .ZN(n788) );
  NAND2_X1 U585 ( .A1(G77), .A2(n788), .ZN(n533) );
  NOR2_X1 U586 ( .A1(G651), .A2(G543), .ZN(n789) );
  NAND2_X1 U587 ( .A1(G90), .A2(n789), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U589 ( .A(n534), .B(KEYINPUT9), .ZN(n536) );
  NAND2_X1 U590 ( .A1(G52), .A2(n784), .ZN(n535) );
  NAND2_X1 U591 ( .A1(n536), .A2(n535), .ZN(n542) );
  NOR2_X1 U592 ( .A1(G543), .A2(n537), .ZN(n538) );
  XOR2_X1 U593 ( .A(KEYINPUT66), .B(n538), .Z(n539) );
  XNOR2_X1 U594 ( .A(KEYINPUT1), .B(n539), .ZN(n785) );
  NAND2_X1 U595 ( .A1(G64), .A2(n785), .ZN(n540) );
  XNOR2_X1 U596 ( .A(KEYINPUT67), .B(n540), .ZN(n541) );
  NOR2_X1 U597 ( .A1(n542), .A2(n541), .ZN(G171) );
  NAND2_X1 U598 ( .A1(n788), .A2(G76), .ZN(n543) );
  XNOR2_X1 U599 ( .A(KEYINPUT74), .B(n543), .ZN(n546) );
  NAND2_X1 U600 ( .A1(n789), .A2(G89), .ZN(n544) );
  XNOR2_X1 U601 ( .A(KEYINPUT4), .B(n544), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U603 ( .A(KEYINPUT5), .B(n547), .ZN(n554) );
  XNOR2_X1 U604 ( .A(KEYINPUT76), .B(KEYINPUT6), .ZN(n552) );
  NAND2_X1 U605 ( .A1(n784), .A2(G51), .ZN(n550) );
  NAND2_X1 U606 ( .A1(G63), .A2(n785), .ZN(n548) );
  XOR2_X1 U607 ( .A(KEYINPUT75), .B(n548), .Z(n549) );
  NAND2_X1 U608 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U609 ( .A(n552), .B(n551), .Z(n553) );
  NAND2_X1 U610 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U611 ( .A(KEYINPUT7), .B(n555), .ZN(G168) );
  NAND2_X1 U612 ( .A1(n784), .A2(G53), .ZN(n557) );
  NAND2_X1 U613 ( .A1(G65), .A2(n785), .ZN(n556) );
  NAND2_X1 U614 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U615 ( .A(KEYINPUT68), .B(n558), .Z(n562) );
  NAND2_X1 U616 ( .A1(n788), .A2(G78), .ZN(n560) );
  NAND2_X1 U617 ( .A1(G91), .A2(n789), .ZN(n559) );
  AND2_X1 U618 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U619 ( .A1(n562), .A2(n561), .ZN(G299) );
  NAND2_X1 U620 ( .A1(n784), .A2(G50), .ZN(n564) );
  NAND2_X1 U621 ( .A1(G62), .A2(n785), .ZN(n563) );
  NAND2_X1 U622 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U623 ( .A1(G75), .A2(n788), .ZN(n566) );
  NAND2_X1 U624 ( .A1(G88), .A2(n789), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U626 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U627 ( .A(n569), .B(KEYINPUT83), .ZN(G303) );
  XOR2_X1 U628 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U629 ( .A1(G87), .A2(n570), .ZN(n572) );
  NAND2_X1 U630 ( .A1(G74), .A2(G651), .ZN(n571) );
  NAND2_X1 U631 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U632 ( .A1(n785), .A2(n573), .ZN(n576) );
  NAND2_X1 U633 ( .A1(G49), .A2(n784), .ZN(n574) );
  XOR2_X1 U634 ( .A(KEYINPUT81), .B(n574), .Z(n575) );
  NAND2_X1 U635 ( .A1(n576), .A2(n575), .ZN(G288) );
  NAND2_X1 U636 ( .A1(G86), .A2(n789), .ZN(n578) );
  NAND2_X1 U637 ( .A1(G61), .A2(n785), .ZN(n577) );
  NAND2_X1 U638 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U639 ( .A(KEYINPUT82), .B(n579), .ZN(n582) );
  NAND2_X1 U640 ( .A1(n788), .A2(G73), .ZN(n580) );
  XOR2_X1 U641 ( .A(KEYINPUT2), .B(n580), .Z(n581) );
  NOR2_X1 U642 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U643 ( .A1(n784), .A2(G48), .ZN(n583) );
  NAND2_X1 U644 ( .A1(n584), .A2(n583), .ZN(G305) );
  NAND2_X1 U645 ( .A1(G85), .A2(n789), .ZN(n586) );
  NAND2_X1 U646 ( .A1(G60), .A2(n785), .ZN(n585) );
  NAND2_X1 U647 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U648 ( .A1(G72), .A2(n788), .ZN(n587) );
  XNOR2_X1 U649 ( .A(KEYINPUT65), .B(n587), .ZN(n588) );
  NOR2_X1 U650 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U651 ( .A1(n784), .A2(G47), .ZN(n590) );
  NAND2_X1 U652 ( .A1(n591), .A2(n590), .ZN(G290) );
  NAND2_X1 U653 ( .A1(G141), .A2(n880), .ZN(n593) );
  NAND2_X1 U654 ( .A1(G117), .A2(n876), .ZN(n592) );
  NAND2_X1 U655 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U656 ( .A1(n879), .A2(G105), .ZN(n594) );
  XOR2_X1 U657 ( .A(KEYINPUT38), .B(n594), .Z(n595) );
  NOR2_X1 U658 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U659 ( .A1(n875), .A2(G129), .ZN(n597) );
  NAND2_X1 U660 ( .A1(n598), .A2(n597), .ZN(n857) );
  AND2_X1 U661 ( .A1(n857), .A2(G1996), .ZN(n606) );
  NAND2_X1 U662 ( .A1(G95), .A2(n879), .ZN(n600) );
  NAND2_X1 U663 ( .A1(G131), .A2(n880), .ZN(n599) );
  NAND2_X1 U664 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U665 ( .A1(G119), .A2(n875), .ZN(n602) );
  NAND2_X1 U666 ( .A1(G107), .A2(n876), .ZN(n601) );
  NAND2_X1 U667 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U668 ( .A1(n604), .A2(n603), .ZN(n870) );
  INV_X1 U669 ( .A(G1991), .ZN(n729) );
  NOR2_X1 U670 ( .A1(n870), .A2(n729), .ZN(n605) );
  NOR2_X1 U671 ( .A1(n606), .A2(n605), .ZN(n987) );
  NOR2_X1 U672 ( .A1(G164), .A2(G1384), .ZN(n622) );
  NAND2_X1 U673 ( .A1(G160), .A2(G40), .ZN(n620) );
  NOR2_X1 U674 ( .A1(n622), .A2(n620), .ZN(n740) );
  INV_X1 U675 ( .A(n740), .ZN(n607) );
  NOR2_X1 U676 ( .A1(n987), .A2(n607), .ZN(n732) );
  INV_X1 U677 ( .A(n732), .ZN(n619) );
  XNOR2_X1 U678 ( .A(G2067), .B(KEYINPUT37), .ZN(n737) );
  NAND2_X1 U679 ( .A1(G104), .A2(n879), .ZN(n609) );
  NAND2_X1 U680 ( .A1(G140), .A2(n880), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U682 ( .A(KEYINPUT34), .B(n610), .ZN(n617) );
  NAND2_X1 U683 ( .A1(n875), .A2(G128), .ZN(n611) );
  XNOR2_X1 U684 ( .A(n611), .B(KEYINPUT92), .ZN(n613) );
  NAND2_X1 U685 ( .A1(G116), .A2(n876), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U687 ( .A(KEYINPUT93), .B(n614), .ZN(n615) );
  XNOR2_X1 U688 ( .A(KEYINPUT35), .B(n615), .ZN(n616) );
  NOR2_X1 U689 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U690 ( .A(KEYINPUT36), .B(n618), .ZN(n890) );
  NOR2_X1 U691 ( .A1(n737), .A2(n890), .ZN(n1003) );
  NAND2_X1 U692 ( .A1(n740), .A2(n1003), .ZN(n735) );
  NAND2_X1 U693 ( .A1(n619), .A2(n735), .ZN(n724) );
  XOR2_X1 U694 ( .A(KEYINPUT94), .B(n620), .Z(n621) );
  INV_X1 U695 ( .A(n677), .ZN(n660) );
  XOR2_X1 U696 ( .A(G1961), .B(KEYINPUT96), .Z(n954) );
  NOR2_X1 U697 ( .A1(n660), .A2(n954), .ZN(n624) );
  XNOR2_X1 U698 ( .A(G2078), .B(KEYINPUT25), .ZN(n912) );
  NOR2_X1 U699 ( .A1(n677), .A2(n912), .ZN(n623) );
  NOR2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n632) );
  NOR2_X1 U701 ( .A1(G171), .A2(n632), .ZN(n629) );
  NOR2_X1 U702 ( .A1(G2084), .A2(n677), .ZN(n692) );
  NOR2_X1 U703 ( .A1(n693), .A2(n692), .ZN(n625) );
  NAND2_X1 U704 ( .A1(G8), .A2(n625), .ZN(n626) );
  XNOR2_X1 U705 ( .A(KEYINPUT30), .B(n626), .ZN(n627) );
  NOR2_X1 U706 ( .A1(G168), .A2(n627), .ZN(n628) );
  XNOR2_X1 U707 ( .A(n630), .B(KEYINPUT31), .ZN(n631) );
  XNOR2_X1 U708 ( .A(n631), .B(KEYINPUT99), .ZN(n691) );
  NAND2_X1 U709 ( .A1(G171), .A2(n632), .ZN(n676) );
  NAND2_X1 U710 ( .A1(n660), .A2(G2072), .ZN(n633) );
  XNOR2_X1 U711 ( .A(n633), .B(KEYINPUT27), .ZN(n635) );
  XNOR2_X1 U712 ( .A(G1956), .B(KEYINPUT97), .ZN(n956) );
  NOR2_X1 U713 ( .A1(n956), .A2(n660), .ZN(n634) );
  NOR2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n668) );
  INV_X1 U715 ( .A(G299), .ZN(n942) );
  NOR2_X1 U716 ( .A1(n668), .A2(n942), .ZN(n637) );
  XOR2_X1 U717 ( .A(KEYINPUT98), .B(KEYINPUT28), .Z(n636) );
  XNOR2_X1 U718 ( .A(n637), .B(n636), .ZN(n672) );
  NAND2_X1 U719 ( .A1(G81), .A2(n789), .ZN(n638) );
  XNOR2_X1 U720 ( .A(n638), .B(KEYINPUT12), .ZN(n639) );
  XNOR2_X1 U721 ( .A(n639), .B(KEYINPUT70), .ZN(n641) );
  NAND2_X1 U722 ( .A1(G68), .A2(n788), .ZN(n640) );
  NAND2_X1 U723 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U724 ( .A(KEYINPUT13), .B(n642), .ZN(n648) );
  NAND2_X1 U725 ( .A1(n785), .A2(G56), .ZN(n643) );
  XOR2_X1 U726 ( .A(KEYINPUT14), .B(n643), .Z(n646) );
  NAND2_X1 U727 ( .A1(G43), .A2(n784), .ZN(n644) );
  XNOR2_X1 U728 ( .A(KEYINPUT71), .B(n644), .ZN(n645) );
  NOR2_X1 U729 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U730 ( .A1(n648), .A2(n647), .ZN(n932) );
  NAND2_X1 U731 ( .A1(n660), .A2(G1996), .ZN(n649) );
  XNOR2_X1 U732 ( .A(n649), .B(KEYINPUT26), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n677), .A2(G1341), .ZN(n650) );
  NAND2_X1 U734 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U735 ( .A1(n932), .A2(n652), .ZN(n664) );
  NAND2_X1 U736 ( .A1(n784), .A2(G54), .ZN(n654) );
  NAND2_X1 U737 ( .A1(G66), .A2(n785), .ZN(n653) );
  NAND2_X1 U738 ( .A1(n654), .A2(n653), .ZN(n658) );
  NAND2_X1 U739 ( .A1(G79), .A2(n788), .ZN(n656) );
  NAND2_X1 U740 ( .A1(G92), .A2(n789), .ZN(n655) );
  NAND2_X1 U741 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U742 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U743 ( .A(n659), .B(KEYINPUT15), .ZN(n933) );
  NAND2_X1 U744 ( .A1(G1348), .A2(n677), .ZN(n662) );
  NAND2_X1 U745 ( .A1(G2067), .A2(n660), .ZN(n661) );
  NAND2_X1 U746 ( .A1(n662), .A2(n661), .ZN(n665) );
  NOR2_X1 U747 ( .A1(n933), .A2(n665), .ZN(n663) );
  OR2_X1 U748 ( .A1(n664), .A2(n663), .ZN(n667) );
  NAND2_X1 U749 ( .A1(n933), .A2(n665), .ZN(n666) );
  NAND2_X1 U750 ( .A1(n667), .A2(n666), .ZN(n670) );
  NAND2_X1 U751 ( .A1(n668), .A2(n942), .ZN(n669) );
  NAND2_X1 U752 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U753 ( .A1(n672), .A2(n671), .ZN(n674) );
  NAND2_X1 U754 ( .A1(n676), .A2(n675), .ZN(n690) );
  INV_X1 U755 ( .A(G8), .ZN(n683) );
  NOR2_X1 U756 ( .A1(G1971), .A2(n717), .ZN(n679) );
  NOR2_X1 U757 ( .A1(G2090), .A2(n677), .ZN(n678) );
  NOR2_X1 U758 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U759 ( .A1(n680), .A2(G303), .ZN(n681) );
  XNOR2_X1 U760 ( .A(n681), .B(KEYINPUT100), .ZN(n682) );
  OR2_X1 U761 ( .A1(n683), .A2(n682), .ZN(n685) );
  NAND2_X1 U762 ( .A1(n691), .A2(n684), .ZN(n688) );
  INV_X1 U763 ( .A(n685), .ZN(n686) );
  OR2_X1 U764 ( .A1(n686), .A2(G286), .ZN(n687) );
  NAND2_X1 U765 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U766 ( .A(n689), .B(KEYINPUT32), .ZN(n698) );
  AND2_X1 U767 ( .A1(n691), .A2(n690), .ZN(n696) );
  AND2_X1 U768 ( .A1(G8), .A2(n692), .ZN(n694) );
  OR2_X1 U769 ( .A1(n694), .A2(n693), .ZN(n695) );
  OR2_X1 U770 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U771 ( .A1(n698), .A2(n697), .ZN(n713) );
  NOR2_X1 U772 ( .A1(G1976), .A2(G288), .ZN(n705) );
  NOR2_X1 U773 ( .A1(G1971), .A2(G303), .ZN(n699) );
  NOR2_X1 U774 ( .A1(n705), .A2(n699), .ZN(n943) );
  NAND2_X1 U775 ( .A1(n713), .A2(n943), .ZN(n702) );
  NAND2_X1 U776 ( .A1(G1976), .A2(G288), .ZN(n937) );
  INV_X1 U777 ( .A(n937), .ZN(n700) );
  NOR2_X1 U778 ( .A1(n717), .A2(n700), .ZN(n701) );
  NAND2_X1 U779 ( .A1(n702), .A2(n701), .ZN(n704) );
  INV_X1 U780 ( .A(KEYINPUT33), .ZN(n703) );
  NAND2_X1 U781 ( .A1(n704), .A2(n703), .ZN(n710) );
  NAND2_X1 U782 ( .A1(n705), .A2(KEYINPUT33), .ZN(n706) );
  NOR2_X1 U783 ( .A1(n706), .A2(n717), .ZN(n708) );
  XOR2_X1 U784 ( .A(G1981), .B(G305), .Z(n929) );
  INV_X1 U785 ( .A(n929), .ZN(n707) );
  NOR2_X1 U786 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U787 ( .A1(n710), .A2(n709), .ZN(n722) );
  NOR2_X1 U788 ( .A1(G2090), .A2(G303), .ZN(n711) );
  NAND2_X1 U789 ( .A1(G8), .A2(n711), .ZN(n712) );
  NAND2_X1 U790 ( .A1(n713), .A2(n712), .ZN(n714) );
  AND2_X1 U791 ( .A1(n714), .A2(n717), .ZN(n720) );
  NOR2_X1 U792 ( .A1(G1981), .A2(G305), .ZN(n715) );
  XNOR2_X1 U793 ( .A(n715), .B(KEYINPUT24), .ZN(n716) );
  XNOR2_X1 U794 ( .A(n716), .B(KEYINPUT95), .ZN(n718) );
  NOR2_X1 U795 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U796 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U797 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U798 ( .A(n726), .B(n725), .ZN(n728) );
  XNOR2_X1 U799 ( .A(G1986), .B(G290), .ZN(n939) );
  NAND2_X1 U800 ( .A1(n939), .A2(n740), .ZN(n727) );
  NAND2_X1 U801 ( .A1(n728), .A2(n727), .ZN(n744) );
  NOR2_X1 U802 ( .A1(G1996), .A2(n857), .ZN(n993) );
  NOR2_X1 U803 ( .A1(G1986), .A2(G290), .ZN(n730) );
  AND2_X1 U804 ( .A1(n729), .A2(n870), .ZN(n999) );
  NOR2_X1 U805 ( .A1(n730), .A2(n999), .ZN(n731) );
  NOR2_X1 U806 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U807 ( .A1(n993), .A2(n733), .ZN(n734) );
  XNOR2_X1 U808 ( .A(n734), .B(KEYINPUT39), .ZN(n736) );
  NAND2_X1 U809 ( .A1(n736), .A2(n735), .ZN(n738) );
  NAND2_X1 U810 ( .A1(n737), .A2(n890), .ZN(n986) );
  NAND2_X1 U811 ( .A1(n738), .A2(n986), .ZN(n739) );
  XNOR2_X1 U812 ( .A(KEYINPUT102), .B(n739), .ZN(n741) );
  NAND2_X1 U813 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U814 ( .A(KEYINPUT103), .B(n742), .Z(n743) );
  NAND2_X1 U815 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U816 ( .A(n745), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U817 ( .A(G2438), .B(G2454), .Z(n747) );
  XNOR2_X1 U818 ( .A(G2435), .B(G2430), .ZN(n746) );
  XNOR2_X1 U819 ( .A(n747), .B(n746), .ZN(n748) );
  XOR2_X1 U820 ( .A(n748), .B(G2427), .Z(n750) );
  XNOR2_X1 U821 ( .A(G1341), .B(G1348), .ZN(n749) );
  XNOR2_X1 U822 ( .A(n750), .B(n749), .ZN(n754) );
  XOR2_X1 U823 ( .A(G2443), .B(G2446), .Z(n752) );
  XNOR2_X1 U824 ( .A(KEYINPUT104), .B(G2451), .ZN(n751) );
  XNOR2_X1 U825 ( .A(n752), .B(n751), .ZN(n753) );
  XOR2_X1 U826 ( .A(n754), .B(n753), .Z(n755) );
  AND2_X1 U827 ( .A1(G14), .A2(n755), .ZN(G401) );
  AND2_X1 U828 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U829 ( .A1(G111), .A2(n876), .ZN(n762) );
  NAND2_X1 U830 ( .A1(G99), .A2(n879), .ZN(n757) );
  NAND2_X1 U831 ( .A1(G135), .A2(n880), .ZN(n756) );
  NAND2_X1 U832 ( .A1(n757), .A2(n756), .ZN(n760) );
  NAND2_X1 U833 ( .A1(n875), .A2(G123), .ZN(n758) );
  XOR2_X1 U834 ( .A(KEYINPUT18), .B(n758), .Z(n759) );
  NOR2_X1 U835 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U836 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U837 ( .A(n763), .B(KEYINPUT80), .ZN(n1001) );
  XNOR2_X1 U838 ( .A(n1001), .B(G2096), .ZN(n764) );
  OR2_X1 U839 ( .A1(G2100), .A2(n764), .ZN(G156) );
  INV_X1 U840 ( .A(G132), .ZN(G219) );
  INV_X1 U841 ( .A(G82), .ZN(G220) );
  INV_X1 U842 ( .A(G57), .ZN(G237) );
  NAND2_X1 U843 ( .A1(G7), .A2(G661), .ZN(n765) );
  XNOR2_X1 U844 ( .A(n765), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U845 ( .A(G223), .B(KEYINPUT69), .ZN(n824) );
  NAND2_X1 U846 ( .A1(n824), .A2(G567), .ZN(n766) );
  XOR2_X1 U847 ( .A(KEYINPUT11), .B(n766), .Z(G234) );
  INV_X1 U848 ( .A(G860), .ZN(n783) );
  OR2_X1 U849 ( .A1(n932), .A2(n783), .ZN(G153) );
  XOR2_X1 U850 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  INV_X1 U851 ( .A(G868), .ZN(n770) );
  NOR2_X1 U852 ( .A1(G301), .A2(n770), .ZN(n768) );
  NOR2_X1 U853 ( .A1(G868), .A2(n933), .ZN(n767) );
  NOR2_X1 U854 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U855 ( .A(KEYINPUT73), .B(n769), .Z(G284) );
  NOR2_X1 U856 ( .A1(G286), .A2(n770), .ZN(n772) );
  NOR2_X1 U857 ( .A1(G868), .A2(G299), .ZN(n771) );
  NOR2_X1 U858 ( .A1(n772), .A2(n771), .ZN(G297) );
  NAND2_X1 U859 ( .A1(n783), .A2(G559), .ZN(n773) );
  INV_X1 U860 ( .A(n933), .ZN(n781) );
  NAND2_X1 U861 ( .A1(n773), .A2(n781), .ZN(n774) );
  XNOR2_X1 U862 ( .A(n774), .B(KEYINPUT16), .ZN(n775) );
  XOR2_X1 U863 ( .A(KEYINPUT77), .B(n775), .Z(G148) );
  NAND2_X1 U864 ( .A1(n781), .A2(G868), .ZN(n776) );
  NOR2_X1 U865 ( .A1(G559), .A2(n776), .ZN(n777) );
  XNOR2_X1 U866 ( .A(n777), .B(KEYINPUT78), .ZN(n779) );
  NOR2_X1 U867 ( .A1(n932), .A2(G868), .ZN(n778) );
  NOR2_X1 U868 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U869 ( .A(KEYINPUT79), .B(n780), .Z(G282) );
  NAND2_X1 U870 ( .A1(G559), .A2(n781), .ZN(n782) );
  XOR2_X1 U871 ( .A(n932), .B(n782), .Z(n804) );
  NAND2_X1 U872 ( .A1(n783), .A2(n804), .ZN(n794) );
  NAND2_X1 U873 ( .A1(n784), .A2(G55), .ZN(n787) );
  NAND2_X1 U874 ( .A1(G67), .A2(n785), .ZN(n786) );
  NAND2_X1 U875 ( .A1(n787), .A2(n786), .ZN(n793) );
  NAND2_X1 U876 ( .A1(G80), .A2(n788), .ZN(n791) );
  NAND2_X1 U877 ( .A1(G93), .A2(n789), .ZN(n790) );
  NAND2_X1 U878 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U879 ( .A1(n793), .A2(n792), .ZN(n806) );
  XOR2_X1 U880 ( .A(n794), .B(n806), .Z(G145) );
  INV_X1 U881 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U882 ( .A(KEYINPUT86), .B(KEYINPUT19), .ZN(n796) );
  XNOR2_X1 U883 ( .A(G288), .B(KEYINPUT87), .ZN(n795) );
  XNOR2_X1 U884 ( .A(n796), .B(n795), .ZN(n797) );
  XOR2_X1 U885 ( .A(n797), .B(KEYINPUT85), .Z(n799) );
  XNOR2_X1 U886 ( .A(G166), .B(KEYINPUT84), .ZN(n798) );
  XNOR2_X1 U887 ( .A(n799), .B(n798), .ZN(n800) );
  XNOR2_X1 U888 ( .A(n806), .B(n800), .ZN(n802) );
  XNOR2_X1 U889 ( .A(G290), .B(n942), .ZN(n801) );
  XNOR2_X1 U890 ( .A(n802), .B(n801), .ZN(n803) );
  XNOR2_X1 U891 ( .A(n803), .B(G305), .ZN(n893) );
  XNOR2_X1 U892 ( .A(n804), .B(n893), .ZN(n805) );
  NAND2_X1 U893 ( .A1(n805), .A2(G868), .ZN(n808) );
  OR2_X1 U894 ( .A1(G868), .A2(n806), .ZN(n807) );
  NAND2_X1 U895 ( .A1(n808), .A2(n807), .ZN(G295) );
  NAND2_X1 U896 ( .A1(G2078), .A2(G2084), .ZN(n809) );
  XOR2_X1 U897 ( .A(KEYINPUT20), .B(n809), .Z(n810) );
  NAND2_X1 U898 ( .A1(G2090), .A2(n810), .ZN(n811) );
  XNOR2_X1 U899 ( .A(KEYINPUT21), .B(n811), .ZN(n812) );
  NAND2_X1 U900 ( .A1(n812), .A2(G2072), .ZN(n813) );
  XNOR2_X1 U901 ( .A(KEYINPUT88), .B(n813), .ZN(G158) );
  XNOR2_X1 U902 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U903 ( .A1(G69), .A2(G120), .ZN(n814) );
  NOR2_X1 U904 ( .A1(G237), .A2(n814), .ZN(n815) );
  NAND2_X1 U905 ( .A1(G108), .A2(n815), .ZN(n904) );
  NAND2_X1 U906 ( .A1(G567), .A2(n904), .ZN(n816) );
  XNOR2_X1 U907 ( .A(n816), .B(KEYINPUT90), .ZN(n822) );
  NOR2_X1 U908 ( .A1(G220), .A2(G219), .ZN(n817) );
  XOR2_X1 U909 ( .A(KEYINPUT22), .B(n817), .Z(n818) );
  NOR2_X1 U910 ( .A1(G218), .A2(n818), .ZN(n819) );
  XOR2_X1 U911 ( .A(KEYINPUT89), .B(n819), .Z(n820) );
  NAND2_X1 U912 ( .A1(G96), .A2(n820), .ZN(n905) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n905), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n822), .A2(n821), .ZN(n830) );
  NAND2_X1 U915 ( .A1(G483), .A2(G661), .ZN(n823) );
  NOR2_X1 U916 ( .A1(n830), .A2(n823), .ZN(n827) );
  NAND2_X1 U917 ( .A1(n827), .A2(G36), .ZN(G176) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n824), .ZN(G217) );
  AND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n825) );
  NAND2_X1 U920 ( .A1(G661), .A2(n825), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n826) );
  XOR2_X1 U922 ( .A(KEYINPUT105), .B(n826), .Z(n828) );
  NAND2_X1 U923 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U924 ( .A(n829), .B(KEYINPUT106), .ZN(G188) );
  XNOR2_X1 U925 ( .A(KEYINPUT107), .B(n830), .ZN(G319) );
  XNOR2_X1 U926 ( .A(G1981), .B(KEYINPUT41), .ZN(n840) );
  XOR2_X1 U927 ( .A(G1976), .B(G1971), .Z(n832) );
  XNOR2_X1 U928 ( .A(G1966), .B(G1961), .ZN(n831) );
  XNOR2_X1 U929 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U930 ( .A(G1956), .B(G1996), .Z(n834) );
  XNOR2_X1 U931 ( .A(G1986), .B(G1991), .ZN(n833) );
  XNOR2_X1 U932 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U933 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U934 ( .A(KEYINPUT108), .B(G2474), .ZN(n837) );
  XNOR2_X1 U935 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n840), .B(n839), .ZN(G229) );
  XOR2_X1 U937 ( .A(G2100), .B(G2096), .Z(n842) );
  XNOR2_X1 U938 ( .A(KEYINPUT42), .B(G2678), .ZN(n841) );
  XNOR2_X1 U939 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U940 ( .A(KEYINPUT43), .B(G2090), .Z(n844) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2072), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U943 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U944 ( .A(G2078), .B(G2084), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(G227) );
  NAND2_X1 U946 ( .A1(G124), .A2(n875), .ZN(n849) );
  XOR2_X1 U947 ( .A(KEYINPUT44), .B(n849), .Z(n850) );
  XNOR2_X1 U948 ( .A(n850), .B(KEYINPUT109), .ZN(n852) );
  NAND2_X1 U949 ( .A1(G100), .A2(n879), .ZN(n851) );
  NAND2_X1 U950 ( .A1(n852), .A2(n851), .ZN(n856) );
  NAND2_X1 U951 ( .A1(G136), .A2(n880), .ZN(n854) );
  NAND2_X1 U952 ( .A1(G112), .A2(n876), .ZN(n853) );
  NAND2_X1 U953 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U954 ( .A1(n856), .A2(n855), .ZN(G162) );
  XNOR2_X1 U955 ( .A(G162), .B(n857), .ZN(n859) );
  XNOR2_X1 U956 ( .A(G164), .B(G160), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n859), .B(n858), .ZN(n874) );
  XOR2_X1 U958 ( .A(KEYINPUT48), .B(KEYINPUT113), .Z(n868) );
  NAND2_X1 U959 ( .A1(G103), .A2(n879), .ZN(n861) );
  NAND2_X1 U960 ( .A1(G139), .A2(n880), .ZN(n860) );
  NAND2_X1 U961 ( .A1(n861), .A2(n860), .ZN(n866) );
  NAND2_X1 U962 ( .A1(G127), .A2(n875), .ZN(n863) );
  NAND2_X1 U963 ( .A1(G115), .A2(n876), .ZN(n862) );
  NAND2_X1 U964 ( .A1(n863), .A2(n862), .ZN(n864) );
  XOR2_X1 U965 ( .A(KEYINPUT47), .B(n864), .Z(n865) );
  NOR2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n988) );
  XNOR2_X1 U967 ( .A(n988), .B(KEYINPUT111), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U969 ( .A(n869), .B(KEYINPUT112), .Z(n872) );
  XNOR2_X1 U970 ( .A(n870), .B(KEYINPUT46), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U972 ( .A(n874), .B(n873), .Z(n889) );
  NAND2_X1 U973 ( .A1(G130), .A2(n875), .ZN(n878) );
  NAND2_X1 U974 ( .A1(G118), .A2(n876), .ZN(n877) );
  NAND2_X1 U975 ( .A1(n878), .A2(n877), .ZN(n886) );
  NAND2_X1 U976 ( .A1(G106), .A2(n879), .ZN(n882) );
  NAND2_X1 U977 ( .A1(G142), .A2(n880), .ZN(n881) );
  NAND2_X1 U978 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U979 ( .A(KEYINPUT45), .B(n883), .Z(n884) );
  XNOR2_X1 U980 ( .A(KEYINPUT110), .B(n884), .ZN(n885) );
  NOR2_X1 U981 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U982 ( .A(n1001), .B(n887), .ZN(n888) );
  XNOR2_X1 U983 ( .A(n889), .B(n888), .ZN(n891) );
  XOR2_X1 U984 ( .A(n891), .B(n890), .Z(n892) );
  NOR2_X1 U985 ( .A1(G37), .A2(n892), .ZN(G395) );
  XNOR2_X1 U986 ( .A(n893), .B(KEYINPUT114), .ZN(n895) );
  XNOR2_X1 U987 ( .A(n933), .B(G286), .ZN(n894) );
  XNOR2_X1 U988 ( .A(n895), .B(n894), .ZN(n897) );
  XOR2_X1 U989 ( .A(n932), .B(G171), .Z(n896) );
  XNOR2_X1 U990 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U991 ( .A1(G37), .A2(n898), .ZN(G397) );
  NOR2_X1 U992 ( .A1(G229), .A2(G227), .ZN(n899) );
  XNOR2_X1 U993 ( .A(KEYINPUT49), .B(n899), .ZN(n900) );
  NOR2_X1 U994 ( .A1(G401), .A2(n900), .ZN(n902) );
  NOR2_X1 U995 ( .A1(G395), .A2(G397), .ZN(n901) );
  AND2_X1 U996 ( .A1(n902), .A2(n901), .ZN(n903) );
  NAND2_X1 U997 ( .A1(G319), .A2(n903), .ZN(G225) );
  XNOR2_X1 U998 ( .A(KEYINPUT115), .B(G225), .ZN(G308) );
  INV_X1 U1000 ( .A(G120), .ZN(G236) );
  INV_X1 U1001 ( .A(G96), .ZN(G221) );
  INV_X1 U1002 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1003 ( .A1(n905), .A2(n904), .ZN(G325) );
  INV_X1 U1004 ( .A(G325), .ZN(G261) );
  INV_X1 U1005 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1006 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n1016) );
  INV_X1 U1007 ( .A(KEYINPUT55), .ZN(n1010) );
  XNOR2_X1 U1008 ( .A(G2084), .B(G34), .ZN(n906) );
  XNOR2_X1 U1009 ( .A(n906), .B(KEYINPUT54), .ZN(n908) );
  XNOR2_X1 U1010 ( .A(G35), .B(G2090), .ZN(n907) );
  NOR2_X1 U1011 ( .A1(n908), .A2(n907), .ZN(n924) );
  XNOR2_X1 U1012 ( .A(G1991), .B(G25), .ZN(n910) );
  XNOR2_X1 U1013 ( .A(G33), .B(G2072), .ZN(n909) );
  NOR2_X1 U1014 ( .A1(n910), .A2(n909), .ZN(n917) );
  XOR2_X1 U1015 ( .A(G2067), .B(G26), .Z(n911) );
  NAND2_X1 U1016 ( .A1(n911), .A2(G28), .ZN(n915) );
  XOR2_X1 U1017 ( .A(G27), .B(n912), .Z(n913) );
  XNOR2_X1 U1018 ( .A(KEYINPUT118), .B(n913), .ZN(n914) );
  NOR2_X1 U1019 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1020 ( .A1(n917), .A2(n916), .ZN(n920) );
  XOR2_X1 U1021 ( .A(G32), .B(G1996), .Z(n918) );
  XNOR2_X1 U1022 ( .A(KEYINPUT119), .B(n918), .ZN(n919) );
  NOR2_X1 U1023 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1024 ( .A(n921), .B(KEYINPUT53), .Z(n922) );
  XNOR2_X1 U1025 ( .A(KEYINPUT120), .B(n922), .ZN(n923) );
  NAND2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1027 ( .A(n1010), .B(n925), .ZN(n927) );
  INV_X1 U1028 ( .A(G29), .ZN(n926) );
  NAND2_X1 U1029 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1030 ( .A1(G11), .A2(n928), .ZN(n985) );
  XNOR2_X1 U1031 ( .A(G16), .B(KEYINPUT56), .ZN(n953) );
  XNOR2_X1 U1032 ( .A(G1966), .B(G168), .ZN(n930) );
  NAND2_X1 U1033 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1034 ( .A(n931), .B(KEYINPUT57), .ZN(n951) );
  XNOR2_X1 U1035 ( .A(n932), .B(G1341), .ZN(n949) );
  XOR2_X1 U1036 ( .A(G171), .B(G1961), .Z(n935) );
  XNOR2_X1 U1037 ( .A(n933), .B(G1348), .ZN(n934) );
  NOR2_X1 U1038 ( .A1(n935), .A2(n934), .ZN(n941) );
  NAND2_X1 U1039 ( .A1(G1971), .A2(G303), .ZN(n936) );
  NAND2_X1 U1040 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1041 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1042 ( .A1(n941), .A2(n940), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(n942), .B(G1956), .ZN(n944) );
  NAND2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1046 ( .A(KEYINPUT121), .B(n947), .ZN(n948) );
  NOR2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n983) );
  INV_X1 U1050 ( .A(G16), .ZN(n981) );
  XNOR2_X1 U1051 ( .A(G5), .B(n954), .ZN(n955) );
  XNOR2_X1 U1052 ( .A(n955), .B(KEYINPUT122), .ZN(n976) );
  XNOR2_X1 U1053 ( .A(n956), .B(G20), .ZN(n965) );
  XOR2_X1 U1054 ( .A(KEYINPUT124), .B(G4), .Z(n958) );
  XNOR2_X1 U1055 ( .A(G1348), .B(KEYINPUT59), .ZN(n957) );
  XNOR2_X1 U1056 ( .A(n958), .B(n957), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(G1341), .B(G19), .ZN(n960) );
  XNOR2_X1 U1058 ( .A(G1981), .B(G6), .ZN(n959) );
  NOR2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1060 ( .A(n961), .B(KEYINPUT123), .ZN(n962) );
  NOR2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1063 ( .A(n966), .B(KEYINPUT60), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n972) );
  XOR2_X1 U1065 ( .A(G1986), .B(G24), .Z(n970) );
  XNOR2_X1 U1066 ( .A(G1971), .B(G22), .ZN(n968) );
  XNOR2_X1 U1067 ( .A(G23), .B(G1976), .ZN(n967) );
  NOR2_X1 U1068 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1069 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1070 ( .A(n972), .B(n971), .Z(n973) );
  NOR2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(G21), .B(G1966), .ZN(n977) );
  NOR2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1075 ( .A(KEYINPUT61), .B(n979), .ZN(n980) );
  NAND2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n1014) );
  NAND2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n1008) );
  XOR2_X1 U1080 ( .A(G2072), .B(n988), .Z(n990) );
  XOR2_X1 U1081 ( .A(G164), .B(G2078), .Z(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1083 ( .A(KEYINPUT50), .B(n991), .Z(n997) );
  XOR2_X1 U1084 ( .A(G2090), .B(G162), .Z(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1086 ( .A(KEYINPUT117), .B(n994), .Z(n995) );
  XNOR2_X1 U1087 ( .A(KEYINPUT51), .B(n995), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n1006) );
  XOR2_X1 U1089 ( .A(G2084), .B(G160), .Z(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(n1004), .B(KEYINPUT116), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(KEYINPUT52), .B(n1009), .ZN(n1011) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(G29), .ZN(n1013) );
  NAND2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1100 ( .A(n1016), .B(n1015), .ZN(G311) );
  XNOR2_X1 U1101 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

