//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n820,
    new_n822, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1026, new_n1027, new_n1028, new_n1029, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1037, new_n1038,
    new_n1039;
  INV_X1    g000(.A(G227gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT27), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT65), .B1(new_n205), .B2(G183gat), .ZN(new_n206));
  AOI21_X1  g005(.A(G190gat), .B1(new_n205), .B2(G183gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n208));
  INV_X1    g007(.A(G183gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT27), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n206), .A2(new_n207), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT28), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n209), .A2(KEYINPUT27), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n207), .A2(KEYINPUT28), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT66), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n207), .A2(new_n217), .A3(KEYINPUT28), .A4(new_n214), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n213), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT26), .ZN(new_n222));
  INV_X1    g021(.A(G169gat), .ZN(new_n223));
  INV_X1    g022(.A(G176gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT67), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(KEYINPUT67), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n223), .A2(new_n224), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n231), .B1(KEYINPUT26), .B2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n221), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT23), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT23), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n237), .B1(G169gat), .B2(G176gat), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n236), .A2(new_n238), .A3(new_n230), .ZN(new_n239));
  NOR2_X1   g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT64), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n220), .A2(KEYINPUT24), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT24), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(G183gat), .A3(G190gat), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g045(.A(KEYINPUT25), .B(new_n239), .C1(new_n242), .C2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n240), .B1(new_n243), .B2(new_n245), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n236), .A2(new_n238), .A3(new_n230), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G127gat), .B(G134gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n254));
  INV_X1    g053(.A(G113gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n255), .A2(G120gat), .ZN(new_n256));
  INV_X1    g055(.A(G120gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n257), .A2(G113gat), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n253), .B(new_n254), .C1(new_n256), .C2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G113gat), .B(G120gat), .ZN(new_n260));
  INV_X1    g059(.A(G127gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(G134gat), .ZN(new_n262));
  INV_X1    g061(.A(G134gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(G127gat), .ZN(new_n264));
  OAI22_X1  g063(.A1(new_n260), .A2(KEYINPUT1), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n235), .A2(new_n252), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n266), .B1(new_n235), .B2(new_n252), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n204), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT33), .ZN(new_n270));
  XNOR2_X1  g069(.A(G15gat), .B(G43gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT70), .ZN(new_n272));
  XNOR2_X1  g071(.A(G71gat), .B(G99gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n269), .B(KEYINPUT32), .C1(new_n270), .C2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n204), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n235), .A2(new_n252), .ZN(new_n277));
  INV_X1    g076(.A(new_n266), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n235), .A2(new_n252), .A3(new_n266), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT68), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n281), .A2(new_n282), .A3(KEYINPUT33), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT68), .B1(new_n269), .B2(new_n270), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT69), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT32), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n286), .B1(new_n281), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n274), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n269), .A2(KEYINPUT69), .A3(KEYINPUT32), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n275), .B1(new_n285), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n267), .A2(new_n268), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(new_n276), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT34), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT34), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n293), .A2(new_n296), .A3(new_n276), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n292), .A2(new_n299), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n298), .B(new_n275), .C1(new_n285), .C2(new_n291), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(KEYINPUT71), .A3(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n282), .B1(new_n281), .B2(KEYINPUT33), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n269), .A2(KEYINPUT68), .A3(new_n270), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n269), .A2(KEYINPUT32), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n274), .B1(new_n306), .B2(new_n286), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n305), .A2(new_n307), .A3(new_n290), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n298), .B1(new_n308), .B2(new_n275), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT71), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G78gat), .B(G106gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT31), .B(G50gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G22gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(G228gat), .A2(G233gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n318));
  AND2_X1   g117(.A1(G211gat), .A2(G218gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(G211gat), .A2(G218gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n318), .B1(new_n321), .B2(KEYINPUT73), .ZN(new_n322));
  INV_X1    g121(.A(G197gat), .ZN(new_n323));
  INV_X1    g122(.A(G204gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G197gat), .A2(G204gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT22), .ZN(new_n327));
  NAND2_X1  g126(.A1(G211gat), .A2(G218gat), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n325), .A2(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n322), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT73), .B1(new_n329), .B2(new_n318), .ZN(new_n332));
  INV_X1    g131(.A(new_n321), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT3), .ZN(new_n336));
  INV_X1    g135(.A(G148gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G141gat), .ZN(new_n338));
  INV_X1    g137(.A(G141gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(G148gat), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT2), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G155gat), .B(G162gat), .ZN(new_n342));
  OAI21_X1  g141(.A(KEYINPUT76), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G155gat), .A2(G162gat), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT76), .ZN(new_n348));
  XNOR2_X1  g147(.A(G141gat), .B(G148gat), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n347), .B(new_n348), .C1(new_n349), .C2(KEYINPUT2), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n343), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT2), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n346), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n339), .ZN(new_n356));
  NAND2_X1  g155(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(G148gat), .A3(new_n357), .ZN(new_n358));
  AOI221_X4 g157(.A(new_n352), .B1(new_n354), .B2(new_n344), .C1(new_n358), .C2(new_n338), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n338), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n354), .A2(new_n344), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT78), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n336), .B(new_n351), .C1(new_n359), .C2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n335), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n338), .ZN(new_n366));
  AND2_X1   g165(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n366), .B1(new_n369), .B2(G148gat), .ZN(new_n370));
  INV_X1    g169(.A(new_n361), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n352), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n360), .A2(KEYINPUT78), .A3(new_n361), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n372), .A2(new_n373), .B1(new_n343), .B2(new_n350), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT29), .B1(new_n330), .B2(new_n333), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n329), .A2(new_n321), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT3), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n317), .B1(new_n365), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT79), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n381), .A3(new_n334), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n336), .B1(new_n334), .B2(KEYINPUT29), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n351), .B1(new_n359), .B2(new_n362), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n317), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n365), .A2(new_n381), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n316), .B(new_n379), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT80), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n315), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n379), .B1(new_n386), .B2(new_n387), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(G22gat), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n394));
  AND3_X1   g193(.A1(new_n393), .A2(new_n394), .A3(new_n388), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n394), .B1(new_n393), .B2(new_n388), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n391), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n388), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n334), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT79), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(new_n382), .A3(new_n385), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n316), .B1(new_n401), .B2(new_n379), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT81), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n393), .A2(new_n394), .A3(new_n388), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(new_n390), .A3(new_n404), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n302), .A2(new_n311), .B1(new_n397), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n384), .A2(KEYINPUT3), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(new_n363), .A3(new_n278), .ZN(new_n408));
  NAND2_X1  g207(.A1(G225gat), .A2(G233gat), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n266), .B(new_n351), .C1(new_n359), .C2(new_n362), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT4), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n374), .A2(KEYINPUT4), .A3(new_n266), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n408), .A2(new_n409), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT5), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n384), .A2(new_n278), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n410), .ZN(new_n417));
  INV_X1    g216(.A(new_n409), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n415), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n413), .A2(new_n412), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n421), .A2(new_n415), .A3(new_n409), .A4(new_n408), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G1gat), .B(G29gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(KEYINPUT0), .ZN(new_n425));
  XNOR2_X1  g224(.A(G57gat), .B(G85gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n420), .A2(new_n427), .A3(new_n422), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n427), .B1(new_n420), .B2(new_n422), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT6), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(G226gat), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n436), .A2(new_n203), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n437), .A2(KEYINPUT29), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n277), .A2(KEYINPUT74), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT74), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n235), .A2(new_n252), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n439), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n277), .A2(new_n436), .A3(new_n203), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n335), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n440), .A2(new_n437), .A3(new_n442), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n277), .A2(new_n438), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(new_n334), .A3(new_n447), .ZN(new_n448));
  XOR2_X1   g247(.A(G8gat), .B(G36gat), .Z(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(KEYINPUT75), .ZN(new_n450));
  XNOR2_X1  g249(.A(G64gat), .B(G92gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n445), .A2(new_n448), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT30), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n445), .A2(KEYINPUT30), .A3(new_n448), .A4(new_n452), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n445), .A2(new_n448), .ZN(new_n457));
  INV_X1    g256(.A(new_n452), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n455), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n435), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n406), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT35), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n429), .A2(KEYINPUT83), .A3(new_n430), .A4(new_n431), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n434), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n433), .A2(KEYINPUT6), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT83), .B1(new_n468), .B2(new_n431), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n461), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT84), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT35), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n300), .A2(new_n472), .A3(new_n301), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n473), .B1(new_n405), .B2(new_n397), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT83), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n432), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n476), .A2(new_n434), .A3(new_n466), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT84), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n478), .A3(new_n461), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n471), .A2(new_n474), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n409), .B1(new_n421), .B2(new_n408), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT39), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n428), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n408), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n413), .A2(new_n412), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n418), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT82), .B1(new_n417), .B2(new_n418), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT82), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n416), .A2(new_n488), .A3(new_n409), .A4(new_n410), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n486), .A2(new_n490), .A3(KEYINPUT39), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n483), .A2(new_n491), .A3(KEYINPUT40), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT40), .B1(new_n483), .B2(new_n491), .ZN(new_n493));
  NOR3_X1   g292(.A1(new_n492), .A2(new_n493), .A3(new_n433), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n494), .A2(new_n460), .B1(new_n397), .B2(new_n405), .ZN(new_n495));
  INV_X1    g294(.A(new_n434), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n420), .A2(new_n427), .A3(new_n422), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n497), .A2(new_n433), .A3(KEYINPUT6), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n496), .B1(new_n498), .B2(KEYINPUT83), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT37), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n445), .A2(new_n500), .A3(new_n448), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n458), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n500), .B1(new_n445), .B2(new_n448), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT38), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n457), .A2(new_n458), .ZN(new_n505));
  INV_X1    g304(.A(new_n502), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n446), .A2(new_n335), .A3(new_n447), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n507), .A2(KEYINPUT37), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n334), .B1(new_n443), .B2(new_n444), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT38), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n505), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n499), .A2(new_n476), .A3(new_n504), .A4(new_n511), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n403), .A2(new_n390), .A3(new_n404), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n390), .B1(new_n403), .B2(new_n404), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n495), .A2(new_n512), .B1(new_n462), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n300), .A2(new_n301), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT36), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI211_X1 g318(.A(KEYINPUT71), .B(new_n298), .C1(new_n308), .C2(new_n275), .ZN(new_n520));
  INV_X1    g319(.A(new_n301), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(new_n309), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n520), .B1(new_n522), .B2(KEYINPUT71), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n519), .B1(new_n523), .B2(new_n518), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n465), .A2(new_n480), .B1(new_n516), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT86), .ZN(new_n527));
  INV_X1    g326(.A(G1gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n526), .A2(KEYINPUT86), .A3(G1gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT16), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT87), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n526), .A2(new_n531), .B1(new_n532), .B2(G8gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n529), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n532), .A2(G8gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G29gat), .A2(G36gat), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NOR3_X1   g339(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G43gat), .B(G50gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(KEYINPUT15), .A3(new_n543), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n543), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(KEYINPUT15), .B2(new_n543), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT85), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n541), .A2(new_n547), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n540), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n544), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n537), .A2(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n551), .A2(KEYINPUT17), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n554), .B(new_n544), .C1(new_n546), .C2(new_n550), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n536), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G229gat), .A2(G233gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n552), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT18), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT88), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n558), .B(KEYINPUT13), .Z(new_n564));
  INV_X1    g363(.A(new_n552), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n537), .A2(new_n551), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n552), .A2(new_n557), .A3(new_n558), .A4(new_n561), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n563), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G113gat), .B(G141gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G197gat), .ZN(new_n571));
  XOR2_X1   g370(.A(KEYINPUT11), .B(G169gat), .Z(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT12), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n563), .A2(new_n567), .A3(new_n574), .A4(new_n568), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n525), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G190gat), .B(G218gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT96), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT93), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(KEYINPUT93), .A2(G99gat), .A3(G106gat), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n587), .A2(KEYINPUT8), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(G85gat), .ZN(new_n590));
  INV_X1    g389(.A(G92gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT94), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT94), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n589), .A2(new_n595), .A3(new_n592), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT95), .ZN(new_n598));
  XOR2_X1   g397(.A(G99gat), .B(G106gat), .Z(new_n599));
  INV_X1    g398(.A(KEYINPUT7), .ZN(new_n600));
  OAI211_X1 g399(.A(G85gat), .B(G92gat), .C1(new_n600), .C2(KEYINPUT92), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(KEYINPUT92), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n597), .A2(new_n598), .A3(new_n599), .A4(new_n603), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n589), .A2(new_n595), .A3(new_n592), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n595), .B1(new_n589), .B2(new_n592), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n599), .A2(new_n598), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n599), .A2(new_n598), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n604), .B(new_n610), .C1(new_n553), .C2(new_n556), .ZN(new_n611));
  AND2_X1   g410(.A1(G232gat), .A2(G233gat), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n581), .A2(new_n582), .B1(KEYINPUT41), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n610), .A2(new_n604), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n614), .B1(new_n615), .B2(new_n551), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n584), .B1(new_n611), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n612), .A2(KEYINPUT41), .ZN(new_n619));
  XNOR2_X1  g418(.A(G134gat), .B(G162gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n611), .A2(new_n616), .A3(new_n584), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n618), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n621), .ZN(new_n624));
  INV_X1    g423(.A(new_n622), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n624), .B1(new_n625), .B2(new_n617), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n629));
  INV_X1    g428(.A(G57gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(G64gat), .ZN(new_n631));
  INV_X1    g430(.A(G64gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(G57gat), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n629), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT89), .ZN(new_n635));
  NAND2_X1  g434(.A1(G71gat), .A2(G78gat), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(G71gat), .A2(G78gat), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OR2_X1    g438(.A1(G71gat), .A2(G78gat), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n640), .A2(KEYINPUT89), .A3(new_n636), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n634), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n636), .ZN(new_n643));
  XNOR2_X1  g442(.A(G57gat), .B(G64gat), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n643), .B(new_n635), .C1(new_n644), .C2(new_n629), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT90), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n642), .A2(new_n645), .A3(KEYINPUT90), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT21), .ZN(new_n651));
  NAND2_X1  g450(.A1(G231gat), .A2(G233gat), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n652), .B1(new_n650), .B2(new_n651), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n261), .ZN(new_n657));
  OAI21_X1  g456(.A(G127gat), .B1(new_n654), .B2(new_n655), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT91), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n642), .A2(KEYINPUT90), .A3(new_n645), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT90), .B1(new_n642), .B2(new_n645), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n648), .A2(KEYINPUT91), .A3(new_n649), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n659), .B(new_n536), .C1(new_n651), .C2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n536), .B1(new_n666), .B2(new_n651), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n657), .A2(new_n668), .A3(new_n658), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n671));
  INV_X1    g470(.A(G155gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(G183gat), .B(G211gat), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n673), .B(new_n674), .Z(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n670), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n667), .A2(new_n669), .A3(new_n675), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n628), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n665), .A2(new_n615), .A3(KEYINPUT10), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT98), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n599), .A2(KEYINPUT97), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n607), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n607), .A2(new_n684), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(new_n646), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT10), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n610), .A2(new_n604), .A3(new_n650), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n665), .A2(new_n615), .A3(KEYINPUT98), .A4(KEYINPUT10), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n683), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(G230gat), .A2(G233gat), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n687), .A2(new_n689), .ZN(new_n695));
  INV_X1    g494(.A(new_n693), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(G120gat), .B(G148gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(G176gat), .B(G204gat), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n699), .B(new_n700), .Z(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n694), .A2(new_n697), .A3(new_n701), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n680), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n580), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n435), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(new_n528), .ZN(G1324gat));
  NAND3_X1  g508(.A1(new_n580), .A2(new_n460), .A3(new_n706), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT42), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT16), .B(G8gat), .ZN(new_n712));
  OR3_X1    g511(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT99), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n710), .A2(G8gat), .ZN(new_n717));
  OAI22_X1  g516(.A1(new_n717), .A2(new_n711), .B1(new_n710), .B2(new_n712), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n715), .B1(new_n716), .B2(new_n718), .ZN(G1325gat));
  INV_X1    g518(.A(KEYINPUT100), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n720), .B(new_n519), .C1(new_n523), .C2(new_n518), .ZN(new_n721));
  INV_X1    g520(.A(new_n519), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n518), .B1(new_n302), .B2(new_n311), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT100), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(G15gat), .B1(new_n707), .B2(new_n726), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n517), .A2(G15gat), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n707), .B2(new_n728), .ZN(G1326gat));
  NAND2_X1  g528(.A1(new_n397), .A2(new_n405), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n707), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g530(.A(KEYINPUT43), .B(G22gat), .Z(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(G1327gat));
  NAND2_X1  g532(.A1(new_n465), .A2(new_n480), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n483), .A2(new_n491), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT40), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n483), .A2(new_n491), .A3(KEYINPUT40), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n460), .A2(new_n737), .A3(new_n429), .A4(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n508), .A2(new_n509), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT38), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n740), .A2(new_n501), .A3(new_n741), .A4(new_n458), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n504), .A2(new_n742), .A3(new_n453), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n730), .B(new_n739), .C1(new_n477), .C2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n515), .A2(new_n462), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n744), .B(new_n745), .C1(new_n722), .C2(new_n723), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n627), .B1(new_n734), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n677), .A2(new_n678), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n705), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(new_n579), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n752), .A2(G29gat), .A3(new_n435), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n753), .B(KEYINPUT45), .Z(new_n754));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT101), .B1(new_n747), .B2(new_n755), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n471), .A2(new_n479), .A3(new_n474), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n472), .B1(new_n406), .B2(new_n463), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n467), .A3(new_n469), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n739), .B1(new_n513), .B2(new_n514), .ZN(new_n761));
  OAI22_X1  g560(.A1(new_n760), .A2(new_n761), .B1(new_n463), .B2(new_n730), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n762), .B1(new_n721), .B2(new_n724), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n755), .B(new_n628), .C1(new_n759), .C2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT101), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n765), .B(KEYINPUT44), .C1(new_n525), .C2(new_n627), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n756), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n751), .ZN(new_n768));
  OAI21_X1  g567(.A(G29gat), .B1(new_n768), .B2(new_n435), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n769), .ZN(G1328gat));
  OAI21_X1  g569(.A(G36gat), .B1(new_n768), .B2(new_n461), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n752), .A2(G36gat), .A3(new_n461), .ZN(new_n772));
  XNOR2_X1  g571(.A(KEYINPUT102), .B(KEYINPUT46), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n771), .A2(new_n774), .ZN(G1329gat));
  OAI21_X1  g574(.A(G43gat), .B1(new_n768), .B2(new_n726), .ZN(new_n776));
  OR3_X1    g575(.A1(new_n752), .A2(G43gat), .A3(new_n517), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT103), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT47), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n778), .B(new_n780), .ZN(G1330gat));
  INV_X1    g580(.A(KEYINPUT48), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n764), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n746), .B1(new_n757), .B2(new_n758), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n628), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n765), .B1(new_n785), .B2(KEYINPUT44), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n515), .B(new_n751), .C1(new_n783), .C2(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n787), .A2(G50gat), .ZN(new_n788));
  NOR4_X1   g587(.A1(new_n750), .A2(G50gat), .A3(new_n730), .A4(new_n627), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n580), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n790), .B(KEYINPUT104), .Z(new_n791));
  OAI21_X1  g590(.A(new_n782), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n580), .A2(KEYINPUT105), .A3(new_n789), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT105), .B1(new_n580), .B2(new_n789), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT48), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(G50gat), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n796), .B1(new_n787), .B2(KEYINPUT106), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT106), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n767), .A2(new_n798), .A3(new_n515), .A4(new_n751), .ZN(new_n799));
  AOI211_X1 g598(.A(KEYINPUT107), .B(new_n795), .C1(new_n797), .C2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT107), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n787), .A2(KEYINPUT106), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(G50gat), .A3(new_n799), .ZN(new_n803));
  INV_X1    g602(.A(new_n795), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n792), .B1(new_n800), .B2(new_n805), .ZN(G1331gat));
  NOR2_X1   g605(.A1(new_n759), .A2(new_n763), .ZN(new_n807));
  INV_X1    g606(.A(new_n705), .ZN(new_n808));
  NOR4_X1   g607(.A1(new_n807), .A2(new_n578), .A3(new_n680), .A4(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n435), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g611(.A(new_n461), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT108), .ZN(new_n815));
  NOR2_X1   g614(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n815), .B(new_n816), .ZN(G1333gat));
  NAND2_X1  g616(.A1(new_n809), .A2(new_n725), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n517), .A2(G71gat), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n818), .A2(G71gat), .B1(new_n809), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g620(.A1(new_n809), .A2(new_n515), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g622(.A1(new_n748), .A2(new_n578), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n628), .B(new_n824), .C1(new_n759), .C2(new_n763), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT109), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n825), .A2(new_n826), .ZN(new_n830));
  OR3_X1    g629(.A1(new_n825), .A2(new_n828), .A3(new_n826), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n705), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n810), .A2(new_n590), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n783), .A2(new_n786), .ZN(new_n835));
  INV_X1    g634(.A(new_n824), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(new_n808), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n835), .A2(new_n435), .A3(new_n838), .ZN(new_n839));
  OAI22_X1  g638(.A1(new_n833), .A2(new_n834), .B1(new_n590), .B2(new_n839), .ZN(G1336gat));
  NOR2_X1   g639(.A1(new_n835), .A2(new_n838), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n460), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(G92gat), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n460), .A2(new_n591), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n833), .A2(new_n846), .ZN(new_n847));
  AOI211_X1 g646(.A(new_n808), .B(new_n846), .C1(new_n827), .C2(new_n830), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n848), .B1(new_n842), .B2(G92gat), .ZN(new_n849));
  OAI22_X1  g648(.A1(new_n845), .A2(new_n847), .B1(new_n849), .B2(new_n844), .ZN(G1337gat));
  NOR3_X1   g649(.A1(new_n835), .A2(new_n726), .A3(new_n838), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n851), .A2(KEYINPUT110), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(KEYINPUT110), .ZN(new_n853));
  XOR2_X1   g652(.A(KEYINPUT111), .B(G99gat), .Z(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n808), .A2(new_n517), .A3(new_n854), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT112), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n832), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n855), .A2(new_n858), .ZN(G1338gat));
  NOR3_X1   g658(.A1(new_n730), .A2(new_n808), .A3(G106gat), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n832), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n515), .B(new_n837), .C1(new_n783), .C2(new_n786), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(G106gat), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n827), .A2(new_n830), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n860), .B(KEYINPUT113), .Z(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT114), .B1(new_n869), .B2(KEYINPUT53), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n871));
  AOI211_X1 g670(.A(new_n871), .B(new_n862), .C1(new_n864), .C2(new_n868), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n865), .B1(new_n870), .B2(new_n872), .ZN(G1339gat));
  INV_X1    g672(.A(new_n748), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n683), .A2(new_n696), .A3(new_n690), .A4(new_n691), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n694), .A2(KEYINPUT54), .A3(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n692), .A2(new_n877), .A3(new_n693), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n876), .A2(KEYINPUT55), .A3(new_n702), .A4(new_n878), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n879), .A2(new_n704), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT55), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n694), .A2(KEYINPUT54), .A3(new_n875), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n878), .A2(new_n702), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n565), .A2(new_n566), .A3(new_n564), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n558), .B1(new_n552), .B2(new_n557), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n573), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AND4_X1   g687(.A1(new_n577), .A2(new_n888), .A3(new_n623), .A4(new_n626), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n880), .A2(new_n881), .A3(new_n885), .A4(new_n889), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n885), .A2(new_n704), .A3(new_n879), .A4(new_n889), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT116), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n885), .A2(new_n578), .A3(new_n704), .A4(new_n879), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n888), .A2(new_n577), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n705), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n628), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n874), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n679), .A2(new_n579), .A3(new_n808), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT115), .ZN(new_n900));
  AOI211_X1 g699(.A(new_n517), .B(new_n515), .C1(new_n898), .C2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n810), .A3(new_n461), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n902), .A2(new_n255), .A3(new_n579), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n435), .B1(new_n898), .B2(new_n900), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n904), .A2(new_n406), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(new_n461), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n578), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n903), .B1(new_n907), .B2(new_n255), .ZN(G1340gat));
  NOR3_X1   g707(.A1(new_n902), .A2(new_n257), .A3(new_n808), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n906), .A2(new_n705), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n257), .ZN(G1341gat));
  NAND3_X1  g710(.A1(new_n906), .A2(new_n261), .A3(new_n748), .ZN(new_n912));
  OAI21_X1  g711(.A(G127gat), .B1(new_n902), .B2(new_n874), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1342gat));
  NOR2_X1   g713(.A1(new_n460), .A2(new_n627), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT117), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n905), .A2(new_n263), .A3(new_n917), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n918), .A2(KEYINPUT56), .ZN(new_n919));
  OAI21_X1  g718(.A(G134gat), .B1(new_n902), .B2(new_n627), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(KEYINPUT56), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(G1343gat));
  NOR3_X1   g721(.A1(new_n725), .A2(new_n435), .A3(new_n460), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n898), .A2(new_n900), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT57), .B1(new_n924), .B2(new_n515), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT115), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n899), .B(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n893), .ZN(new_n928));
  INV_X1    g727(.A(new_n896), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n879), .A2(new_n704), .A3(new_n578), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT119), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n931), .B1(new_n883), .B2(new_n884), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n876), .A2(KEYINPUT119), .A3(new_n702), .A4(new_n878), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n932), .A2(new_n882), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n930), .B1(new_n934), .B2(KEYINPUT120), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT120), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n932), .A2(new_n936), .A3(new_n882), .A4(new_n933), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n929), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n928), .B1(new_n938), .B2(new_n628), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n927), .B1(new_n939), .B2(new_n874), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n515), .A2(KEYINPUT57), .ZN(new_n941));
  OAI22_X1  g740(.A1(new_n925), .A2(KEYINPUT118), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT118), .ZN(new_n943));
  AOI211_X1 g742(.A(new_n943), .B(KEYINPUT57), .C1(new_n924), .C2(new_n515), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n578), .B(new_n923), .C1(new_n942), .C2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n369), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT121), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n725), .A2(new_n730), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n904), .A2(new_n949), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n950), .A2(new_n461), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n951), .A2(new_n339), .A3(new_n578), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n947), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n948), .A2(new_n953), .A3(KEYINPUT58), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT58), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n947), .B(new_n952), .C1(KEYINPUT121), .C2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1344gat));
  INV_X1    g756(.A(KEYINPUT59), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n923), .B1(new_n942), .B2(new_n944), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n958), .B(G148gat), .C1(new_n959), .C2(new_n808), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT122), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n705), .B1(new_n923), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n962), .B1(new_n961), .B2(new_n923), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n891), .B1(new_n938), .B2(new_n628), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(new_n874), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(new_n899), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n730), .A2(KEYINPUT57), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n924), .A2(new_n515), .ZN(new_n968));
  AOI22_X1  g767(.A1(new_n966), .A2(new_n967), .B1(KEYINPUT57), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n337), .B1(new_n963), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n960), .B1(new_n970), .B2(new_n958), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n951), .A2(new_n337), .A3(new_n705), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1345gat));
  OAI21_X1  g772(.A(G155gat), .B1(new_n959), .B2(new_n874), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n951), .A2(new_n672), .A3(new_n748), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1346gat));
  OAI21_X1  g775(.A(G162gat), .B1(new_n959), .B2(new_n627), .ZN(new_n977));
  INV_X1    g776(.A(G162gat), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n950), .A2(new_n978), .A3(new_n917), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(G1347gat));
  AOI21_X1  g779(.A(new_n810), .B1(new_n898), .B2(new_n900), .ZN(new_n981));
  NOR3_X1   g780(.A1(new_n523), .A2(new_n461), .A3(new_n515), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g782(.A(new_n983), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n984), .A2(new_n223), .A3(new_n578), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT124), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n810), .A2(new_n461), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n901), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(KEYINPUT123), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT123), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n901), .A2(new_n990), .A3(new_n987), .ZN(new_n991));
  AND2_X1   g790(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(new_n578), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n986), .B1(new_n993), .B2(G169gat), .ZN(new_n994));
  AOI211_X1 g793(.A(KEYINPUT124), .B(new_n223), .C1(new_n992), .C2(new_n578), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n985), .B1(new_n994), .B2(new_n995), .ZN(G1348gat));
  NAND2_X1  g795(.A1(new_n989), .A2(new_n991), .ZN(new_n997));
  OAI21_X1  g796(.A(G176gat), .B1(new_n997), .B2(new_n808), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n984), .A2(new_n224), .A3(new_n705), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(G1349gat));
  OAI21_X1  g799(.A(G183gat), .B1(new_n997), .B2(new_n874), .ZN(new_n1001));
  INV_X1    g800(.A(new_n214), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n209), .A2(KEYINPUT27), .ZN(new_n1003));
  NOR4_X1   g802(.A1(new_n983), .A2(new_n1002), .A3(new_n1003), .A4(new_n874), .ZN(new_n1004));
  INV_X1    g803(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1006), .A2(KEYINPUT60), .ZN(new_n1007));
  INV_X1    g806(.A(KEYINPUT60), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n1001), .A2(new_n1008), .A3(new_n1005), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1007), .A2(new_n1009), .ZN(G1350gat));
  OR3_X1    g809(.A1(new_n983), .A2(G190gat), .A3(new_n627), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n989), .A2(new_n628), .A3(new_n991), .ZN(new_n1012));
  INV_X1    g811(.A(KEYINPUT61), .ZN(new_n1013));
  AND4_X1   g812(.A1(KEYINPUT125), .A2(new_n1012), .A3(new_n1013), .A4(G190gat), .ZN(new_n1014));
  OAI21_X1  g813(.A(G190gat), .B1(new_n1013), .B2(KEYINPUT125), .ZN(new_n1015));
  INV_X1    g814(.A(new_n1015), .ZN(new_n1016));
  AOI22_X1  g815(.A1(new_n1012), .A2(new_n1016), .B1(KEYINPUT125), .B2(new_n1013), .ZN(new_n1017));
  OAI21_X1  g816(.A(new_n1011), .B1(new_n1014), .B2(new_n1017), .ZN(G1351gat));
  AND3_X1   g817(.A1(new_n981), .A2(new_n460), .A3(new_n949), .ZN(new_n1019));
  AOI21_X1  g818(.A(G197gat), .B1(new_n1019), .B2(new_n578), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n726), .A2(new_n987), .ZN(new_n1021));
  INV_X1    g820(.A(new_n1021), .ZN(new_n1022));
  AND2_X1   g821(.A1(new_n969), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g822(.A1(new_n579), .A2(new_n323), .ZN(new_n1024));
  AOI21_X1  g823(.A(new_n1020), .B1(new_n1023), .B2(new_n1024), .ZN(G1352gat));
  NAND3_X1  g824(.A1(new_n1019), .A2(new_n324), .A3(new_n705), .ZN(new_n1026));
  XOR2_X1   g825(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1027));
  XNOR2_X1  g826(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  AND2_X1   g827(.A1(new_n1023), .A2(new_n705), .ZN(new_n1029));
  OAI21_X1  g828(.A(new_n1028), .B1(new_n1029), .B2(new_n324), .ZN(G1353gat));
  INV_X1    g829(.A(G211gat), .ZN(new_n1031));
  NAND3_X1  g830(.A1(new_n1019), .A2(new_n1031), .A3(new_n748), .ZN(new_n1032));
  NAND2_X1  g831(.A1(new_n1023), .A2(new_n748), .ZN(new_n1033));
  AND3_X1   g832(.A1(new_n1033), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1034));
  AOI21_X1  g833(.A(KEYINPUT63), .B1(new_n1033), .B2(G211gat), .ZN(new_n1035));
  OAI21_X1  g834(.A(new_n1032), .B1(new_n1034), .B2(new_n1035), .ZN(G1354gat));
  AOI21_X1  g835(.A(G218gat), .B1(new_n1019), .B2(new_n628), .ZN(new_n1037));
  NAND2_X1  g836(.A1(new_n628), .A2(G218gat), .ZN(new_n1038));
  XNOR2_X1  g837(.A(new_n1038), .B(KEYINPUT127), .ZN(new_n1039));
  AOI21_X1  g838(.A(new_n1037), .B1(new_n1023), .B2(new_n1039), .ZN(G1355gat));
endmodule


