//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT30), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  OAI211_X1 g004(.A(new_n189), .B(G146), .C1(new_n190), .C2(KEYINPUT1), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(new_n192), .A3(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT67), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT67), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n191), .A2(new_n196), .A3(new_n193), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n192), .A2(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n189), .A2(G146), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n198), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n195), .A2(new_n197), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT11), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G137), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT11), .A3(G134), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n204), .A2(G137), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n205), .A2(new_n207), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n204), .A2(G137), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n206), .A2(G134), .ZN(new_n212));
  OAI21_X1  g026(.A(G131), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G143), .B(G146), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT0), .ZN(new_n216));
  OAI22_X1  g030(.A1(new_n215), .A2(KEYINPUT66), .B1(new_n216), .B2(new_n190), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n199), .A2(new_n200), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n216), .A2(new_n190), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n216), .A2(new_n190), .A3(KEYINPUT65), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n223), .B1(KEYINPUT0), .B2(G128), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n218), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n217), .A2(new_n221), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n205), .A2(new_n209), .A3(new_n207), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G131), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n210), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n202), .A2(new_n214), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n187), .B(new_n188), .C1(new_n230), .C2(KEYINPUT64), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n202), .A2(new_n214), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n226), .A2(new_n229), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT64), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT70), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT30), .B1(new_n230), .B2(new_n187), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n231), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT2), .ZN(new_n240));
  INV_X1    g054(.A(G113), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n242), .A2(new_n243), .B1(KEYINPUT2), .B2(G113), .ZN(new_n244));
  INV_X1    g058(.A(G116), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(G119), .ZN(new_n246));
  INV_X1    g060(.A(G119), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT69), .B1(new_n247), .B2(G116), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(new_n245), .A3(G119), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n246), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n244), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n244), .A2(new_n251), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n238), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n232), .A2(new_n254), .A3(new_n233), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G953), .ZN(new_n260));
  AND2_X1   g074(.A1(KEYINPUT71), .A2(G237), .ZN(new_n261));
  NOR2_X1   g075(.A1(KEYINPUT71), .A2(G237), .ZN(new_n262));
  OAI211_X1 g076(.A(G210), .B(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT26), .B(G101), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n263), .A2(new_n264), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n259), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OR2_X1    g081(.A1(new_n263), .A2(new_n264), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n263), .A2(new_n264), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n258), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n256), .A2(new_n257), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT31), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n232), .A2(new_n254), .A3(new_n233), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n254), .B1(new_n233), .B2(new_n232), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n257), .A2(new_n278), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n271), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n275), .B1(new_n238), .B2(new_n255), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT31), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(new_n284), .A3(new_n272), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n274), .A2(new_n282), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G472), .ZN(new_n287));
  INV_X1    g101(.A(G902), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n289), .B(KEYINPUT73), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT32), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT75), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT29), .ZN(new_n296));
  AOI211_X1 g110(.A(new_n296), .B(new_n271), .C1(new_n257), .C2(new_n278), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n298), .B(KEYINPUT28), .C1(new_n275), .C2(new_n276), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n234), .A2(new_n255), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n257), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n298), .B1(new_n302), .B2(KEYINPUT28), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n288), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n188), .B1(new_n234), .B2(KEYINPUT70), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n187), .B1(new_n230), .B2(KEYINPUT64), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n254), .B1(new_n307), .B2(new_n231), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n271), .B1(new_n308), .B2(new_n275), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n280), .A2(new_n272), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n302), .A2(KEYINPUT28), .ZN(new_n312));
  AOI21_X1  g126(.A(KEYINPUT29), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n304), .B1(new_n309), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n295), .B1(new_n314), .B2(new_n287), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n296), .B1(new_n279), .B2(new_n310), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n256), .A2(new_n257), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(new_n271), .ZN(new_n318));
  OAI211_X1 g132(.A(KEYINPUT75), .B(G472), .C1(new_n318), .C2(new_n304), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n286), .A2(KEYINPUT32), .A3(new_n291), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n294), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(G234), .A2(G237), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(G952), .A3(new_n260), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(G902), .A3(G953), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT21), .B(G898), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n325), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(G214), .B1(G237), .B2(G902), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n251), .A2(KEYINPUT5), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n247), .A2(G116), .ZN(new_n333));
  OAI21_X1  g147(.A(G113), .B1(new_n333), .B2(KEYINPUT5), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G104), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT3), .B1(new_n337), .B2(G107), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n339));
  INV_X1    g153(.A(G107), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n340), .A3(G104), .ZN(new_n341));
  INV_X1    g155(.A(G101), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n337), .A2(G107), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n338), .A2(new_n341), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n337), .A2(G107), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n340), .A2(G104), .ZN(new_n346));
  OAI21_X1  g160(.A(G101), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n244), .A2(new_n251), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n336), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n338), .A2(new_n341), .A3(new_n343), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n353), .A3(G101), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n252), .B2(new_n253), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(G101), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(KEYINPUT4), .A3(new_n344), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n351), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(G110), .B(G122), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  AND2_X1   g175(.A1(KEYINPUT84), .A2(KEYINPUT6), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n359), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n351), .B(new_n360), .C1(new_n355), .C2(new_n358), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n364), .A2(new_n362), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n359), .A2(new_n361), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n363), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G125), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n202), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n226), .A2(G125), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n260), .A2(G224), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n371), .B1(new_n369), .B2(new_n370), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(G902), .B1(new_n367), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT85), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT7), .B1(new_n260), .B2(G224), .ZN(new_n377));
  NOR3_X1   g191(.A1(new_n372), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n334), .B1(new_n251), .B2(KEYINPUT5), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n348), .B1(new_n252), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n351), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n360), .B(KEYINPUT8), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n369), .A2(new_n370), .A3(new_n377), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n376), .B1(new_n378), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n373), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n388));
  INV_X1    g202(.A(new_n377), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n390), .A2(KEYINPUT85), .A3(new_n384), .A4(new_n383), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n386), .A2(new_n391), .A3(new_n364), .ZN(new_n392));
  OAI21_X1  g206(.A(G210), .B1(G237), .B2(G902), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n375), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n375), .B2(new_n392), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n330), .B(new_n331), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G469), .ZN(new_n397));
  XNOR2_X1  g211(.A(G110), .B(G140), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n260), .A2(G227), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n201), .A2(KEYINPUT81), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT81), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n215), .A2(new_n402), .A3(new_n198), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n401), .A2(new_n403), .A3(new_n191), .A4(new_n193), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n349), .ZN(new_n405));
  XOR2_X1   g219(.A(KEYINPUT82), .B(KEYINPUT10), .Z(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n229), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n357), .A2(new_n226), .A3(new_n354), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n202), .A2(new_n349), .A3(KEYINPUT10), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n408), .A2(new_n409), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n348), .A2(new_n197), .A3(new_n195), .A4(new_n201), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n405), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(KEYINPUT12), .B1(new_n414), .B2(new_n229), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT12), .ZN(new_n416));
  AOI211_X1 g230(.A(new_n416), .B(new_n409), .C1(new_n405), .C2(new_n413), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n400), .B(new_n412), .C1(new_n415), .C2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n194), .B1(KEYINPUT81), .B2(new_n201), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n348), .B1(new_n419), .B2(new_n403), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n410), .B(new_n411), .C1(new_n420), .C2(new_n406), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n229), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n400), .B1(new_n422), .B2(new_n412), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT83), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n418), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI211_X1 g239(.A(KEYINPUT83), .B(new_n400), .C1(new_n422), .C2(new_n412), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n397), .B(new_n288), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n397), .A2(new_n288), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n412), .B1(new_n415), .B2(new_n417), .ZN(new_n429));
  XOR2_X1   g243(.A(new_n400), .B(KEYINPUT80), .Z(new_n430));
  AND2_X1   g244(.A1(new_n412), .A2(new_n400), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n429), .A2(new_n430), .B1(new_n431), .B2(new_n422), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n428), .B1(new_n432), .B2(G469), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT9), .B(G234), .ZN(new_n435));
  OAI21_X1  g249(.A(G221), .B1(new_n435), .B2(G902), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AND2_X1   g251(.A1(KEYINPUT86), .A2(G143), .ZN(new_n438));
  NOR2_X1   g252(.A1(KEYINPUT86), .A2(G143), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OR2_X1    g254(.A1(KEYINPUT71), .A2(G237), .ZN(new_n441));
  NAND2_X1  g255(.A1(KEYINPUT71), .A2(G237), .ZN(new_n442));
  AOI21_X1  g256(.A(G953), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n440), .B1(new_n443), .B2(G214), .ZN(new_n444));
  OAI211_X1 g258(.A(G214), .B(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(new_n439), .ZN(new_n446));
  OAI21_X1  g260(.A(G131), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT17), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT86), .B(G143), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT71), .B(G237), .ZN(new_n451));
  INV_X1    g265(.A(new_n439), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n451), .A2(G214), .A3(new_n260), .A4(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n450), .A2(new_n453), .A3(new_n208), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n447), .A2(new_n448), .A3(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(G125), .B(G140), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT77), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT16), .ZN(new_n458));
  INV_X1    g272(.A(G140), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(G125), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n456), .A2(KEYINPUT16), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT77), .A4(G125), .ZN(new_n462));
  AOI21_X1  g276(.A(G146), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n459), .A2(G125), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n368), .A2(G140), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT16), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n460), .A2(new_n457), .ZN(new_n467));
  AND4_X1   g281(.A1(G146), .A2(new_n466), .A3(new_n467), .A4(new_n462), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n450), .A2(new_n453), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(KEYINPUT17), .A3(G131), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n455), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(G113), .B(G122), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(new_n337), .ZN(new_n474));
  NAND2_X1  g288(.A1(KEYINPUT18), .A2(G131), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n450), .A2(new_n453), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n464), .A2(new_n465), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G146), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n456), .A2(new_n192), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT87), .ZN(new_n482));
  INV_X1    g296(.A(new_n475), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n482), .B1(new_n470), .B2(new_n483), .ZN(new_n484));
  AOI211_X1 g298(.A(KEYINPUT87), .B(new_n475), .C1(new_n450), .C2(new_n453), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n481), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n472), .A2(new_n474), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n474), .B1(new_n472), .B2(new_n486), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n288), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(G475), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT20), .ZN(new_n491));
  INV_X1    g305(.A(new_n474), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n476), .A2(new_n480), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n470), .A2(new_n483), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT87), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n470), .A2(new_n482), .A3(new_n483), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n456), .A2(KEYINPUT19), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n456), .A2(KEYINPUT19), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n192), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n461), .A2(G146), .A3(new_n462), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n502), .B1(new_n447), .B2(new_n454), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n492), .B1(new_n497), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n472), .A2(new_n474), .A3(new_n486), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(G475), .A2(G902), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n491), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n507), .ZN(new_n509));
  AOI211_X1 g323(.A(KEYINPUT20), .B(new_n509), .C1(new_n504), .C2(new_n505), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n490), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(G128), .B(G143), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(new_n204), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n245), .A2(KEYINPUT14), .A3(G122), .ZN(new_n515));
  XNOR2_X1  g329(.A(G116), .B(G122), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(G107), .B(new_n515), .C1(new_n517), .C2(KEYINPUT14), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n514), .B(new_n518), .C1(G107), .C2(new_n517), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n513), .A2(KEYINPUT13), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n189), .A2(G128), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n520), .B(G134), .C1(KEYINPUT13), .C2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n516), .B(new_n340), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n513), .A2(new_n204), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G217), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n435), .A2(new_n526), .A3(G953), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n519), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n527), .B1(new_n519), .B2(new_n525), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n288), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G478), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(KEYINPUT15), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n530), .B(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n512), .A2(new_n534), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n396), .A2(new_n437), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n526), .B1(G234), .B2(new_n288), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n190), .A2(G119), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n247), .A2(G128), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT24), .B(G110), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT23), .B1(new_n190), .B2(G119), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(KEYINPUT76), .A3(new_n539), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT76), .B1(new_n247), .B2(G128), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n247), .A2(G128), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(KEYINPUT23), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n543), .B1(new_n549), .B2(G110), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n463), .B2(new_n468), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n541), .A2(new_n542), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(new_n549), .B2(G110), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(new_n501), .A3(new_n479), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n260), .A2(G221), .A3(G234), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(KEYINPUT22), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(new_n206), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n558), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(new_n551), .A3(new_n554), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n288), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n538), .B1(new_n562), .B2(KEYINPUT25), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT78), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT25), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n559), .A2(new_n565), .A3(new_n561), .A4(new_n288), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n564), .B1(new_n563), .B2(new_n566), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n537), .A2(G902), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(KEYINPUT79), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n559), .A2(new_n561), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n322), .A2(new_n536), .A3(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(G101), .ZN(G3));
  INV_X1    g390(.A(new_n292), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n577), .A2(new_n437), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n287), .B1(new_n286), .B2(new_n288), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(new_n573), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n530), .A2(new_n531), .ZN(new_n582));
  XOR2_X1   g396(.A(KEYINPUT88), .B(KEYINPUT33), .Z(new_n583));
  OR3_X1    g397(.A1(new_n528), .A2(new_n529), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(KEYINPUT88), .A2(KEYINPUT33), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n585), .B1(new_n528), .B2(new_n529), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n288), .A2(G478), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n582), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n511), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n396), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n581), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(KEYINPUT34), .B(G104), .Z(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(G6));
  INV_X1    g408(.A(new_n331), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n375), .A2(new_n392), .ZN(new_n596));
  INV_X1    g410(.A(new_n393), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n375), .A2(new_n392), .A3(new_n393), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n595), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n512), .A2(KEYINPUT89), .A3(new_n330), .A4(new_n533), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT89), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n490), .B(new_n533), .C1(new_n508), .C2(new_n510), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n602), .B1(new_n603), .B2(new_n329), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n600), .A2(new_n601), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n581), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT35), .B(G107), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G9));
  INV_X1    g422(.A(new_n568), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n558), .A2(KEYINPUT36), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n555), .B(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT90), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n611), .A2(new_n612), .A3(new_n571), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n612), .B1(new_n611), .B2(new_n571), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n609), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n617), .A2(new_n434), .A3(new_n436), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n618), .A2(new_n396), .A3(new_n535), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n286), .A2(new_n288), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(G472), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n619), .A2(new_n292), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT37), .B(G110), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G12));
  AND3_X1   g438(.A1(new_n286), .A2(KEYINPUT32), .A3(new_n291), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT32), .B1(new_n286), .B2(new_n291), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n618), .B1(new_n627), .B2(new_n320), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT92), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n324), .B(KEYINPUT91), .Z(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(G900), .B2(new_n326), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n603), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n600), .A2(new_n629), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n629), .B1(new_n600), .B2(new_n633), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n628), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G128), .ZN(G30));
  NOR2_X1   g452(.A1(new_n394), .A2(new_n395), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT38), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n512), .A2(new_n534), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n617), .A2(new_n595), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n273), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n277), .A2(new_n272), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT93), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n288), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(G472), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n627), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT94), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n644), .A2(KEYINPUT94), .A3(new_n650), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n631), .B(KEYINPUT39), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n434), .A2(new_n436), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT95), .B(KEYINPUT40), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n653), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G143), .ZN(G45));
  NAND3_X1  g474(.A1(new_n511), .A2(new_n589), .A3(new_n631), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT96), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT96), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n511), .A2(new_n589), .A3(new_n663), .A4(new_n631), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n665), .A2(new_n595), .A3(new_n639), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n628), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT97), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(new_n192), .ZN(G48));
  OAI21_X1  g483(.A(new_n288), .B1(new_n425), .B2(new_n426), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(G469), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n436), .A3(new_n427), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT98), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n671), .A2(KEYINPUT98), .A3(new_n436), .A4(new_n427), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n676), .A2(new_n322), .A3(new_n574), .A4(new_n591), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT41), .B(G113), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G15));
  NAND4_X1  g493(.A1(new_n676), .A2(new_n322), .A3(new_n605), .A4(new_n574), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G116), .ZN(G18));
  AND3_X1   g495(.A1(new_n674), .A2(new_n600), .A3(new_n675), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n617), .A2(new_n330), .A3(new_n534), .A4(new_n512), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n682), .A2(new_n322), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G119), .ZN(G21));
  NAND2_X1  g500(.A1(new_n299), .A2(new_n280), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n271), .B1(new_n687), .B2(new_n303), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n274), .A2(new_n285), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n291), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n691), .A2(new_n579), .A3(new_n573), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n600), .A2(new_n330), .A3(new_n642), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n676), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G122), .ZN(G24));
  NAND2_X1  g509(.A1(new_n690), .A2(new_n617), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n665), .A2(new_n696), .A3(new_n579), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT99), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n682), .A3(new_n698), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n291), .A2(new_n689), .B1(new_n569), .B2(new_n615), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n621), .A2(new_n700), .A3(new_n664), .A4(new_n662), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n674), .A2(new_n600), .A3(new_n675), .ZN(new_n702));
  OAI21_X1  g516(.A(KEYINPUT99), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT100), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n368), .ZN(G27));
  INV_X1    g520(.A(new_n665), .ZN(new_n707));
  INV_X1    g521(.A(new_n436), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n595), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n598), .A2(new_n599), .A3(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT101), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n427), .A2(new_n433), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n434), .A2(KEYINPUT101), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n710), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n707), .A2(new_n714), .A3(KEYINPUT42), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n322), .A2(new_n574), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT102), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n322), .A2(KEYINPUT102), .A3(new_n574), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n715), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n322), .A2(new_n707), .A3(new_n574), .A4(new_n714), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT42), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n208), .ZN(G33));
  NAND4_X1  g540(.A1(new_n322), .A2(new_n714), .A3(new_n574), .A4(new_n633), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G134), .ZN(G36));
  OAI21_X1  g542(.A(G469), .B1(new_n432), .B2(KEYINPUT45), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n429), .A2(new_n430), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n431), .A2(new_n422), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n730), .A2(new_n731), .A3(KEYINPUT45), .ZN(new_n732));
  OAI22_X1  g546(.A1(new_n729), .A2(new_n732), .B1(new_n397), .B2(new_n288), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n734), .A2(KEYINPUT46), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n427), .B1(new_n734), .B2(KEYINPUT46), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n436), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n738), .A2(new_n655), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n617), .B1(new_n577), .B2(new_n579), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT43), .B1(new_n512), .B2(new_n589), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT103), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n511), .B(new_n742), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n589), .A2(KEYINPUT43), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n746), .A2(KEYINPUT44), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(KEYINPUT44), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n598), .A2(new_n331), .A3(new_n599), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n739), .A2(new_n747), .A3(new_n748), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT104), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n206), .ZN(G39));
  OR4_X1    g567(.A1(new_n574), .A2(new_n322), .A3(new_n665), .A4(new_n749), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  XOR2_X1   g569(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n756));
  OR2_X1    g570(.A1(new_n737), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n737), .B1(KEYINPUT105), .B2(KEYINPUT47), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n755), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT106), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(new_n459), .ZN(G42));
  NOR2_X1   g575(.A1(G952), .A2(G953), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n631), .A2(new_n436), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n617), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n765), .A2(new_n600), .A3(new_n642), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n713), .A2(new_n712), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI22_X1  g582(.A1(new_n628), .A2(new_n666), .B1(new_n650), .B2(new_n768), .ZN(new_n769));
  AND4_X1   g583(.A1(KEYINPUT52), .A2(new_n704), .A3(new_n769), .A4(new_n637), .ZN(new_n770));
  AOI22_X1  g584(.A1(new_n699), .A2(new_n703), .B1(new_n628), .B2(new_n636), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT52), .B1(new_n771), .B2(new_n769), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n396), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n590), .A2(KEYINPUT108), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT108), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n776), .B1(new_n511), .B2(new_n589), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n578), .A2(new_n580), .A3(new_n774), .A4(new_n778), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n575), .A2(new_n779), .A3(KEYINPUT109), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT109), .B1(new_n575), .B2(new_n779), .ZN(new_n781));
  INV_X1    g595(.A(new_n603), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n578), .A2(new_n580), .A3(new_n774), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n622), .A2(new_n783), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n780), .A2(new_n781), .A3(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n677), .A2(new_n685), .A3(new_n680), .A4(new_n694), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n511), .A2(new_n533), .A3(new_n632), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n750), .A2(KEYINPUT110), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n618), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT110), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n512), .A2(new_n534), .A3(new_n631), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n792), .B1(new_n749), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n322), .A2(new_n790), .A3(new_n791), .A4(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n696), .A2(new_n579), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(new_n707), .A3(new_n714), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(new_n727), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n715), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n322), .A2(KEYINPUT102), .A3(new_n574), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT102), .B1(new_n322), .B2(new_n574), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n798), .B1(new_n802), .B2(new_n723), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n785), .A2(new_n788), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n763), .B1(new_n773), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n698), .B1(new_n697), .B2(new_n682), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n701), .A2(new_n702), .A3(KEYINPUT99), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n637), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n769), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n806), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n771), .A2(KEYINPUT52), .A3(new_n769), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n683), .B1(new_n627), .B2(new_n320), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n621), .A2(new_n574), .A3(new_n690), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n674), .A2(new_n675), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n682), .A2(new_n814), .B1(new_n817), .B2(new_n693), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n818), .A2(KEYINPUT53), .A3(new_n677), .A4(new_n680), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n575), .A2(new_n779), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT109), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n575), .A2(new_n779), .A3(KEYINPUT109), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n622), .A2(new_n783), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n819), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n813), .A2(new_n826), .A3(KEYINPUT111), .A4(new_n803), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n805), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT107), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n818), .A2(new_n830), .A3(new_n677), .A4(new_n680), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n786), .A2(KEYINPUT107), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n785), .A2(new_n803), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n787), .B1(new_n773), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n828), .A2(new_n829), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT53), .B1(new_n773), .B2(new_n833), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n785), .A2(new_n831), .A3(new_n832), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(new_n813), .A3(new_n787), .A4(new_n803), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n836), .A2(new_n838), .A3(KEYINPUT54), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n745), .A2(new_n630), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n817), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n600), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n843), .B(KEYINPUT114), .Z(new_n844));
  NOR3_X1   g658(.A1(new_n650), .A2(new_n573), .A3(new_n324), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n816), .A2(new_n749), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g661(.A(G952), .B(new_n260), .C1(new_n847), .C2(new_n590), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n641), .A2(new_n331), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n842), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT50), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n841), .A2(new_n846), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n796), .ZN(new_n855));
  INV_X1    g669(.A(new_n589), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n845), .A2(new_n512), .A3(new_n856), .A4(new_n846), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n671), .A2(new_n427), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n436), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n757), .B2(new_n758), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n841), .A2(new_n692), .A3(new_n750), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n855), .B(new_n857), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n850), .B1(new_n853), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n718), .A2(new_n719), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n854), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT48), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n849), .A2(new_n863), .A3(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n857), .A2(KEYINPUT112), .A3(new_n855), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT112), .B1(new_n857), .B2(new_n855), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT113), .ZN(new_n871));
  OR3_X1    g685(.A1(new_n870), .A2(new_n871), .A3(new_n853), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n871), .B1(new_n870), .B2(new_n853), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n860), .A2(new_n861), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n850), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n867), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n762), .B1(new_n840), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n858), .B(KEYINPUT49), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n743), .A2(new_n574), .A3(new_n589), .A4(new_n709), .ZN(new_n880));
  NOR4_X1   g694(.A1(new_n650), .A2(new_n641), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n878), .A2(new_n881), .ZN(G75));
  NOR2_X1   g696(.A1(new_n260), .A2(G952), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n773), .A2(new_n804), .A3(new_n763), .ZN(new_n885));
  INV_X1    g699(.A(new_n798), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n886), .B1(new_n720), .B2(new_n724), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n887), .A2(new_n819), .A3(new_n825), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT111), .B1(new_n888), .B2(new_n813), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n834), .B1(new_n885), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(G210), .A3(G902), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT56), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n367), .B(new_n374), .Z(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT55), .Z(new_n895));
  OAI21_X1  g709(.A(new_n884), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT115), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n893), .A2(new_n897), .A3(new_n895), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n288), .B1(new_n828), .B2(new_n834), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT56), .B1(new_n899), .B2(G210), .ZN(new_n900));
  INV_X1    g714(.A(new_n895), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT115), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n896), .B1(new_n898), .B2(new_n902), .ZN(G51));
  NAND2_X1  g717(.A1(new_n890), .A2(KEYINPUT54), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n835), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n428), .B(KEYINPUT57), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n425), .A2(new_n426), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT116), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n729), .A2(new_n732), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n899), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n910), .B1(new_n899), .B2(new_n911), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n883), .B1(new_n909), .B2(new_n914), .ZN(G54));
  NAND2_X1  g729(.A1(KEYINPUT58), .A2(G475), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n890), .A2(G902), .A3(new_n506), .A4(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT117), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n899), .A2(KEYINPUT117), .A3(new_n506), .A4(new_n917), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n883), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI211_X1 g736(.A(new_n288), .B(new_n916), .C1(new_n828), .C2(new_n834), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT118), .B1(new_n923), .B2(new_n506), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n890), .A2(G902), .A3(new_n917), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT118), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n925), .A2(new_n926), .A3(new_n505), .A4(new_n504), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n922), .A2(new_n928), .ZN(G60));
  NAND2_X1  g743(.A1(G478), .A2(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT59), .Z(new_n931));
  OAI211_X1 g745(.A(KEYINPUT119), .B(new_n587), .C1(new_n840), .C2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n587), .A2(new_n931), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n883), .B1(new_n905), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT119), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n931), .B1(new_n835), .B2(new_n839), .ZN(new_n936));
  INV_X1    g750(.A(new_n587), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n932), .A2(new_n934), .A3(new_n938), .ZN(G63));
  NAND2_X1  g753(.A1(G217), .A2(G902), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT120), .Z(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT60), .Z(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n828), .B2(new_n834), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n559), .A2(new_n561), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n883), .B1(new_n944), .B2(new_n611), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT121), .B1(new_n944), .B2(new_n611), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n950), .A2(KEYINPUT61), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n947), .B(new_n948), .C1(new_n950), .C2(KEYINPUT61), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(G66));
  NAND3_X1  g768(.A1(new_n785), .A2(new_n831), .A3(new_n832), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n260), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT122), .Z(new_n957));
  INV_X1    g771(.A(G224), .ZN(new_n958));
  OAI21_X1  g772(.A(G953), .B1(new_n328), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(G898), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n367), .B1(new_n961), .B2(G953), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n960), .B(new_n962), .Z(G69));
  NOR2_X1   g777(.A1(new_n498), .A2(new_n499), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n238), .B(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(G900), .B2(G953), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n727), .B1(new_n720), .B2(new_n724), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT125), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n771), .A2(new_n667), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n739), .A2(new_n600), .A3(new_n642), .A4(new_n864), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n970), .A2(new_n759), .A3(new_n751), .A4(new_n971), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n968), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n966), .B1(new_n973), .B2(G953), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n970), .A2(new_n659), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(KEYINPUT62), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT62), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n970), .A2(new_n659), .A3(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n778), .A2(new_n782), .ZN(new_n979));
  OR4_X1    g793(.A1(new_n716), .A2(new_n979), .A3(new_n656), .A4(new_n749), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n759), .A2(new_n751), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n976), .A2(new_n978), .A3(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT123), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n976), .A2(KEYINPUT123), .A3(new_n978), .A4(new_n981), .ZN(new_n985));
  AOI21_X1  g799(.A(G953), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n965), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n974), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n260), .B1(G227), .B2(G900), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT124), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n989), .B1(new_n974), .B2(new_n990), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n988), .A2(new_n991), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n992), .A2(new_n993), .ZN(G72));
  NAND2_X1  g808(.A1(G472), .A2(G902), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT63), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT126), .Z(new_n997));
  OAI21_X1  g811(.A(new_n997), .B1(new_n973), .B2(new_n955), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n998), .A2(new_n271), .A3(new_n283), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n309), .A2(KEYINPUT127), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n1000), .A2(new_n645), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n309), .A2(KEYINPUT127), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n996), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n836), .A2(new_n838), .A3(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n999), .A2(new_n884), .A3(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n984), .A2(new_n837), .A3(new_n985), .ZN(new_n1006));
  AOI211_X1 g820(.A(new_n271), .B(new_n283), .C1(new_n1006), .C2(new_n997), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1005), .A2(new_n1007), .ZN(G57));
endmodule


