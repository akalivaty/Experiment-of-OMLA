//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(new_n214), .A2(KEYINPUT0), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n219), .B1(KEYINPUT0), .B2(new_n214), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT64), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n211), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n221), .A2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  NAND2_X1  g0038(.A1(G68), .A2(G77), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n203), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT65), .ZN(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  NAND2_X1  g0047(.A1(new_n208), .A2(G274), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G41), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT66), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT66), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n249), .B1(new_n254), .B2(G45), .ZN(new_n255));
  INV_X1    g0055(.A(G226), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n255), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(G222), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n262), .A2(G223), .A3(G1698), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n264), .B(new_n265), .C1(new_n202), .C2(new_n262), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT67), .ZN(new_n267));
  OR2_X1    g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n258), .B1(new_n266), .B2(new_n267), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n261), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(G179), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(G50), .ZN(new_n274));
  NAND3_X1  g0074(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n275), .A2(new_n215), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n276), .B1(G1), .B2(new_n209), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n274), .B1(new_n278), .B2(G50), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT68), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G58), .ZN(new_n282));
  XNOR2_X1  g0082(.A(new_n282), .B(KEYINPUT8), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n209), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G150), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT69), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n286), .A2(KEYINPUT69), .A3(new_n288), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G50), .A2(G58), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n209), .B1(new_n293), .B2(new_n201), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT70), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n291), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n275), .A2(new_n215), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n280), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n270), .A2(G169), .ZN(new_n299));
  NOR3_X1   g0099(.A1(new_n272), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n296), .A2(new_n297), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n279), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT9), .ZN(new_n303));
  INV_X1    g0103(.A(G200), .ZN(new_n304));
  OAI22_X1  g0104(.A1(new_n302), .A2(new_n303), .B1(new_n304), .B2(new_n270), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n298), .A2(KEYINPUT9), .B1(new_n271), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT10), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n302), .A2(new_n303), .B1(G190), .B2(new_n270), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n298), .A2(KEYINPUT9), .B1(new_n271), .B2(G200), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT10), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n300), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT17), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n262), .A2(G223), .A3(new_n263), .ZN(new_n315));
  INV_X1    g0115(.A(G33), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT3), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT3), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G33), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n317), .A2(new_n319), .A3(G226), .A4(G1698), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G33), .A2(G87), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n315), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT76), .ZN(new_n323));
  INV_X1    g0123(.A(new_n258), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n323), .B1(new_n322), .B2(new_n324), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT77), .ZN(new_n328));
  INV_X1    g0128(.A(G232), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n260), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT66), .B(G41), .ZN(new_n331));
  INV_X1    g0131(.A(G45), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n248), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n328), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n255), .B(KEYINPUT77), .C1(new_n329), .C2(new_n260), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n334), .A2(new_n335), .A3(new_n306), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n322), .A2(new_n324), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n338), .A2(new_n334), .A3(new_n335), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n327), .A2(new_n337), .B1(new_n304), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n283), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n273), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n277), .A2(new_n283), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G58), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(new_n201), .ZN(new_n346));
  NOR2_X1   g0146(.A1(G58), .A2(G68), .ZN(new_n347));
  OAI21_X1  g0147(.A(G20), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n287), .A2(G159), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n317), .A2(new_n319), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n209), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n354), .A2(G20), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n353), .A2(new_n354), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  OAI211_X1 g0156(.A(KEYINPUT16), .B(new_n351), .C1(new_n356), .C2(new_n201), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n297), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT75), .ZN(new_n359));
  AND3_X1   g0159(.A1(new_n317), .A2(new_n319), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n316), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n355), .ZN(new_n362));
  AOI21_X1  g0162(.A(G20), .B1(new_n317), .B2(new_n319), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n360), .A2(new_n362), .B1(new_n363), .B2(KEYINPUT7), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G68), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT16), .B1(new_n365), .B2(new_n351), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n344), .B1(new_n358), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n314), .B1(new_n340), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G169), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n339), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n338), .A2(KEYINPUT76), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G179), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n334), .A2(new_n335), .A3(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n370), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n344), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n354), .B1(new_n262), .B2(G20), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n352), .A2(new_n355), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n350), .B1(new_n380), .B2(G68), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n276), .B1(new_n381), .B2(KEYINPUT16), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT16), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n355), .B(new_n361), .C1(new_n352), .C2(KEYINPUT75), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n201), .B1(new_n384), .B2(new_n378), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n383), .B1(new_n385), .B2(new_n350), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n377), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT18), .B1(new_n376), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n375), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n327), .A2(new_n389), .B1(new_n369), .B2(new_n339), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT18), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n367), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n339), .A2(new_n304), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n373), .B2(new_n336), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n394), .A2(new_n387), .A3(KEYINPUT17), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n368), .A2(new_n388), .A3(new_n392), .A4(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT8), .B(G58), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n399), .A2(new_n287), .B1(G20), .B2(G77), .ZN(new_n400));
  XNOR2_X1  g0200(.A(KEYINPUT15), .B(G87), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n285), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n276), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n273), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n202), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n277), .B2(new_n202), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n262), .A2(G232), .A3(new_n263), .ZN(new_n409));
  INV_X1    g0209(.A(G107), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n409), .B1(new_n410), .B2(new_n262), .ZN(new_n411));
  INV_X1    g0211(.A(G238), .ZN(new_n412));
  NOR3_X1   g0212(.A1(new_n352), .A2(new_n412), .A3(new_n263), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n324), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n260), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n333), .B1(G244), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n408), .B1(new_n417), .B2(new_n369), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(G179), .B2(new_n417), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(G200), .ZN(new_n420));
  OR3_X1    g0220(.A1(new_n404), .A2(KEYINPUT71), .A3(new_n407), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n414), .A2(G190), .A3(new_n416), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT71), .B1(new_n407), .B2(new_n404), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n420), .A2(new_n421), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT72), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n255), .B1(new_n412), .B2(new_n260), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n256), .A2(new_n263), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n329), .A2(G1698), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n317), .A2(new_n429), .A3(new_n319), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G97), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n258), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT13), .B1(new_n428), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n432), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n324), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT13), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n415), .A2(G238), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n436), .A2(new_n437), .A3(new_n255), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(G169), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT14), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT14), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n440), .A2(new_n443), .A3(G169), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n442), .B(new_n444), .C1(new_n374), .C2(new_n440), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n287), .A2(G50), .B1(G20), .B2(new_n201), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n202), .B2(new_n284), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n447), .A2(KEYINPUT11), .A3(new_n297), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT12), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n449), .B1(new_n405), .B2(new_n201), .ZN(new_n450));
  NOR3_X1   g0250(.A1(new_n273), .A2(KEYINPUT12), .A3(G68), .ZN(new_n451));
  OAI22_X1  g0251(.A1(new_n277), .A2(new_n201), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT11), .B1(new_n447), .B2(new_n297), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n448), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n445), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n419), .A2(KEYINPUT72), .A3(new_n424), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n427), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n434), .A2(new_n439), .A3(G190), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n459), .A2(new_n454), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT73), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n461), .B1(new_n440), .B2(G200), .ZN(new_n462));
  AOI211_X1 g0262(.A(KEYINPUT73), .B(new_n304), .C1(new_n434), .C2(new_n439), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT74), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n460), .B(KEYINPUT74), .C1(new_n463), .C2(new_n462), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AND4_X1   g0268(.A1(new_n313), .A2(new_n397), .A3(new_n458), .A4(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT80), .ZN(new_n471));
  INV_X1    g0271(.A(G97), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n405), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n208), .A2(G33), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n276), .A2(new_n474), .A3(new_n273), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n473), .B1(new_n476), .B2(new_n472), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n364), .A2(G107), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT78), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT6), .ZN(new_n480));
  AND2_X1   g0280(.A1(G97), .A2(G107), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n480), .B1(new_n481), .B2(new_n205), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n410), .A2(KEYINPUT6), .A3(G97), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n209), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n287), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(new_n202), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n479), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n486), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n410), .A2(KEYINPUT6), .A3(G97), .ZN(new_n489));
  XNOR2_X1  g0289(.A(G97), .B(G107), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(new_n480), .ZN(new_n491));
  OAI211_X1 g0291(.A(KEYINPUT78), .B(new_n488), .C1(new_n491), .C2(new_n209), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n478), .A2(new_n487), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n297), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT79), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT79), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n493), .A2(new_n496), .A3(new_n297), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n477), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n317), .A2(new_n319), .A3(G244), .A4(new_n263), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n262), .A2(KEYINPUT4), .A3(G244), .A4(new_n263), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n262), .A2(G250), .A3(G1698), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G283), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n501), .A2(new_n502), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT5), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n208), .B(G45), .C1(new_n506), .C2(G41), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n507), .B1(new_n254), .B2(new_n506), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(new_n324), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n505), .A2(new_n324), .B1(new_n509), .B2(G257), .ZN(new_n510));
  INV_X1    g0310(.A(G274), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n324), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n508), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n510), .A2(new_n374), .A3(new_n513), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n510), .A2(new_n513), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n514), .B1(new_n515), .B2(G169), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n471), .B1(new_n498), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n477), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n493), .A2(new_n496), .A3(new_n297), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n496), .B1(new_n493), .B2(new_n297), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n510), .A2(new_n374), .A3(new_n513), .ZN(new_n522));
  AOI21_X1  g0322(.A(G169), .B1(new_n510), .B2(new_n513), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n521), .A2(KEYINPUT80), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n510), .A2(new_n513), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G200), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n515), .A2(G190), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n498), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n517), .A2(new_n525), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n475), .A2(G116), .ZN(new_n531));
  INV_X1    g0331(.A(G116), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n405), .A2(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n275), .A2(new_n215), .B1(G20), .B2(new_n532), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n504), .B(new_n209), .C1(G33), .C2(new_n472), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT20), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n534), .A2(KEYINPUT20), .A3(new_n535), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n531), .B(new_n533), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT5), .B1(new_n251), .B2(new_n253), .ZN(new_n540));
  OAI211_X1 g0340(.A(G270), .B(new_n258), .C1(new_n540), .C2(new_n507), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT81), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n332), .A2(G1), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n250), .A2(KEYINPUT5), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n543), .B(new_n544), .C1(new_n331), .C2(KEYINPUT5), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT81), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(G270), .A4(new_n258), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n317), .A2(new_n319), .A3(G264), .A4(G1698), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n317), .A2(new_n319), .A3(G257), .A4(new_n263), .ZN(new_n550));
  INV_X1    g0350(.A(G303), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n549), .B(new_n550), .C1(new_n551), .C2(new_n262), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n324), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n513), .ZN(new_n554));
  OAI211_X1 g0354(.A(KEYINPUT21), .B(G169), .C1(new_n548), .C2(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n552), .A2(new_n324), .B1(new_n508), .B2(new_n512), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n556), .A2(G179), .A3(new_n542), .A4(new_n547), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n539), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n538), .B(G169), .C1(new_n548), .C2(new_n554), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT21), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT82), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT82), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n559), .A2(new_n563), .A3(new_n560), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n558), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n262), .A2(new_n209), .A3(G68), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT19), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n209), .B1(new_n432), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(G87), .B2(new_n206), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n567), .B1(new_n284), .B2(new_n472), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n566), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n297), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n401), .A2(new_n405), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n572), .B(new_n573), .C1(new_n476), .C2(new_n401), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n543), .A2(new_n511), .ZN(new_n575));
  INV_X1    g0375(.A(G250), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n332), .B2(G1), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n575), .A2(new_n258), .A3(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n317), .A2(new_n319), .A3(G238), .A4(new_n263), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n317), .A2(new_n319), .A3(G244), .A4(G1698), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n579), .B(new_n580), .C1(new_n316), .C2(new_n532), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n578), .B1(new_n581), .B2(new_n324), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n374), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n574), .B(new_n583), .C1(G169), .C2(new_n582), .ZN(new_n584));
  OR2_X1    g0384(.A1(new_n582), .A2(new_n304), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n475), .A2(G87), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n572), .A2(new_n573), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n582), .A2(G190), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT25), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n273), .B2(G107), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n273), .A2(new_n591), .A3(G107), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT84), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(KEYINPUT84), .B(new_n591), .C1(new_n273), .C2(G107), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n595), .A2(new_n596), .B1(new_n475), .B2(G107), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n317), .A2(new_n319), .A3(new_n209), .A4(G87), .ZN(new_n599));
  XOR2_X1   g0399(.A(KEYINPUT83), .B(KEYINPUT22), .Z(new_n600));
  XNOR2_X1  g0400(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NOR3_X1   g0401(.A1(new_n316), .A2(new_n532), .A3(G20), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT23), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n209), .B2(G107), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n410), .A2(KEYINPUT23), .A3(G20), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n602), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(KEYINPUT24), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT24), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n601), .A2(new_n609), .A3(new_n606), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n598), .B1(new_n611), .B2(new_n297), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n545), .A2(G264), .A3(new_n258), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n613), .A2(new_n513), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n262), .A2(G257), .A3(G1698), .ZN(new_n615));
  NAND2_X1  g0415(.A1(G33), .A2(G294), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n317), .A2(new_n319), .A3(G250), .A4(new_n263), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n324), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n614), .A2(G190), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n513), .A3(new_n613), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G200), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n590), .B1(new_n612), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n612), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT85), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n626), .B1(new_n621), .B2(G169), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT86), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n621), .B2(new_n374), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n614), .A2(KEYINPUT86), .A3(G179), .A4(new_n619), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n621), .A2(new_n626), .A3(G169), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n628), .A2(new_n630), .A3(new_n631), .A4(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n625), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n542), .A2(new_n547), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n556), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n538), .B1(new_n636), .B2(G200), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n306), .B2(new_n636), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n565), .A2(new_n624), .A3(new_n634), .A4(new_n638), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n470), .A2(new_n530), .A3(new_n639), .ZN(G372));
  INV_X1    g0440(.A(new_n419), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n455), .A2(new_n445), .B1(new_n641), .B2(new_n464), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n368), .A2(new_n395), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n388), .B(new_n392), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n308), .A2(new_n312), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n300), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n555), .A2(new_n557), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n538), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n559), .A2(new_n563), .A3(new_n560), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n563), .B1(new_n559), .B2(new_n560), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n630), .A2(new_n631), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n621), .A2(new_n626), .A3(G169), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(new_n627), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n612), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n624), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n584), .B1(new_n656), .B2(new_n530), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n498), .A2(new_n516), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n584), .A2(new_n589), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n590), .B1(new_n517), .B2(new_n525), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n661), .B1(new_n662), .B2(new_n659), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n646), .B1(new_n470), .B2(new_n664), .ZN(G369));
  INV_X1    g0465(.A(G13), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n666), .A2(G1), .A3(G20), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT27), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT87), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n667), .A2(KEYINPUT87), .A3(new_n668), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G213), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(new_n667), .B2(new_n668), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G343), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n538), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(KEYINPUT88), .B1(new_n651), .B2(new_n679), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n638), .B(new_n648), .C1(new_n649), .C2(new_n650), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n680), .B1(new_n681), .B2(new_n679), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n651), .A2(KEYINPUT88), .A3(new_n679), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G330), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n610), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n609), .B1(new_n601), .B2(new_n606), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n297), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(new_n620), .A3(new_n597), .A4(new_n622), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n612), .B2(new_n676), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(new_n655), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n634), .B2(new_n676), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n686), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n565), .A2(new_n677), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n696), .A2(new_n692), .B1(new_n655), .B2(new_n676), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT89), .ZN(G399));
  INV_X1    g0499(.A(new_n212), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(new_n254), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n217), .B2(new_n702), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n659), .B1(new_n658), .B2(new_n660), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n521), .A2(KEYINPUT80), .A3(new_n524), .ZN(new_n709));
  AOI21_X1  g0509(.A(KEYINPUT80), .B1(new_n521), .B2(new_n524), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n660), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n708), .B1(new_n711), .B2(KEYINPUT26), .ZN(new_n712));
  OAI211_X1 g0512(.A(KEYINPUT29), .B(new_n676), .C1(new_n712), .C2(new_n657), .ZN(new_n713));
  INV_X1    g0513(.A(new_n584), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n517), .A2(new_n525), .A3(new_n529), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n660), .A2(new_n690), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n716), .B1(new_n565), .B2(new_n634), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n714), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  NOR4_X1   g0518(.A1(new_n498), .A2(new_n590), .A3(new_n516), .A4(KEYINPUT26), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n719), .B1(new_n711), .B2(KEYINPUT26), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n677), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n713), .B1(new_n721), .B2(KEYINPUT29), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n582), .A2(new_n513), .A3(new_n619), .A4(new_n613), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n505), .A2(new_n324), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n509), .A2(G257), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT90), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n557), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n635), .A2(KEYINPUT90), .A3(G179), .A4(new_n556), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n727), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(KEYINPUT91), .A2(KEYINPUT30), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n582), .B(KEYINPUT92), .ZN(new_n734));
  AOI21_X1  g0534(.A(G179), .B1(new_n614), .B2(new_n619), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n734), .A2(new_n735), .A3(new_n636), .A4(new_n526), .ZN(new_n736));
  INV_X1    g0536(.A(new_n732), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n727), .A2(new_n729), .A3(new_n730), .A4(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n733), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n740));
  AOI21_X1  g0540(.A(KEYINPUT31), .B1(new_n739), .B2(new_n677), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n681), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n655), .A2(new_n716), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n715), .A2(new_n743), .A3(new_n744), .A4(new_n676), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n685), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n722), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n706), .B1(new_n748), .B2(G1), .ZN(G364));
  NOR2_X1   g0549(.A1(new_n666), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n208), .B1(new_n750), .B2(G45), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n702), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT93), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n686), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n684), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G330), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT94), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n209), .A2(new_n374), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G200), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT97), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n306), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G326), .ZN(new_n769));
  AOI21_X1  g0569(.A(KEYINPUT98), .B1(new_n374), .B2(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n209), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n374), .A2(KEYINPUT98), .A3(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n306), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n768), .A2(new_n769), .B1(new_n775), .B2(new_n551), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G283), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n773), .A2(G190), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n766), .A2(G190), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  XOR2_X1   g0582(.A(KEYINPUT33), .B(G317), .Z(new_n783));
  OAI221_X1 g0583(.A(new_n777), .B1(new_n778), .B2(new_n780), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n763), .A2(G190), .A3(new_n304), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n785), .A2(KEYINPUT96), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(KEYINPUT96), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G322), .ZN(new_n790));
  INV_X1    g0590(.A(new_n763), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n791), .A2(G190), .A3(G200), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G311), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n352), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G179), .A2(G200), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n796), .A2(G20), .A3(new_n306), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n795), .B1(G329), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G294), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n209), .B1(new_n796), .B2(G190), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n790), .B(new_n799), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n472), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n352), .B(new_n803), .C1(new_n792), .C2(G77), .ZN(new_n804));
  INV_X1    g0604(.A(G159), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n797), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT32), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n804), .B(new_n807), .C1(new_n345), .C2(new_n788), .ZN(new_n808));
  INV_X1    g0608(.A(G50), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n768), .A2(new_n809), .B1(new_n780), .B2(new_n410), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n774), .A2(G87), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n811), .B(new_n812), .C1(new_n201), .C2(new_n782), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n784), .A2(new_n802), .B1(new_n808), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n215), .B1(G20), .B2(new_n369), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n815), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n761), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT95), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n700), .A2(new_n262), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(G45), .B2(new_n217), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n243), .B2(G45), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n700), .A2(new_n352), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(G355), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(G116), .B2(new_n212), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n820), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n816), .A2(new_n753), .A3(new_n827), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n755), .A2(new_n757), .B1(new_n762), .B2(new_n828), .ZN(G396));
  OAI221_X1 g0629(.A(new_n352), .B1(new_n797), .B2(new_n794), .C1(new_n793), .C2(new_n532), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n803), .B(new_n830), .C1(new_n789), .C2(G294), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n768), .A2(new_n551), .B1(new_n775), .B2(new_n410), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n779), .A2(G87), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n781), .A2(G283), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n831), .A2(new_n833), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT99), .Z(new_n837));
  AOI22_X1  g0637(.A1(new_n789), .A2(G143), .B1(G159), .B2(new_n792), .ZN(new_n838));
  INV_X1    g0638(.A(G137), .ZN(new_n839));
  INV_X1    g0639(.A(G150), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n838), .B1(new_n839), .B2(new_n768), .C1(new_n840), .C2(new_n782), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT34), .Z(new_n842));
  NAND2_X1  g0642(.A1(new_n779), .A2(G68), .ZN(new_n843));
  INV_X1    g0643(.A(G132), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n262), .B1(new_n797), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n801), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n845), .B1(G58), .B2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n843), .B(new_n847), .C1(new_n775), .C2(new_n809), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT100), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n842), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n815), .B1(new_n837), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n753), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n815), .A2(new_n758), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n852), .B1(new_n202), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n419), .A2(new_n677), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n424), .B1(new_n408), .B2(new_n676), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n855), .B1(new_n856), .B2(new_n419), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n851), .B(new_n854), .C1(new_n857), .C2(new_n759), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  OR2_X1    g0659(.A1(new_n721), .A2(new_n857), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n419), .A2(new_n424), .A3(new_n676), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n657), .B2(new_n663), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n860), .A2(new_n746), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT101), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n860), .A2(new_n863), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n753), .B1(new_n866), .B2(new_n747), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n859), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(G384));
  INV_X1    g0669(.A(new_n491), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n870), .A2(KEYINPUT35), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(KEYINPUT35), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n871), .A2(new_n872), .A3(G116), .A4(new_n216), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT36), .Z(new_n874));
  OAI211_X1 g0674(.A(new_n218), .B(G77), .C1(new_n345), .C2(new_n201), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n809), .A2(G68), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n208), .B(G13), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n677), .A2(new_n455), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n464), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n456), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n445), .B1(new_n466), .B2(new_n467), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n881), .B1(new_n882), .B2(new_n879), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n857), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n745), .B2(new_n742), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n351), .B1(new_n356), .B2(new_n201), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n383), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n377), .B1(new_n382), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n675), .ZN(new_n889));
  OAI22_X1  g0689(.A1(new_n340), .A2(new_n367), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n376), .A2(new_n888), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n390), .A2(new_n367), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n394), .A2(new_n387), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n367), .A2(new_n675), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n893), .A2(new_n894), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n888), .A2(new_n889), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n396), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT38), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n898), .A2(new_n900), .A3(KEYINPUT38), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT40), .B1(new_n885), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT40), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n897), .ZN(new_n910));
  INV_X1    g0710(.A(new_n895), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n396), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  XOR2_X1   g0713(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n907), .B1(new_n915), .B2(new_n904), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n906), .B1(new_n885), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n470), .B1(new_n745), .B2(new_n742), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n685), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n917), .B2(new_n918), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n861), .B1(new_n718), .B2(new_n720), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n905), .B(new_n883), .C1(new_n921), .C2(new_n855), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  INV_X1    g0723(.A(new_n904), .ZN(new_n924));
  INV_X1    g0724(.A(new_n914), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n910), .B2(new_n912), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n923), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n903), .A2(KEYINPUT39), .A3(new_n904), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n445), .A2(new_n455), .A3(new_n676), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n388), .A2(new_n392), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n889), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n922), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n713), .B(new_n469), .C1(new_n721), .C2(KEYINPUT29), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n646), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n934), .B(new_n936), .Z(new_n937));
  NAND2_X1  g0737(.A1(new_n920), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n208), .B2(new_n750), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n920), .A2(new_n937), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n878), .B1(new_n939), .B2(new_n940), .ZN(G367));
  OAI21_X1  g0741(.A(new_n715), .B1(new_n498), .B2(new_n676), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n658), .A2(new_n677), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(new_n692), .A3(new_n696), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT42), .Z(new_n946));
  INV_X1    g0746(.A(new_n944), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(new_n634), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n517), .A2(new_n525), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n676), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n676), .A2(new_n587), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(new_n584), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n660), .A2(new_n951), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n946), .A2(new_n950), .B1(KEYINPUT43), .B2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n954), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT43), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n695), .A2(new_n947), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n946), .A2(new_n957), .A3(new_n956), .A4(new_n950), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n960), .B1(new_n959), .B2(new_n961), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n701), .B(KEYINPUT41), .Z(new_n965));
  INV_X1    g0765(.A(KEYINPUT45), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n944), .A2(new_n697), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(KEYINPUT103), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n967), .A2(KEYINPUT103), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n970), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(KEYINPUT45), .A3(new_n968), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n944), .A2(new_n697), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT44), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n971), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n976), .A2(new_n686), .A3(new_n694), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n696), .A2(new_n692), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n694), .B2(new_n696), .ZN(new_n979));
  INV_X1    g0779(.A(new_n686), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n979), .B1(new_n980), .B2(KEYINPUT104), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT104), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n686), .B(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n981), .B1(new_n983), .B2(new_n979), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n748), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT105), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n971), .A2(new_n973), .A3(new_n975), .A4(new_n695), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n984), .A2(KEYINPUT105), .A3(new_n748), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n977), .A2(new_n987), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n965), .B1(new_n990), .B2(new_n748), .ZN(new_n991));
  INV_X1    g0791(.A(new_n751), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n964), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n821), .A2(new_n237), .B1(new_n700), .B2(new_n402), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n852), .B1(new_n820), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n775), .A2(new_n345), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n779), .A2(G77), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n782), .B2(new_n805), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n996), .B(new_n998), .C1(G143), .C2(new_n767), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n801), .A2(new_n201), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n262), .B1(new_n797), .B2(new_n839), .C1(new_n793), .C2(new_n809), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(new_n789), .C2(G150), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n779), .A2(G97), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n768), .B2(new_n794), .C1(new_n800), .C2(new_n782), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n801), .A2(new_n410), .ZN(new_n1007));
  INV_X1    g0807(.A(G317), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n352), .B1(new_n797), .B2(new_n1008), .C1(new_n793), .C2(new_n778), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1007), .B(new_n1009), .C1(new_n789), .C2(G303), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n775), .A2(new_n532), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1006), .B(new_n1010), .C1(KEYINPUT46), .C2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(KEYINPUT46), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT106), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1003), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT47), .Z(new_n1016));
  OAI221_X1 g0816(.A(new_n995), .B1(new_n761), .B2(new_n954), .C1(new_n1016), .C2(new_n817), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT107), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n993), .A2(new_n1018), .ZN(G387));
  INV_X1    g0819(.A(new_n703), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n824), .A2(new_n1020), .B1(new_n410), .B2(new_n700), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n234), .A2(new_n332), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n399), .A2(new_n809), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT50), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n703), .A2(new_n332), .A3(new_n239), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n821), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1021), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n852), .B1(new_n1027), .B2(new_n820), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n694), .B2(new_n761), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n801), .A2(new_n401), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n262), .B1(new_n797), .B2(new_n840), .C1(new_n793), .C2(new_n201), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1030), .B(new_n1031), .C1(new_n789), .C2(G50), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n805), .A2(new_n768), .B1(new_n782), .B2(new_n341), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n775), .A2(new_n202), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1032), .A2(new_n1034), .A3(new_n1004), .A4(new_n1036), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n788), .A2(new_n1008), .B1(new_n551), .B2(new_n793), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1038), .A2(KEYINPUT108), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(KEYINPUT108), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G311), .A2(new_n781), .B1(new_n767), .B2(G322), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT109), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT48), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n775), .A2(new_n800), .B1(new_n778), .B2(new_n801), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(KEYINPUT49), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n262), .B1(new_n798), .B2(G326), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(new_n532), .C2(new_n780), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1048), .A2(KEYINPUT49), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1037), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1029), .B1(new_n1053), .B2(new_n815), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT110), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n992), .B2(new_n984), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n984), .A2(new_n748), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n1057), .A2(KEYINPUT111), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(KEYINPUT111), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1058), .A2(new_n701), .A3(new_n985), .A4(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1056), .A2(new_n1060), .ZN(G393));
  AND2_X1   g0861(.A1(new_n977), .A2(new_n988), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n985), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n990), .B(new_n701), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n947), .A2(new_n760), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT112), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n768), .A2(new_n840), .B1(new_n788), .B2(new_n805), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT51), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n801), .A2(new_n202), .ZN(new_n1069));
  INV_X1    g0869(.A(G143), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n262), .B1(new_n797), .B2(new_n1070), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1069), .B(new_n1071), .C1(new_n399), .C2(new_n792), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n782), .A2(new_n809), .B1(new_n775), .B2(new_n201), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1068), .A2(new_n834), .A3(new_n1072), .A4(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n262), .B1(new_n798), .B2(G322), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1076), .B1(new_n532), .B2(new_n801), .C1(new_n793), .C2(new_n800), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n782), .A2(new_n551), .B1(new_n775), .B2(new_n778), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(G107), .C2(new_n779), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n768), .A2(new_n1008), .B1(new_n788), .B2(new_n794), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT52), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n817), .B1(new_n1075), .B2(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n821), .A2(new_n246), .B1(G97), .B2(new_n700), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n852), .B(new_n1083), .C1(new_n820), .C2(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1062), .A2(new_n992), .B1(new_n1066), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1064), .A2(new_n1086), .ZN(G390));
  INV_X1    g0887(.A(new_n741), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NOR3_X1   g0890(.A1(new_n639), .A2(new_n530), .A3(new_n677), .ZN(new_n1091));
  OAI211_X1 g0891(.A(G330), .B(new_n857), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n883), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n883), .B1(new_n921), .B2(new_n855), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1095), .A2(new_n929), .B1(new_n927), .B2(new_n928), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n929), .B1(new_n924), .B2(new_n926), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n856), .A2(new_n419), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n676), .B(new_n1098), .C1(new_n712), .C2(new_n657), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n855), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1097), .B1(new_n1101), .B2(new_n883), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1094), .B1(new_n1096), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1097), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n707), .B1(new_n662), .B2(new_n659), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n677), .B1(new_n718), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n855), .B1(new_n1106), .B2(new_n1098), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1104), .B1(new_n1107), .B2(new_n1093), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n927), .A2(new_n928), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1093), .B1(new_n863), .B2(new_n1100), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1109), .B1(new_n1110), .B2(new_n930), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n746), .A2(new_n857), .A3(new_n883), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1108), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1103), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n883), .B1(new_n746), .B2(new_n857), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1094), .A2(new_n1115), .B1(new_n921), .B2(new_n855), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1117), .A2(new_n1107), .A3(new_n1112), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n746), .A2(new_n469), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n935), .A2(new_n646), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1114), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1103), .A2(new_n1119), .A3(new_n1113), .A4(new_n1122), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1124), .A2(new_n701), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n759), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1109), .A2(new_n1127), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n352), .B1(new_n797), .B2(new_n800), .C1(new_n793), .C2(new_n472), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1069), .B(new_n1129), .C1(new_n789), .C2(G116), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(G107), .A2(new_n781), .B1(new_n767), .B2(G283), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1130), .A2(new_n812), .A3(new_n843), .A4(new_n1131), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n782), .A2(new_n839), .B1(new_n780), .B2(new_n809), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n801), .A2(new_n805), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n798), .A2(G125), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT54), .B(G143), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1136), .B(new_n262), .C1(new_n793), .C2(new_n1137), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1135), .B(new_n1138), .C1(new_n789), .C2(G132), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n774), .A2(G150), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1140), .B(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n767), .A2(G128), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1134), .A2(new_n1139), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n817), .B1(new_n1132), .B2(new_n1144), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n852), .B(new_n1145), .C1(new_n341), .C2(new_n853), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1128), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n1114), .B2(new_n751), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1126), .A2(new_n1149), .ZN(G378));
  INV_X1    g0950(.A(new_n934), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n905), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n857), .B(new_n883), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n907), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n685), .B1(new_n885), .B2(new_n916), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n300), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n645), .A2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n298), .A2(new_n889), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1160), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n313), .A2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1157), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n313), .A2(new_n1162), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1165), .A2(new_n1166), .A3(new_n1156), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1154), .A2(new_n1155), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1151), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1172));
  OAI21_X1  g0972(.A(KEYINPUT40), .B1(new_n924), .B2(new_n926), .ZN(new_n1173));
  OAI21_X1  g0973(.A(G330), .B1(new_n1153), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1172), .B1(new_n906), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1154), .A2(new_n1155), .A3(new_n1168), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1175), .A2(new_n1176), .A3(new_n934), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1171), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1172), .A2(new_n1127), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n853), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n753), .B1(G50), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1000), .B1(new_n767), .B2(G116), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT115), .Z(new_n1183));
  AOI211_X1 g0983(.A(new_n262), .B(new_n254), .C1(new_n798), .C2(G283), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n401), .B2(new_n793), .C1(new_n788), .C2(new_n410), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n782), .A2(new_n472), .B1(new_n780), .B2(new_n345), .ZN(new_n1186));
  NOR4_X1   g0986(.A1(new_n1183), .A2(new_n1035), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT116), .B(KEYINPUT58), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1187), .B(new_n1188), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(G33), .A2(G41), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT114), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1191), .B(new_n809), .C1(new_n262), .C2(new_n254), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n782), .A2(new_n844), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n792), .A2(G137), .B1(G150), .B2(new_n846), .ZN(new_n1194));
  INV_X1    g0994(.A(G128), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1194), .B1(new_n775), .B2(new_n1137), .C1(new_n788), .C2(new_n1195), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1193), .B(new_n1196), .C1(G125), .C2(new_n767), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1191), .B1(G124), .B2(new_n798), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT59), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1200), .B1(new_n805), .B2(new_n780), .C1(new_n1197), .C2(new_n1201), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1189), .B(new_n1192), .C1(new_n1199), .C2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1181), .B1(new_n1203), .B2(new_n815), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1178), .A2(new_n992), .B1(new_n1179), .B2(new_n1204), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1096), .A2(new_n1102), .A3(new_n1094), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1112), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1121), .B1(new_n1208), .B2(new_n1119), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1175), .A2(new_n1176), .A3(new_n934), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n934), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1211));
  OAI21_X1  g1011(.A(KEYINPUT57), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n701), .B1(new_n1209), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1125), .A2(new_n1122), .ZN(new_n1214));
  AOI21_X1  g1014(.A(KEYINPUT57), .B1(new_n1214), .B2(new_n1178), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1205), .B1(new_n1213), .B2(new_n1215), .ZN(G375));
  AND2_X1   g1016(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1093), .A2(new_n758), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n767), .A2(G294), .B1(G107), .B2(new_n792), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n532), .B2(new_n782), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT118), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n262), .B(new_n1030), .C1(G303), .C2(new_n798), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1223), .B(new_n997), .C1(new_n778), .C2(new_n788), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G97), .B2(new_n774), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n801), .A2(new_n809), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n262), .B1(new_n1195), .B2(new_n797), .C1(new_n793), .C2(new_n840), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1226), .B(new_n1227), .C1(new_n789), .C2(G137), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n844), .A2(new_n768), .B1(new_n782), .B2(new_n1137), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n345), .A2(new_n780), .B1(new_n775), .B2(new_n805), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1222), .A2(new_n1225), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n753), .B1(G68), .B2(new_n1180), .C1(new_n1232), .C2(new_n817), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1217), .A2(new_n751), .B1(new_n1219), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1217), .A2(new_n1121), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n965), .B(KEYINPUT117), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(new_n1123), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1235), .A2(new_n1238), .ZN(new_n1239));
  XOR2_X1   g1039(.A(new_n1239), .B(KEYINPUT119), .Z(G381));
  XOR2_X1   g1040(.A(G375), .B(KEYINPUT120), .Z(new_n1241));
  NOR2_X1   g1041(.A1(G393), .A2(G396), .ZN(new_n1242));
  INV_X1    g1042(.A(G390), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n702), .B1(new_n1114), .B2(new_n1123), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1148), .B1(new_n1125), .B2(new_n1244), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1242), .A2(new_n1243), .A3(new_n868), .A4(new_n1245), .ZN(new_n1246));
  OR4_X1    g1046(.A1(G387), .A2(new_n1241), .A3(G381), .A4(new_n1246), .ZN(G407));
  NOR2_X1   g1047(.A1(new_n673), .A2(G343), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1245), .A2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G407), .B(G213), .C1(new_n1241), .C2(new_n1249), .ZN(G409));
  AOI21_X1  g1050(.A(G390), .B1(new_n993), .B2(new_n1018), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(G396), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1242), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n993), .A2(new_n1018), .A3(G390), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1252), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1255), .B1(new_n1252), .B2(new_n1256), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(G378), .B(new_n1205), .C1(new_n1213), .C2(new_n1215), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1214), .A2(new_n1178), .A3(new_n1237), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1178), .A2(new_n992), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1179), .A2(new_n1204), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1245), .B1(new_n1261), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1260), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1217), .A2(KEYINPUT60), .A3(new_n1121), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1267), .A2(new_n701), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1123), .A2(KEYINPUT60), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1236), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(G384), .B1(new_n1271), .B2(new_n1235), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n868), .B(new_n1234), .C1(new_n1268), .C2(new_n1270), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1248), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1266), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT121), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT62), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1248), .B1(new_n1260), .B2(new_n1265), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1280), .A2(KEYINPUT121), .A3(new_n1274), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1278), .A2(new_n1279), .A3(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT122), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1278), .A2(KEYINPUT122), .A3(new_n1279), .A4(new_n1281), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1266), .A2(new_n1274), .A3(KEYINPUT62), .A4(new_n1275), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT123), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1280), .A2(KEYINPUT123), .A3(KEYINPUT62), .A4(new_n1274), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1284), .A2(new_n1285), .A3(new_n1291), .ZN(new_n1292));
  OR2_X1    g1092(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1248), .A2(G2897), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(new_n1293), .B(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1280), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT61), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1259), .B1(new_n1292), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT63), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1278), .A2(new_n1299), .A3(new_n1281), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1280), .A2(KEYINPUT63), .A3(new_n1274), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1297), .A2(new_n1259), .A3(new_n1300), .A4(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(KEYINPUT124), .B1(new_n1298), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT124), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1297), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1280), .A2(KEYINPUT121), .A3(new_n1274), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT121), .B1(new_n1280), .B2(new_n1274), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1307), .A2(new_n1308), .A3(KEYINPUT62), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1290), .B1(new_n1309), .B2(KEYINPUT122), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1306), .B1(new_n1310), .B2(new_n1284), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1305), .B(new_n1302), .C1(new_n1311), .C2(new_n1259), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1304), .A2(new_n1312), .ZN(G405));
  NAND2_X1  g1113(.A1(new_n1293), .A2(KEYINPUT125), .ZN(new_n1314));
  XOR2_X1   g1114(.A(new_n1314), .B(KEYINPUT126), .Z(new_n1315));
  XNOR2_X1  g1115(.A(new_n1315), .B(new_n1259), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(G375), .A2(new_n1245), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1260), .B(new_n1317), .C1(new_n1293), .C2(KEYINPUT125), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(new_n1316), .B(new_n1318), .ZN(G402));
endmodule


