//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1254, new_n1255,
    new_n1256, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n208), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT65), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n210), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n213), .B(new_n218), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G50), .B(G68), .Z(new_n236));
  XNOR2_X1  g0036(.A(G58), .B(G77), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G97), .B(G107), .Z(new_n239));
  XNOR2_X1  g0039(.A(G87), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  NAND3_X1  g0042(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(new_n216), .ZN(new_n244));
  NOR2_X1   g0044(.A1(KEYINPUT8), .A2(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT69), .B(G58), .ZN(new_n246));
  AOI21_X1  g0046(.A(new_n245), .B1(new_n246), .B2(KEYINPUT8), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n208), .A2(G33), .ZN(new_n249));
  INV_X1    g0049(.A(G150), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  OAI22_X1  g0052(.A1(new_n248), .A2(new_n249), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  AND2_X1   g0053(.A1(new_n253), .A2(KEYINPUT70), .ZN(new_n254));
  OAI21_X1  g0054(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(new_n253), .B2(KEYINPUT70), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n244), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G50), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n244), .B1(new_n207), .B2(G20), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n259), .B1(new_n260), .B2(G50), .ZN(new_n261));
  AOI21_X1  g0061(.A(KEYINPUT9), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT66), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT66), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G45), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n207), .A2(G274), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT67), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT67), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n269), .A2(new_n273), .A3(new_n270), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n275));
  AOI21_X1  g0075(.A(G1), .B1(new_n268), .B2(new_n264), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n272), .A2(new_n274), .B1(G226), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G222), .ZN(new_n282));
  INV_X1    g0082(.A(G77), .ZN(new_n283));
  OAI22_X1  g0083(.A1(new_n281), .A2(new_n282), .B1(new_n283), .B2(new_n279), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT68), .ZN(new_n285));
  AND2_X1   g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NOR2_X1   g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n285), .B1(new_n288), .B2(new_n280), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n279), .A2(KEYINPUT68), .A3(G1698), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n284), .B1(new_n291), .B2(G223), .ZN(new_n292));
  INV_X1    g0092(.A(G33), .ZN(new_n293));
  OAI211_X1 g0093(.A(G1), .B(G13), .C1(new_n293), .C2(new_n268), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n278), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n295), .A2(G200), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  AND2_X1   g0098(.A1(KEYINPUT77), .A2(KEYINPUT10), .ZN(new_n299));
  NOR3_X1   g0099(.A1(new_n296), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n257), .A2(KEYINPUT9), .A3(new_n261), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n263), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(KEYINPUT77), .A2(KEYINPUT10), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n303), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n263), .A2(new_n300), .A3(new_n305), .A4(new_n301), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n257), .A2(new_n261), .ZN(new_n308));
  AND2_X1   g0108(.A1(KEYINPUT71), .A2(G179), .ZN(new_n309));
  NOR2_X1   g0109(.A1(KEYINPUT71), .A2(G179), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  OR2_X1    g0112(.A1(new_n295), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n295), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n308), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G50), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n252), .A2(new_n317), .B1(new_n208), .B2(G68), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n249), .A2(new_n283), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n244), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT11), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n260), .ZN(new_n324));
  INV_X1    g0124(.A(G68), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT12), .ZN(new_n326));
  INV_X1    g0126(.A(new_n258), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n326), .B1(new_n327), .B2(new_n325), .ZN(new_n328));
  NOR3_X1   g0128(.A1(new_n258), .A2(KEYINPUT12), .A3(G68), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n324), .A2(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n320), .A2(new_n321), .ZN(new_n331));
  NOR3_X1   g0131(.A1(new_n323), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n272), .A2(new_n274), .B1(G238), .B2(new_n277), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n279), .A2(G232), .A3(G1698), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n279), .A2(G226), .A3(new_n280), .ZN(new_n336));
  INV_X1    g0136(.A(G97), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n335), .B(new_n336), .C1(new_n293), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n275), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT13), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n334), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n340), .B1(new_n334), .B2(new_n339), .ZN(new_n342));
  OAI21_X1  g0142(.A(G169), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n334), .A2(new_n339), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT13), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n334), .A2(new_n339), .A3(new_n340), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G179), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n343), .A2(KEYINPUT14), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT14), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n350), .B1(new_n347), .B2(G169), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n333), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n347), .A2(G200), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n345), .A2(G190), .A3(new_n346), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n353), .A2(new_n332), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT78), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n352), .A2(KEYINPUT78), .A3(new_n355), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n307), .A2(new_n316), .A3(new_n358), .A4(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n244), .ZN(new_n361));
  XNOR2_X1  g0161(.A(KEYINPUT15), .B(G87), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n362), .A2(new_n249), .ZN(new_n363));
  OR2_X1    g0163(.A1(KEYINPUT8), .A2(G58), .ZN(new_n364));
  NAND2_X1  g0164(.A1(KEYINPUT8), .A2(G58), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(KEYINPUT72), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT72), .ZN(new_n367));
  AND2_X1   g0167(.A1(KEYINPUT8), .A2(G58), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n367), .B1(new_n368), .B2(new_n245), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n366), .A2(new_n369), .A3(new_n251), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G20), .A2(G77), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n363), .B1(new_n372), .B2(KEYINPUT73), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT73), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n370), .A2(new_n374), .A3(new_n371), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n361), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  OR3_X1    g0176(.A1(new_n258), .A2(KEYINPUT74), .A3(G77), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT74), .B1(new_n258), .B2(G77), .ZN(new_n378));
  AOI22_X1  g0178(.A1(G77), .A2(new_n260), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT75), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT75), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n370), .A2(new_n374), .A3(new_n371), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n374), .B1(new_n370), .B2(new_n371), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n383), .A2(new_n384), .A3(new_n363), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n382), .B(new_n379), .C1(new_n385), .C2(new_n361), .ZN(new_n386));
  INV_X1    g0186(.A(G238), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n289), .B2(new_n290), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n279), .A2(G232), .A3(new_n280), .ZN(new_n389));
  INV_X1    g0189(.A(G107), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n389), .B1(new_n390), .B2(new_n279), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n275), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n272), .A2(new_n274), .B1(G244), .B2(new_n277), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G200), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n381), .A2(new_n386), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT76), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT76), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n381), .A2(new_n386), .A3(new_n395), .A4(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n392), .A2(G190), .A3(new_n393), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n397), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n247), .A2(new_n327), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(new_n324), .B2(new_n247), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT7), .B1(new_n288), .B2(new_n208), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT3), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n293), .ZN(new_n406));
  NAND2_X1  g0206(.A1(KEYINPUT3), .A2(G33), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n406), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(G68), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(G159), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n252), .A2(new_n411), .ZN(new_n412));
  AND2_X1   g0212(.A1(KEYINPUT69), .A2(G58), .ZN(new_n413));
  NOR2_X1   g0213(.A1(KEYINPUT69), .A2(G58), .ZN(new_n414));
  OAI21_X1  g0214(.A(G68), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n202), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n412), .B1(new_n416), .B2(G20), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n410), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT16), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n361), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n410), .A2(new_n417), .A3(KEYINPUT16), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n403), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n272), .A2(new_n274), .B1(G232), .B2(new_n277), .ZN(new_n423));
  OAI211_X1 g0223(.A(G223), .B(new_n280), .C1(new_n286), .C2(new_n287), .ZN(new_n424));
  OAI211_X1 g0224(.A(G226), .B(G1698), .C1(new_n286), .C2(new_n287), .ZN(new_n425));
  INV_X1    g0225(.A(G87), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n424), .B(new_n425), .C1(new_n293), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n275), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n423), .A2(new_n311), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n272), .A2(new_n274), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n277), .A2(G232), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n430), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n429), .B1(new_n432), .B2(G169), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT18), .B1(new_n422), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n412), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n201), .B1(new_n246), .B2(G68), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n435), .B1(new_n436), .B2(new_n208), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n406), .A2(new_n208), .A3(new_n407), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT7), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n325), .B1(new_n440), .B2(new_n408), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n419), .B1(new_n437), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n442), .A2(new_n244), .A3(new_n421), .ZN(new_n443));
  INV_X1    g0243(.A(new_n403), .ZN(new_n444));
  AND4_X1   g0244(.A1(new_n297), .A2(new_n430), .A3(new_n428), .A4(new_n431), .ZN(new_n445));
  AOI21_X1  g0245(.A(G200), .B1(new_n423), .B2(new_n428), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n443), .B(new_n444), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT17), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n423), .A2(new_n311), .A3(new_n428), .ZN(new_n450));
  AOI21_X1  g0250(.A(G169), .B1(new_n423), .B2(new_n428), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n443), .A2(new_n444), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT18), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n423), .A2(new_n297), .A3(new_n428), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(new_n432), .B2(G200), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n422), .A2(KEYINPUT17), .A3(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n434), .A2(new_n449), .A3(new_n455), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n381), .A2(new_n386), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n394), .A2(new_n312), .ZN(new_n461));
  AOI21_X1  g0261(.A(G169), .B1(new_n392), .B2(new_n393), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  OR3_X1    g0265(.A1(new_n401), .A2(new_n459), .A3(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n360), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT6), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n469), .A2(new_n337), .A3(G107), .ZN(new_n470));
  XNOR2_X1  g0270(.A(G97), .B(G107), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n470), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  OAI22_X1  g0272(.A1(new_n472), .A2(new_n208), .B1(new_n283), .B2(new_n252), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n390), .B1(new_n440), .B2(new_n408), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n244), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n258), .A2(G97), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n293), .A2(G1), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n327), .A2(new_n244), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n476), .B1(new_n478), .B2(G97), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT81), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n475), .A2(KEYINPUT81), .A3(new_n479), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g0284(.A(G244), .B(new_n280), .C1(new_n286), .C2(new_n287), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G250), .A2(G1698), .ZN(new_n490));
  NAND2_X1  g0290(.A1(KEYINPUT4), .A2(G244), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n490), .B1(new_n491), .B2(G1698), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n489), .B1(new_n279), .B2(new_n492), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n487), .A2(new_n493), .A3(KEYINPUT79), .ZN(new_n494));
  AOI21_X1  g0294(.A(KEYINPUT79), .B1(new_n487), .B2(new_n493), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n275), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n264), .A2(G1), .ZN(new_n497));
  XNOR2_X1  g0297(.A(KEYINPUT5), .B(G41), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n275), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G257), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(G274), .A3(new_n497), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n496), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n314), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n487), .A2(new_n493), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT79), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n487), .A2(new_n493), .A3(KEYINPUT79), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT80), .B1(new_n510), .B2(new_n275), .ZN(new_n511));
  OAI211_X1 g0311(.A(KEYINPUT80), .B(new_n275), .C1(new_n494), .C2(new_n495), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n503), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n484), .B(new_n505), .C1(new_n514), .C2(new_n312), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n502), .B1(new_n510), .B2(new_n275), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n480), .B1(new_n516), .B2(G190), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT80), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n496), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n502), .B1(new_n519), .B2(new_n512), .ZN(new_n520));
  INV_X1    g0320(.A(G200), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n270), .A2(G45), .ZN(new_n523));
  OAI21_X1  g0323(.A(G250), .B1(new_n264), .B2(G1), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n523), .B1(new_n275), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n279), .A2(G244), .A3(G1698), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n279), .A2(G238), .A3(new_n280), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G116), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n525), .B1(new_n529), .B2(new_n275), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT83), .B1(new_n530), .B2(G190), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n275), .ZN(new_n532));
  INV_X1    g0332(.A(new_n525), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n521), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n279), .A2(new_n208), .A3(G68), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT19), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n249), .B2(new_n337), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g0338(.A(KEYINPUT82), .B(G87), .ZN(new_n539));
  NOR2_X1   g0339(.A1(G97), .A2(G107), .ZN(new_n540));
  NAND3_X1  g0340(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n539), .A2(new_n540), .B1(new_n208), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n244), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n362), .A2(new_n327), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n478), .A2(G87), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n531), .A2(new_n534), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n530), .A2(KEYINPUT83), .A3(G190), .ZN(new_n548));
  AOI211_X1 g0348(.A(new_n312), .B(new_n525), .C1(new_n529), .C2(new_n275), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n532), .A2(new_n533), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n549), .B1(new_n314), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n362), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n478), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n543), .A2(new_n544), .A3(new_n553), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n547), .A2(new_n548), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n515), .A2(new_n522), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n499), .A2(G264), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n557), .A2(new_n501), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n279), .A2(G257), .A3(G1698), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n279), .A2(G250), .A3(new_n280), .ZN(new_n560));
  INV_X1    g0360(.A(G294), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n559), .B(new_n560), .C1(new_n293), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n275), .ZN(new_n563));
  AND3_X1   g0363(.A1(new_n558), .A2(new_n348), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(G169), .B1(new_n558), .B2(new_n563), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT86), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n208), .A2(KEYINPUT23), .A3(G107), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT23), .ZN(new_n569));
  OAI22_X1  g0369(.A1(new_n568), .A2(KEYINPUT85), .B1(new_n569), .B2(new_n390), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n390), .A3(G20), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT85), .ZN(new_n572));
  AOI21_X1  g0372(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n573));
  OAI22_X1  g0373(.A1(new_n571), .A2(new_n572), .B1(new_n573), .B2(G20), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n567), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n528), .A2(new_n569), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n568), .A2(KEYINPUT85), .B1(new_n576), .B2(new_n208), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n571), .A2(new_n572), .B1(KEYINPUT23), .B2(G107), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n577), .A2(KEYINPUT86), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n279), .A2(new_n208), .A3(G87), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT22), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT22), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n279), .A2(new_n583), .A3(new_n208), .A4(G87), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT24), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT24), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n580), .A2(new_n588), .A3(new_n585), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n361), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT25), .B1(new_n327), .B2(new_n390), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n327), .A2(KEYINPUT25), .A3(new_n390), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n592), .A2(new_n593), .B1(new_n478), .B2(G107), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n566), .B1(new_n590), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n558), .A2(new_n297), .A3(new_n563), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n563), .A2(new_n501), .A3(new_n557), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n597), .B1(new_n598), .B2(G200), .ZN(new_n599));
  INV_X1    g0399(.A(new_n589), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n588), .B1(new_n580), .B2(new_n585), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n244), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n602), .A3(new_n594), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n596), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(G264), .B(G1698), .C1(new_n286), .C2(new_n287), .ZN(new_n605));
  OAI211_X1 g0405(.A(G257), .B(new_n280), .C1(new_n286), .C2(new_n287), .ZN(new_n606));
  INV_X1    g0406(.A(G303), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n605), .B(new_n606), .C1(new_n607), .C2(new_n279), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n275), .ZN(new_n609));
  AND2_X1   g0409(.A1(KEYINPUT5), .A2(G41), .ZN(new_n610));
  NOR2_X1   g0410(.A1(KEYINPUT5), .A2(G41), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n497), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(G270), .A3(new_n294), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT84), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT84), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n612), .A2(new_n615), .A3(G270), .A4(new_n294), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n609), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(G190), .A3(new_n501), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n488), .B(new_n208), .C1(G33), .C2(new_n337), .ZN(new_n619));
  INV_X1    g0419(.A(G116), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G20), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n244), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT20), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n619), .A2(KEYINPUT20), .A3(new_n244), .A4(new_n621), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n258), .A2(G116), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n478), .B2(G116), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n609), .A2(new_n614), .A3(new_n501), .A4(new_n616), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n629), .B1(new_n630), .B2(G200), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n618), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n617), .A2(G179), .A3(new_n501), .A4(new_n629), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT21), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n314), .B1(new_n626), .B2(new_n628), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n634), .B1(new_n635), .B2(new_n630), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n635), .A2(new_n630), .A3(new_n634), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n632), .B(new_n633), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  NOR4_X1   g0438(.A1(new_n468), .A2(new_n556), .A3(new_n604), .A4(new_n638), .ZN(G372));
  INV_X1    g0439(.A(new_n316), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n343), .A2(KEYINPUT14), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n347), .A2(new_n350), .A3(G169), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n641), .B(new_n642), .C1(new_n348), .C2(new_n347), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n333), .A2(new_n643), .B1(new_n465), .B2(new_n355), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n449), .A2(new_n458), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n434), .B(new_n455), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n640), .B1(new_n646), .B2(new_n307), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n530), .A2(new_n311), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n648), .B(new_n554), .C1(G169), .C2(new_n530), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n534), .A2(new_n546), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n530), .A2(G190), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n652), .A2(new_n649), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n515), .A2(new_n522), .A3(new_n603), .A4(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n558), .A2(new_n348), .A3(new_n563), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n598), .B2(G169), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n602), .B2(new_n594), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n633), .B1(new_n637), .B2(new_n636), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT87), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT87), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n660), .B(new_n633), .C1(new_n637), .C2(new_n636), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n657), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n649), .B1(new_n654), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n505), .B1(new_n514), .B2(new_n312), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n652), .A2(new_n649), .A3(new_n480), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n520), .A2(new_n311), .B1(new_n314), .B2(new_n504), .ZN(new_n668));
  XOR2_X1   g0468(.A(KEYINPUT88), .B(KEYINPUT26), .Z(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n668), .A2(new_n555), .A3(new_n484), .A4(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n663), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n647), .B1(new_n468), .B2(new_n673), .ZN(G369));
  NAND3_X1  g0474(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AND4_X1   g0480(.A1(new_n629), .A2(new_n659), .A3(new_n661), .A4(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT89), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n638), .B1(new_n629), .B2(new_n680), .ZN(new_n683));
  OR3_X1    g0483(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n681), .A2(new_n682), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(G330), .A3(new_n685), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n596), .A2(new_n603), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n680), .B1(new_n590), .B2(new_n595), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n687), .A2(new_n688), .B1(new_n657), .B2(new_n680), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n680), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n658), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT90), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n596), .A2(new_n680), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n691), .A2(new_n697), .ZN(G399));
  NAND3_X1  g0498(.A1(new_n539), .A2(new_n620), .A3(new_n540), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT91), .Z(new_n700));
  INV_X1    g0500(.A(new_n211), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n700), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n214), .B2(new_n703), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n692), .B1(new_n663), .B2(new_n672), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(KEYINPUT93), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT93), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n709), .B(new_n692), .C1(new_n663), .C2(new_n672), .ZN(new_n710));
  XNOR2_X1  g0510(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n708), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n657), .A2(new_n658), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n654), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n547), .A2(new_n548), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n649), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n669), .B1(new_n515), .B2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n668), .A2(new_n653), .A3(KEYINPUT26), .A4(new_n480), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n717), .A2(new_n718), .B1(new_n554), .B2(new_n551), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n680), .B1(new_n714), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n712), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n550), .A2(new_n348), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n724), .A2(new_n598), .A3(new_n617), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n723), .B1(new_n725), .B2(new_n504), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n617), .A2(new_n563), .A3(new_n558), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n727), .A2(KEYINPUT30), .A3(new_n516), .A4(new_n724), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n630), .A2(new_n550), .A3(new_n311), .ZN(new_n730));
  INV_X1    g0530(.A(new_n598), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n514), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT92), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n730), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n514), .A2(KEYINPUT92), .A3(new_n731), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n729), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n680), .A2(KEYINPUT31), .ZN(new_n737));
  INV_X1    g0537(.A(new_n632), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n658), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n739), .A2(new_n596), .A3(new_n603), .A4(new_n692), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n736), .A2(new_n737), .B1(new_n556), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n733), .B1(new_n520), .B2(new_n598), .ZN(new_n742));
  INV_X1    g0542(.A(new_n730), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n735), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n726), .A2(new_n728), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(KEYINPUT31), .B1(new_n746), .B2(new_n680), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n741), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G330), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n722), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(KEYINPUT95), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT95), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n722), .A2(new_n754), .A3(new_n751), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n706), .B1(new_n756), .B2(G1), .ZN(G364));
  INV_X1    g0557(.A(G13), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n207), .B1(new_n759), .B2(G45), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OR3_X1    g0561(.A1(new_n702), .A2(KEYINPUT96), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(KEYINPUT96), .B1(new_n702), .B2(new_n761), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n216), .B1(G20), .B2(new_n314), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n211), .A2(new_n288), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT98), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n265), .A2(new_n267), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n773), .B1(new_n214), .B2(new_n774), .C1(new_n238), .C2(new_n264), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n701), .A2(new_n288), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n776), .A2(G355), .B1(new_n620), .B2(new_n701), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n777), .A2(KEYINPUT97), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(KEYINPUT97), .B2(new_n777), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n208), .A2(G190), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G179), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n411), .ZN(new_n784));
  XNOR2_X1  g0584(.A(KEYINPUT99), .B(KEYINPUT32), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n208), .A2(new_n521), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n312), .A2(G190), .A3(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n246), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n208), .A2(new_n297), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n312), .A2(new_n521), .A3(new_n790), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n786), .B1(new_n317), .B2(new_n788), .C1(new_n789), .C2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n781), .A2(new_n348), .A3(G200), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT100), .Z(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n312), .A2(new_n521), .A3(new_n781), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n795), .A2(new_n390), .B1(new_n283), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n312), .A2(new_n297), .A3(new_n787), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n325), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n208), .B1(new_n782), .B2(G190), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n790), .A2(new_n348), .A3(G200), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n279), .B1(new_n800), .B2(new_n337), .C1(new_n801), .C2(new_n539), .ZN(new_n802));
  NOR4_X1   g0602(.A1(new_n792), .A2(new_n797), .A3(new_n799), .A4(new_n802), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n803), .A2(KEYINPUT101), .ZN(new_n804));
  INV_X1    g0604(.A(G311), .ZN(new_n805));
  INV_X1    g0605(.A(G322), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n805), .A2(new_n796), .B1(new_n791), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n798), .ZN(new_n808));
  XNOR2_X1  g0608(.A(KEYINPUT33), .B(G317), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G329), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n288), .B1(new_n783), .B2(new_n811), .C1(new_n801), .C2(new_n607), .ZN(new_n812));
  INV_X1    g0612(.A(new_n800), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n812), .B1(G294), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n788), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n794), .A2(G283), .B1(G326), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n810), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n804), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(KEYINPUT101), .B2(new_n803), .ZN(new_n819));
  INV_X1    g0619(.A(new_n769), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n765), .B1(new_n771), .B2(new_n780), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n684), .A2(new_n685), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n821), .B1(new_n822), .B2(new_n768), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n686), .A2(new_n764), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n749), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G396));
  NAND2_X1  g0627(.A1(new_n465), .A2(new_n680), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT103), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n464), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n460), .A2(new_n680), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n460), .A2(new_n463), .A3(KEYINPUT103), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n828), .B1(new_n833), .B2(new_n401), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n708), .A2(new_n710), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n833), .A2(new_n401), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n837), .B(new_n692), .C1(new_n663), .C2(new_n672), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n765), .B1(new_n839), .B2(new_n751), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n751), .B2(new_n839), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n769), .A2(new_n766), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n764), .B1(new_n283), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n791), .ZN(new_n844));
  AOI22_X1  g0644(.A1(G137), .A2(new_n815), .B1(new_n844), .B2(G143), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n845), .B1(new_n250), .B2(new_n798), .C1(new_n411), .C2(new_n796), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT34), .ZN(new_n847));
  INV_X1    g0647(.A(G132), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n279), .B1(new_n783), .B2(new_n848), .C1(new_n801), .C2(new_n317), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n795), .A2(new_n325), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n849), .B(new_n850), .C1(new_n246), .C2(new_n813), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n288), .B1(new_n800), .B2(new_n337), .C1(new_n801), .C2(new_n390), .ZN(new_n852));
  INV_X1    g0652(.A(new_n796), .ZN(new_n853));
  AOI22_X1  g0653(.A1(G116), .A2(new_n853), .B1(new_n844), .B2(G294), .ZN(new_n854));
  INV_X1    g0654(.A(G283), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n854), .B1(new_n855), .B2(new_n798), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n852), .B(new_n856), .C1(G303), .C2(new_n815), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n794), .A2(G87), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n805), .B2(new_n783), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT102), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n847), .A2(new_n851), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n843), .B1(new_n820), .B2(new_n861), .C1(new_n834), .C2(new_n767), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n841), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(G384));
  INV_X1    g0664(.A(new_n472), .ZN(new_n865));
  OR2_X1    g0665(.A1(new_n865), .A2(KEYINPUT35), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(KEYINPUT35), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n866), .A2(G116), .A3(new_n217), .A4(new_n867), .ZN(new_n868));
  XNOR2_X1  g0668(.A(KEYINPUT104), .B(KEYINPUT36), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n868), .B(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n215), .A2(G77), .A3(new_n415), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n871), .A2(KEYINPUT105), .B1(G50), .B2(new_n325), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(KEYINPUT105), .B2(new_n871), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n758), .A2(G1), .ZN(new_n874));
  XOR2_X1   g0674(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n875));
  AND3_X1   g0675(.A1(new_n353), .A2(new_n332), .A3(new_n354), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n333), .B(new_n680), .C1(new_n643), .C2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n333), .A2(new_n680), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n352), .A2(new_n355), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n452), .A2(new_n453), .ZN(new_n881));
  INV_X1    g0681(.A(new_n678), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n453), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n881), .A2(new_n883), .A3(new_n447), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT37), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n881), .A2(new_n883), .A3(new_n886), .A4(new_n447), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n883), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n459), .A2(new_n889), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n888), .A2(new_n890), .A3(KEYINPUT38), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT38), .B1(new_n888), .B2(new_n890), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n834), .B(new_n880), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(KEYINPUT107), .B(new_n875), .C1(new_n893), .C2(new_n748), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n834), .A2(new_n880), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n888), .A2(new_n890), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n888), .A2(new_n890), .A3(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n746), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n604), .A2(new_n638), .A3(new_n680), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n515), .A2(new_n522), .A3(new_n555), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n692), .B1(new_n744), .B2(new_n745), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n901), .B(new_n904), .C1(KEYINPUT31), .C2(new_n905), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n895), .A2(new_n900), .A3(new_n906), .A4(KEYINPUT40), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n894), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n895), .A2(new_n900), .A3(new_n906), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT107), .B1(new_n909), .B2(new_n875), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n468), .A2(new_n748), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n749), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n912), .B2(new_n911), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n882), .B1(new_n434), .B2(new_n455), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n891), .B2(new_n892), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n898), .A2(KEYINPUT39), .A3(new_n899), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n643), .A2(new_n333), .A3(new_n692), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n915), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n880), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n680), .B1(new_n830), .B2(new_n832), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n924), .B1(new_n838), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n900), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n923), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n712), .A2(new_n467), .A3(new_n721), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n647), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n929), .B(new_n931), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n914), .A2(new_n932), .B1(new_n207), .B2(new_n759), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT108), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n914), .A2(new_n932), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n933), .B2(new_n934), .ZN(new_n937));
  OAI221_X1 g0737(.A(new_n870), .B1(new_n873), .B2(new_n874), .C1(new_n935), .C2(new_n937), .ZN(G367));
  NOR2_X1   g0738(.A1(new_n800), .A2(new_n325), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n844), .B2(G150), .ZN(new_n940));
  INV_X1    g0740(.A(G143), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n940), .B1(new_n941), .B2(new_n788), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT114), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n808), .A2(G159), .ZN(new_n946));
  INV_X1    g0746(.A(G137), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n279), .B1(new_n783), .B2(new_n947), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n789), .A2(new_n801), .B1(new_n793), .B2(new_n283), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n948), .B(new_n949), .C1(G50), .C2(new_n853), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n944), .A2(new_n945), .A3(new_n946), .A4(new_n950), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n607), .A2(new_n791), .B1(new_n788), .B2(new_n805), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT113), .Z(new_n953));
  INV_X1    g0753(.A(new_n801), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT46), .B1(new_n954), .B2(G116), .ZN(new_n955));
  INV_X1    g0755(.A(new_n793), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n279), .B1(new_n956), .B2(G97), .ZN(new_n957));
  INV_X1    g0757(.A(G317), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n957), .B1(new_n958), .B2(new_n783), .C1(new_n855), .C2(new_n796), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n954), .A2(KEYINPUT46), .A3(G116), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n390), .B2(new_n800), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n798), .A2(new_n561), .ZN(new_n962));
  OR4_X1    g0762(.A1(new_n955), .A2(new_n959), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n951), .B1(new_n953), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT47), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n769), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n546), .A2(new_n680), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n653), .A2(new_n967), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n968), .B(new_n768), .C1(new_n649), .C2(new_n967), .ZN(new_n969));
  INV_X1    g0769(.A(new_n773), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n770), .B1(new_n211), .B2(new_n362), .C1(new_n970), .C2(new_n234), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT112), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n971), .A2(new_n972), .ZN(new_n974));
  NOR3_X1   g0774(.A1(new_n973), .A2(new_n974), .A3(new_n764), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n966), .A2(new_n969), .A3(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n689), .ZN(new_n977));
  INV_X1    g0777(.A(new_n694), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n979), .A2(KEYINPUT111), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n686), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n980), .A2(new_n686), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n982), .A2(new_n983), .B1(new_n977), .B2(new_n978), .ZN(new_n984));
  INV_X1    g0784(.A(new_n983), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n977), .A2(new_n978), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n985), .A2(new_n986), .A3(new_n981), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n696), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n979), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n515), .A2(new_n522), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n480), .A2(new_n680), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n665), .A2(new_n480), .A3(new_n680), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n990), .A2(new_n991), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  OAI211_X1 g0799(.A(KEYINPUT110), .B(KEYINPUT44), .C1(new_n697), .C2(new_n996), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n979), .A2(new_n989), .A3(new_n996), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT45), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(KEYINPUT45), .B1(new_n697), .B2(new_n996), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n999), .B(new_n1000), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n690), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n697), .A2(KEYINPUT45), .A3(new_n996), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1009), .A2(new_n691), .A3(new_n999), .A4(new_n1000), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n756), .B1(new_n988), .B2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n702), .B(KEYINPUT41), .Z(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n761), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n695), .A2(new_n996), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT42), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n515), .B1(new_n997), .B2(new_n596), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n692), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT109), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n968), .B1(new_n649), .B2(new_n967), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT43), .Z(new_n1024));
  NAND3_X1  g0824(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1023), .A2(KEYINPUT43), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1018), .A2(new_n1020), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1022), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n1028), .A2(new_n1029), .B1(new_n691), .B2(new_n997), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1029), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n691), .A2(new_n997), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1031), .A2(new_n1032), .A3(new_n1027), .A4(new_n1025), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n976), .B1(new_n1015), .B2(new_n1034), .ZN(G387));
  NAND3_X1  g0835(.A1(new_n988), .A2(new_n755), .A3(new_n753), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n984), .A2(new_n987), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n756), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1036), .A2(new_n1038), .A3(new_n702), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n689), .A2(new_n768), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n231), .B1(new_n265), .B2(new_n267), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n776), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n1041), .A2(new_n970), .B1(new_n700), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n366), .A2(new_n369), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1044), .A2(G50), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT50), .ZN(new_n1046));
  AOI21_X1  g0846(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1046), .A2(new_n700), .A3(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1043), .A2(new_n1048), .B1(new_n390), .B2(new_n701), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n765), .B1(new_n1049), .B2(new_n771), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n794), .A2(G97), .B1(G50), .B2(new_n844), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n808), .A2(new_n247), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G68), .A2(new_n853), .B1(new_n815), .B2(G159), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n279), .B1(new_n783), .B2(new_n250), .C1(new_n801), .C2(new_n283), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n552), .B2(new_n813), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n783), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n279), .B1(new_n1057), .B2(G326), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n801), .A2(new_n561), .B1(new_n800), .B2(new_n855), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G317), .A2(new_n844), .B1(new_n815), .B2(G322), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n607), .B2(new_n796), .C1(new_n805), .C2(new_n798), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT48), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n1062), .B2(new_n1061), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT49), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1058), .B1(new_n620), .B2(new_n793), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1056), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1050), .B1(new_n1068), .B2(new_n769), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1037), .A2(new_n761), .B1(new_n1040), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1039), .A2(new_n1070), .ZN(G393));
  NAND2_X1  g0871(.A1(new_n1038), .A2(new_n1011), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1011), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1073), .A2(new_n756), .A3(new_n1037), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1072), .A2(new_n702), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n997), .A2(new_n768), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n770), .B1(new_n337), .B2(new_n211), .C1(new_n970), .C2(new_n241), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n765), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n858), .B1(new_n317), .B2(new_n798), .C1(new_n1044), .C2(new_n796), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n800), .A2(new_n283), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n279), .B1(new_n783), .B2(new_n941), .C1(new_n801), .C2(new_n325), .ZN(new_n1081));
  OR3_X1    g0881(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n250), .A2(new_n788), .B1(new_n791), .B2(new_n411), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT51), .Z(new_n1084));
  AOI22_X1  g0884(.A1(new_n808), .A2(G303), .B1(G116), .B2(new_n813), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n561), .B2(new_n796), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT115), .Z(new_n1087));
  OAI22_X1  g0887(.A1(new_n805), .A2(new_n791), .B1(new_n788), .B2(new_n958), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT52), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n288), .B1(new_n783), .B2(new_n806), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G283), .B2(new_n954), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1089), .B(new_n1091), .C1(new_n390), .C2(new_n795), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n1082), .A2(new_n1084), .B1(new_n1087), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1078), .B1(new_n1093), .B2(new_n769), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1073), .A2(new_n761), .B1(new_n1076), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1075), .A2(new_n1095), .ZN(G390));
  OAI21_X1  g0896(.A(new_n919), .B1(new_n927), .B2(new_n922), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n922), .B1(new_n898), .B2(new_n899), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n925), .B1(new_n720), .B2(new_n837), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1098), .B1(new_n1099), .B2(new_n924), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n906), .A2(G330), .A3(new_n834), .A4(new_n880), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1103), .A2(KEYINPUT116), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(KEYINPUT116), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1101), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1097), .A2(new_n1100), .A3(KEYINPUT116), .A4(new_n1103), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n920), .A2(new_n767), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n288), .B1(new_n783), .B2(new_n561), .C1(new_n801), .C2(new_n426), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1110), .A2(new_n1080), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n855), .B2(new_n788), .C1(new_n795), .C2(new_n325), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G97), .A2(new_n853), .B1(new_n808), .B2(G107), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n620), .B2(new_n791), .ZN(new_n1114));
  XOR2_X1   g0914(.A(KEYINPUT54), .B(G143), .Z(new_n1115));
  AOI22_X1  g0915(.A1(G128), .A2(new_n815), .B1(new_n853), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n848), .B2(new_n791), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n793), .A2(new_n317), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n288), .B(new_n1118), .C1(G125), .C2(new_n1057), .ZN(new_n1119));
  OAI21_X1  g0919(.A(KEYINPUT53), .B1(new_n801), .B2(new_n250), .ZN(new_n1120));
  NOR3_X1   g0920(.A1(new_n801), .A2(KEYINPUT53), .A3(new_n250), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(G159), .B2(new_n813), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n808), .A2(G137), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1119), .A2(new_n1120), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1112), .A2(new_n1114), .B1(new_n1117), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n769), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n842), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1126), .B(new_n765), .C1(new_n247), .C2(new_n1127), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n1108), .A2(new_n760), .B1(new_n1109), .B2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g0929(.A(G330), .B(new_n834), .C1(new_n741), .C2(new_n747), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n924), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1131), .A2(KEYINPUT117), .A3(new_n1102), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n838), .A2(new_n926), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT117), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1130), .A2(new_n1134), .A3(new_n924), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1132), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1131), .A2(new_n1099), .A3(new_n1102), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n467), .A2(new_n750), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n930), .A2(new_n647), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(KEYINPUT118), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT119), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT118), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1138), .A2(new_n1140), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1142), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n703), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1142), .A2(new_n1108), .A3(new_n1143), .A4(new_n1145), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1129), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(G378));
  INV_X1    g0951(.A(KEYINPUT57), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n304), .A2(new_n306), .A3(new_n316), .ZN(new_n1153));
  XOR2_X1   g0953(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1154));
  XNOR2_X1  g0954(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n308), .A2(new_n882), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT121), .Z(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1155), .B(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n911), .B2(G330), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n875), .B1(new_n893), .B2(new_n748), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT107), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1163), .A2(G330), .A3(new_n907), .A4(new_n894), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1155), .B(new_n1157), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n929), .B1(new_n1160), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n911), .A2(G330), .A3(new_n1159), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1168), .A2(new_n1169), .A3(new_n928), .A4(new_n923), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1152), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1108), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1140), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT123), .B1(new_n923), .B2(new_n928), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n1160), .B2(new_n1166), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1168), .A2(new_n1169), .A3(new_n1175), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1138), .A2(new_n1144), .A3(new_n1140), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1144), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1147), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1179), .B1(new_n1140), .B2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1174), .B(new_n702), .C1(new_n1183), .C2(KEYINPUT57), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1168), .A2(new_n1169), .A3(new_n1175), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1175), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n761), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n288), .A2(new_n268), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1189), .B(new_n317), .C1(G33), .C2(G41), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G97), .A2(new_n808), .B1(new_n815), .B2(G116), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n801), .A2(new_n283), .B1(new_n783), .B2(new_n855), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n789), .A2(new_n793), .ZN(new_n1193));
  NOR4_X1   g0993(.A1(new_n1192), .A2(new_n1193), .A3(new_n939), .A4(new_n1189), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n844), .A2(G107), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n853), .A2(new_n552), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1191), .A2(new_n1194), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1190), .B1(new_n1198), .B2(KEYINPUT58), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT120), .Z(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(KEYINPUT58), .ZN(new_n1201));
  INV_X1    g1001(.A(G128), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n1202), .A2(new_n791), .B1(new_n796), .B2(new_n947), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n954), .A2(new_n1115), .B1(new_n813), .B2(G150), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n848), .B2(new_n798), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1203), .B(new_n1205), .C1(G125), .C2(new_n815), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1207), .A2(KEYINPUT59), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(KEYINPUT59), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n956), .A2(G159), .ZN(new_n1210));
  AOI211_X1 g1010(.A(G33), .B(G41), .C1(new_n1057), .C2(G124), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1200), .B(new_n1201), .C1(new_n1208), .C2(new_n1212), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1213), .A2(new_n769), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n765), .B1(G50), .B2(new_n1127), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(new_n1165), .C2(new_n766), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT122), .Z(new_n1217));
  NAND2_X1  g1017(.A1(new_n1188), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1184), .A2(new_n1219), .ZN(G375));
  NAND2_X1  g1020(.A1(new_n1138), .A2(new_n761), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n765), .B1(G68), .B2(new_n1127), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n853), .A2(G150), .B1(new_n808), .B2(new_n1115), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(G132), .A2(new_n815), .B1(new_n844), .B2(G137), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n801), .A2(new_n411), .B1(new_n783), .B2(new_n1202), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n800), .A2(new_n317), .ZN(new_n1226));
  NOR4_X1   g1026(.A1(new_n1225), .A2(new_n1193), .A3(new_n288), .A4(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1223), .A2(new_n1224), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n279), .B1(new_n794), .B2(G77), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT124), .Z(new_n1230));
  AOI22_X1  g1030(.A1(new_n954), .A2(G97), .B1(new_n1057), .B2(G303), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n362), .B2(new_n800), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G283), .B2(new_n844), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(G107), .A2(new_n853), .B1(new_n808), .B2(G116), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1233), .B(new_n1234), .C1(new_n561), .C2(new_n788), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1228), .B1(new_n1230), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1222), .B1(new_n1236), .B2(new_n769), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n880), .B2(new_n767), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1221), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  OR2_X1    g1040(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1142), .A2(new_n1145), .A3(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1240), .B1(new_n1242), .B2(new_n1013), .ZN(G381));
  OAI21_X1  g1043(.A(new_n1187), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1152), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1182), .A2(new_n1140), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n703), .B1(new_n1246), .B2(new_n1171), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1218), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1150), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1039), .A2(new_n826), .A3(new_n1070), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1251), .A2(new_n863), .A3(new_n1075), .A4(new_n1095), .ZN(new_n1252));
  OR4_X1    g1052(.A1(G387), .A2(new_n1249), .A3(G381), .A4(new_n1252), .ZN(G407));
  NAND2_X1  g1053(.A1(new_n679), .A2(G213), .ZN(new_n1254));
  XOR2_X1   g1054(.A(new_n1254), .B(KEYINPUT125), .Z(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  OAI211_X1 g1056(.A(G407), .B(G213), .C1(new_n1249), .C2(new_n1256), .ZN(G409));
  NAND2_X1  g1057(.A1(new_n1255), .A2(G2897), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n702), .B1(new_n1260), .B2(KEYINPUT60), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1180), .A2(new_n1181), .A3(new_n1260), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT60), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1262), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT126), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1261), .B1(new_n1242), .B2(KEYINPUT60), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(KEYINPUT126), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(G384), .B1(new_n1270), .B2(new_n1240), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n863), .B(new_n1239), .C1(new_n1267), .C2(new_n1269), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1259), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1268), .A2(KEYINPUT126), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n1266), .B(new_n1261), .C1(new_n1242), .C2(KEYINPUT60), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1240), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n863), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1270), .A2(G384), .A3(new_n1240), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1277), .A2(new_n1278), .A3(new_n1258), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1280), .A2(new_n702), .A3(new_n1149), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1187), .B(new_n1014), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1129), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1216), .B1(new_n1284), .B2(new_n761), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .A4(new_n1285), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1256), .B(new_n1286), .C1(new_n1248), .C2(new_n1150), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1273), .A2(new_n1279), .A3(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1290));
  OAI21_X1  g1090(.A(KEYINPUT62), .B1(new_n1290), .B2(new_n1287), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1150), .B1(new_n1184), .B2(new_n1219), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1286), .A2(new_n1256), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT62), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1294), .A2(new_n1295), .A3(new_n1277), .A4(new_n1278), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1288), .A2(new_n1289), .A3(new_n1291), .A4(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n976), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n760), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1034), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1298), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n826), .B1(new_n1039), .B2(new_n1070), .ZN(new_n1303));
  OAI22_X1  g1103(.A1(new_n1302), .A2(KEYINPUT127), .B1(new_n1251), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1303), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1305), .A2(G387), .A3(new_n1250), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1304), .A2(G390), .A3(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(G390), .B1(new_n1304), .B2(new_n1306), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1297), .A2(new_n1309), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1290), .A2(new_n1287), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1309), .B1(new_n1311), .B2(KEYINPUT63), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT63), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1313), .B1(new_n1290), .B2(new_n1287), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1312), .A2(new_n1289), .A3(new_n1288), .A4(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1310), .A2(new_n1315), .ZN(G405));
  NAND2_X1  g1116(.A1(G375), .A2(G378), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1249), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1318), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1290), .A2(new_n1249), .A3(new_n1317), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1309), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1321), .B(new_n1322), .ZN(G402));
endmodule


