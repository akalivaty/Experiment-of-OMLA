//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1195, new_n1196, new_n1197, new_n1199, new_n1200, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT65), .ZN(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  AND2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(G58), .ZN(new_n209));
  INV_X1    g0009(.A(G232), .ZN(new_n210));
  INV_X1    g0010(.A(G116), .ZN(new_n211));
  INV_X1    g0011(.A(G270), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G87), .B2(G250), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G97), .A2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G68), .A2(G238), .ZN(new_n220));
  XOR2_X1   g0020(.A(KEYINPUT66), .B(G77), .Z(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G244), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n214), .A2(new_n219), .A3(new_n220), .A4(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT1), .Z(new_n226));
  NOR2_X1   g0026(.A1(new_n224), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT0), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n203), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G50), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n226), .B(new_n229), .C1(new_n233), .C2(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n210), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT2), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n217), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT67), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G264), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n212), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n241), .B(new_n245), .Z(G358));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G107), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n211), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G68), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(new_n216), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(new_n209), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT72), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n255), .A2(KEYINPUT72), .A3(G13), .A4(G20), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G50), .ZN(new_n261));
  NAND3_X1  g0061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n230), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n260), .B(new_n264), .C1(G1), .C2(new_n231), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n216), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G150), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(G20), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT8), .B(G58), .ZN(new_n272));
  OAI221_X1 g0072(.A(new_n268), .B1(new_n271), .B2(new_n272), .C1(new_n205), .C2(new_n231), .ZN(new_n273));
  AOI211_X1 g0073(.A(new_n261), .B(new_n266), .C1(new_n273), .C2(new_n263), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n278), .B1(G222), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G223), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n280), .B1(new_n281), .B2(new_n279), .ZN(new_n282));
  AND2_X1   g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(new_n230), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT3), .B(G33), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n282), .B(new_n284), .C1(new_n221), .C2(new_n285), .ZN(new_n286));
  OR2_X1    g0086(.A1(KEYINPUT69), .A2(G41), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT69), .A2(G41), .ZN(new_n288));
  AOI21_X1  g0088(.A(G45), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(KEYINPUT70), .B1(new_n289), .B2(G1), .ZN(new_n290));
  INV_X1    g0090(.A(G274), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT71), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(new_n283), .B2(new_n230), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G41), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n294), .A2(KEYINPUT71), .A3(G1), .A4(G13), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n291), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G45), .ZN(new_n297));
  INV_X1    g0097(.A(new_n288), .ZN(new_n298));
  NOR2_X1   g0098(.A1(KEYINPUT69), .A2(G41), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT70), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n300), .A2(new_n301), .A3(new_n255), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n290), .A2(new_n296), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n293), .A2(new_n295), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n255), .B1(G41), .B2(G45), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n286), .B(new_n303), .C1(new_n217), .C2(new_n306), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n274), .A2(KEYINPUT9), .B1(G200), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n261), .B1(new_n273), .B2(new_n263), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(new_n216), .B2(new_n265), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT9), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n308), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT10), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT10), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n308), .A2(new_n312), .A3(new_n317), .A4(new_n314), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n307), .A2(new_n320), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n307), .A2(G179), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n310), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT77), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT17), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n304), .A2(G232), .A3(new_n305), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n275), .A2(new_n277), .A3(G223), .A4(new_n279), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n275), .A2(new_n277), .A3(G226), .A4(G1698), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G33), .A2(G87), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n284), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n303), .A2(new_n328), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G200), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n303), .A2(new_n333), .A3(new_n313), .A4(new_n328), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n260), .ZN(new_n340));
  INV_X1    g0140(.A(new_n272), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(new_n265), .B2(new_n341), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT7), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n285), .B2(G20), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n276), .A2(G33), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n348));
  OAI211_X1 g0148(.A(KEYINPUT7), .B(new_n231), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G68), .ZN(new_n351));
  INV_X1    g0151(.A(G68), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n209), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(G20), .B1(new_n353), .B2(new_n203), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n267), .A2(G159), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n351), .A2(KEYINPUT16), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n263), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n346), .A2(KEYINPUT76), .A3(new_n349), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT76), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n278), .A2(new_n361), .A3(KEYINPUT7), .A4(new_n231), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(G68), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT16), .B1(new_n363), .B2(new_n357), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n344), .B1(new_n359), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n327), .B1(new_n339), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(KEYINPUT77), .A2(KEYINPUT17), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n363), .A2(new_n357), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT16), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n356), .B1(new_n350), .B2(G68), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n264), .B1(new_n371), .B2(KEYINPUT16), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n343), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n367), .B1(new_n373), .B2(new_n338), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n366), .B1(new_n374), .B2(new_n327), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n334), .A2(G169), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n303), .A2(new_n333), .A3(G179), .A4(new_n328), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n365), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT18), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n365), .A2(KEYINPUT18), .A3(new_n379), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n376), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G238), .A2(G1698), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n285), .B(new_n387), .C1(new_n210), .C2(G1698), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n388), .B(new_n284), .C1(G107), .C2(new_n285), .ZN(new_n389));
  INV_X1    g0189(.A(G244), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n303), .B(new_n389), .C1(new_n390), .C2(new_n306), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n320), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n341), .A2(new_n267), .B1(new_n221), .B2(G20), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT15), .B(G87), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n393), .B1(new_n271), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n265), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n395), .A2(new_n263), .B1(new_n396), .B2(G77), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT73), .ZN(new_n398));
  INV_X1    g0198(.A(new_n221), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n340), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n397), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n398), .B1(new_n397), .B2(new_n400), .ZN(new_n403));
  OAI221_X1 g0203(.A(new_n392), .B1(G179), .B2(new_n391), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n397), .A2(new_n400), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT73), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n391), .A2(G200), .ZN(new_n407));
  OR2_X1    g0207(.A1(new_n391), .A2(new_n313), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n401), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n386), .B1(KEYINPUT74), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n324), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(KEYINPUT74), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G33), .A2(G97), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n210), .A2(G1698), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(G226), .B2(G1698), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n414), .B1(new_n416), .B2(new_n278), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n284), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n304), .A2(G238), .A3(new_n305), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n303), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT13), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT75), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT13), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n303), .A2(new_n418), .A3(new_n423), .A4(new_n419), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n303), .A2(new_n419), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n426), .A2(KEYINPUT75), .A3(new_n423), .A4(new_n418), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(G200), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n340), .A2(new_n352), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT12), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n270), .A2(G77), .B1(new_n267), .B2(G50), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n231), .B2(G68), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n432), .A2(new_n263), .ZN(new_n433));
  OR2_X1    g0233(.A1(new_n433), .A2(KEYINPUT11), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n396), .A2(G68), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(KEYINPUT11), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n430), .A2(new_n434), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n421), .A2(G190), .A3(new_n424), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n428), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n425), .A2(G169), .A3(new_n427), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT14), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n421), .A2(G179), .A3(new_n424), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT14), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n425), .A2(new_n445), .A3(G169), .A4(new_n427), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n443), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n441), .B1(new_n447), .B2(new_n437), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n413), .A2(new_n448), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n412), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n360), .A2(G107), .A3(new_n362), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n267), .A2(G77), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n453), .A2(KEYINPUT78), .ZN(new_n454));
  INV_X1    g0254(.A(G107), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(KEYINPUT6), .A3(G97), .ZN(new_n456));
  XOR2_X1   g0256(.A(G97), .B(G107), .Z(new_n457));
  OAI21_X1  g0257(.A(new_n456), .B1(new_n457), .B2(KEYINPUT6), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n458), .A2(G20), .B1(KEYINPUT78), .B2(new_n453), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n452), .A2(new_n454), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n263), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n260), .A2(G97), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n255), .A2(G33), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n260), .A2(new_n264), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G97), .ZN(new_n466));
  OR2_X1    g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n461), .A2(new_n463), .A3(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n275), .A2(new_n277), .A3(G244), .A4(new_n279), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT4), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n470), .A2(new_n390), .A3(G1698), .ZN(new_n472));
  AND2_X1   g0272(.A1(G250), .A2(G1698), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n285), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n471), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT5), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n287), .A2(new_n477), .A3(new_n288), .ZN(new_n478));
  OR2_X1    g0278(.A1(new_n477), .A2(G41), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n297), .A2(G1), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n476), .A2(new_n284), .B1(new_n482), .B2(new_n296), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n481), .A2(G257), .A3(new_n304), .ZN(new_n484));
  AOI21_X1  g0284(.A(G169), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G179), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n476), .A2(new_n284), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n482), .A2(new_n296), .ZN(new_n489));
  AND4_X1   g0289(.A1(new_n487), .A2(new_n488), .A3(new_n489), .A4(new_n484), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n468), .A2(new_n486), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n483), .A2(new_n484), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G190), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n462), .B1(new_n460), .B2(new_n263), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(G200), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n467), .A4(new_n497), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n275), .A2(new_n277), .A3(new_n231), .A4(G87), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT22), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT22), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n285), .A2(new_n502), .A3(new_n231), .A4(G87), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n270), .A2(G116), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n231), .A2(G107), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n506), .B(KEYINPUT23), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT24), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n504), .A2(KEYINPUT24), .A3(new_n505), .A4(new_n507), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n263), .A3(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT25), .B1(new_n260), .B2(G107), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n260), .A2(new_n264), .A3(G107), .A4(new_n464), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT25), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n258), .A2(new_n515), .A3(new_n455), .A4(new_n259), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n513), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT83), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT83), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n513), .A2(new_n514), .A3(new_n519), .A4(new_n516), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n512), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n285), .A2(G257), .A3(G1698), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n285), .A2(G250), .A3(new_n279), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G294), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n284), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n481), .A2(G264), .A3(new_n304), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(new_n489), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n335), .ZN(new_n530));
  OR2_X1    g0330(.A1(new_n530), .A2(KEYINPUT84), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n530), .B(KEYINPUT84), .C1(G190), .C2(new_n529), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n522), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n512), .A2(new_n521), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n529), .A2(new_n320), .ZN(new_n535));
  OR2_X1    g0335(.A1(new_n529), .A2(G179), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n499), .A2(new_n533), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n465), .A2(new_n211), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n262), .A2(new_n230), .B1(G20), .B2(new_n211), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n475), .B(new_n231), .C1(G33), .C2(new_n466), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n541), .A2(KEYINPUT20), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT20), .B1(new_n541), .B2(new_n542), .ZN(new_n544));
  OR2_X1    g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n340), .A2(new_n211), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n540), .A2(KEYINPUT81), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT81), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n546), .B1(new_n543), .B2(new_n544), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n548), .B1(new_n549), .B2(new_n539), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n275), .A2(new_n277), .A3(G257), .A4(new_n279), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT80), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT80), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n285), .A2(new_n554), .A3(G257), .A4(new_n279), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n278), .A2(G303), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n285), .A2(G264), .A3(G1698), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n553), .A2(new_n555), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n558), .A2(new_n284), .B1(new_n296), .B2(new_n482), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n481), .A2(G270), .A3(new_n304), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n320), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT21), .B1(new_n551), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT82), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n558), .A2(new_n284), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n564), .A2(new_n489), .A3(new_n560), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n561), .A2(KEYINPUT21), .B1(new_n565), .B2(G179), .ZN(new_n566));
  INV_X1    g0366(.A(new_n551), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n563), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT21), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n565), .A2(new_n569), .A3(new_n320), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n564), .A2(new_n489), .A3(new_n560), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n571), .A2(new_n487), .ZN(new_n572));
  OAI211_X1 g0372(.A(KEYINPUT82), .B(new_n551), .C1(new_n570), .C2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n562), .B1(new_n568), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n571), .A2(G200), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n567), .B(new_n575), .C1(new_n313), .C2(new_n571), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n275), .A2(new_n277), .A3(G244), .A4(G1698), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n275), .A2(new_n277), .A3(G238), .A4(new_n279), .ZN(new_n578));
  NAND2_X1  g0378(.A1(G33), .A2(G116), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n284), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n480), .A2(new_n292), .A3(G274), .ZN(new_n582));
  INV_X1    g0382(.A(new_n480), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n304), .A2(G250), .A3(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n581), .A2(G190), .A3(new_n582), .A4(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n586), .B1(G200), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT19), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n231), .B1(new_n414), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(G87), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n591), .A2(new_n466), .A3(new_n455), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n275), .A2(new_n277), .A3(new_n231), .A4(G68), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n589), .B1(new_n414), .B2(G20), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n263), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n340), .A2(new_n394), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n260), .A2(new_n264), .A3(G87), .A4(new_n464), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n587), .A2(new_n320), .ZN(new_n601));
  XNOR2_X1  g0401(.A(new_n394), .B(KEYINPUT79), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n597), .B(new_n598), .C1(new_n465), .C2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n581), .A2(new_n487), .A3(new_n582), .A4(new_n584), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n588), .A2(new_n600), .B1(new_n601), .B2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n538), .A2(new_n574), .A3(new_n576), .A4(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n451), .A2(new_n607), .ZN(G372));
  NAND3_X1  g0408(.A1(new_n584), .A2(KEYINPUT86), .A3(new_n582), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT86), .B1(new_n584), .B2(new_n582), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT85), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n580), .A2(new_n612), .A3(new_n284), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n612), .B1(new_n580), .B2(new_n284), .ZN(new_n615));
  OAI22_X1  g0415(.A1(new_n610), .A2(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n586), .B1(new_n616), .B2(G200), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT87), .ZN(new_n618));
  XNOR2_X1  g0418(.A(new_n600), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n616), .A2(new_n320), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n617), .A2(new_n619), .B1(new_n620), .B2(new_n605), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n621), .A2(new_n533), .A3(new_n492), .A4(new_n498), .ZN(new_n622));
  INV_X1    g0422(.A(new_n562), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n551), .B1(new_n570), .B2(new_n572), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n622), .B1(new_n537), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n584), .A2(new_n582), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT86), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n581), .A2(KEYINPUT85), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n629), .A2(new_n609), .B1(new_n630), .B2(new_n613), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n605), .B1(new_n631), .B2(G169), .ZN(new_n632));
  AOI211_X1 g0432(.A(new_n485), .B(new_n490), .C1(new_n496), .C2(new_n467), .ZN(new_n633));
  XNOR2_X1  g0433(.A(KEYINPUT88), .B(KEYINPUT26), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n633), .A2(new_n606), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT26), .B1(new_n621), .B2(new_n633), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n626), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n450), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n323), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n447), .A2(new_n437), .ZN(new_n641));
  AOI211_X1 g0441(.A(new_n441), .B(new_n376), .C1(new_n641), .C2(new_n404), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(new_n385), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n640), .B1(new_n643), .B2(new_n319), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n639), .A2(new_n644), .ZN(G369));
  INV_X1    g0445(.A(G13), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n646), .A2(G1), .A3(G20), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT27), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g0449(.A(new_n649), .B(KEYINPUT89), .Z(new_n650));
  OR2_X1    g0450(.A1(new_n647), .A2(new_n648), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(G213), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G343), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OR3_X1    g0455(.A1(new_n625), .A2(new_n567), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n574), .A2(new_n576), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n567), .A2(new_n655), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G330), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n537), .A2(new_n654), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n533), .B1(new_n522), .B2(new_n655), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n662), .B1(new_n663), .B2(new_n537), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n574), .A2(new_n654), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n664), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(new_n662), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n665), .A2(new_n669), .ZN(G399));
  NAND2_X1  g0470(.A1(new_n287), .A2(new_n288), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n227), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n592), .A2(G116), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G1), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n235), .B2(new_n675), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT28), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n572), .A2(KEYINPUT90), .ZN(new_n680));
  INV_X1    g0480(.A(new_n587), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT90), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n571), .B2(new_n487), .ZN(new_n683));
  OAI211_X1 g0483(.A(new_n527), .B(new_n528), .C1(KEYINPUT91), .C2(KEYINPUT30), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n493), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n680), .A2(new_n681), .A3(new_n683), .A4(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(KEYINPUT91), .A2(KEYINPUT30), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n494), .A2(new_n631), .A3(G179), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n690), .A2(new_n529), .A3(new_n571), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n654), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT31), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n692), .A2(KEYINPUT31), .A3(new_n654), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT92), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n695), .A2(KEYINPUT92), .A3(new_n696), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n699), .B(new_n700), .C1(new_n607), .C2(new_n654), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G330), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n622), .B1(new_n574), .B2(new_n537), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n585), .B1(new_n631), .B2(new_n335), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n600), .B(KEYINPUT87), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n632), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT26), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n706), .A2(new_n492), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n634), .B1(new_n633), .B2(new_n606), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n632), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n703), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n711), .A2(new_n712), .A3(new_n654), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n713), .A2(KEYINPUT93), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n638), .A2(new_n655), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n712), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n713), .A2(KEYINPUT93), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n702), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n679), .B1(new_n720), .B2(G1), .ZN(G364));
  NOR2_X1   g0521(.A1(new_n646), .A2(G20), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n255), .B1(new_n722), .B2(G45), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n675), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n724), .B(KEYINPUT94), .Z(new_n725));
  NOR2_X1   g0525(.A1(new_n661), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(G330), .B2(new_n659), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n253), .A2(G45), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n673), .A2(new_n285), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n728), .B(new_n729), .C1(G45), .C2(new_n235), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n285), .A2(G355), .A3(new_n227), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n730), .B(new_n731), .C1(G116), .C2(new_n227), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT95), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G13), .A2(G33), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n230), .B1(G20), .B2(new_n320), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n734), .A2(new_n735), .A3(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n725), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n231), .A2(new_n487), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(new_n313), .A3(G200), .ZN(new_n744));
  INV_X1    g0544(.A(G317), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n744), .B1(KEYINPUT33), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(KEYINPUT33), .B2(new_n745), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n743), .A2(G190), .A3(G200), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n285), .B1(new_n749), .B2(G326), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n487), .A2(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n231), .A2(G190), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n751), .B1(G311), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n231), .A2(new_n313), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n752), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G322), .ZN(new_n760));
  OR3_X1    g0560(.A1(KEYINPUT96), .A2(G179), .A3(G200), .ZN(new_n761));
  OAI21_X1  g0561(.A(KEYINPUT96), .B1(G179), .B2(G200), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n313), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n231), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G294), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n335), .A2(G179), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n757), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G303), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n753), .A2(new_n767), .ZN(new_n770));
  INV_X1    g0570(.A(G283), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n768), .A2(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n231), .B(G190), .C1(new_n761), .C2(new_n762), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n772), .B1(G329), .B2(new_n773), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n756), .A2(new_n760), .A3(new_n766), .A4(new_n774), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n285), .B1(new_n744), .B2(new_n352), .C1(new_n216), .C2(new_n748), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n399), .A2(new_n754), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n768), .A2(new_n591), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n770), .A2(new_n455), .ZN(new_n779));
  NOR4_X1   g0579(.A1(new_n776), .A2(new_n777), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n780), .B1(new_n209), .B2(new_n758), .C1(new_n466), .C2(new_n764), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n773), .A2(G159), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT32), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n775), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n742), .B1(new_n784), .B2(new_n739), .ZN(new_n785));
  INV_X1    g0585(.A(new_n738), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n741), .B(new_n785), .C1(new_n659), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n727), .A2(new_n787), .ZN(G396));
  NOR2_X1   g0588(.A1(new_n404), .A2(new_n654), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n654), .B1(new_n402), .B2(new_n403), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT100), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g0592(.A(KEYINPUT100), .B(new_n654), .C1(new_n402), .C2(new_n403), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n792), .A2(new_n793), .A3(new_n409), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n789), .B1(new_n794), .B2(new_n404), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n715), .A2(new_n796), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n795), .B(new_n655), .C1(new_n637), .C2(new_n626), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n702), .B(new_n799), .Z(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n742), .ZN(new_n801));
  INV_X1    g0601(.A(G294), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n758), .A2(new_n802), .B1(new_n770), .B2(new_n591), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n285), .B1(new_n749), .B2(G303), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n804), .B1(new_n455), .B2(new_n768), .C1(new_n771), .C2(new_n744), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n803), .B(new_n805), .C1(G311), .C2(new_n773), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n806), .B1(new_n466), .B2(new_n764), .C1(new_n211), .C2(new_n754), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT97), .Z(new_n808));
  NOR2_X1   g0608(.A1(new_n768), .A2(new_n216), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n749), .A2(G137), .B1(new_n755), .B2(G159), .ZN(new_n810));
  INV_X1    g0610(.A(G143), .ZN(new_n811));
  INV_X1    g0611(.A(G150), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n810), .B1(new_n811), .B2(new_n758), .C1(new_n812), .C2(new_n744), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT98), .Z(new_n814));
  OR2_X1    g0614(.A1(new_n814), .A2(KEYINPUT34), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(KEYINPUT34), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n278), .B1(new_n773), .B2(G132), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT99), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n764), .A2(new_n209), .B1(new_n352), .B2(new_n770), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n815), .A2(new_n816), .A3(new_n819), .A4(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n808), .B1(new_n809), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n742), .B1(new_n824), .B2(new_n739), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n739), .A2(new_n736), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n825), .B1(G77), .B2(new_n827), .C1(new_n737), .C2(new_n795), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n801), .A2(new_n828), .ZN(G384));
  INV_X1    g0629(.A(KEYINPUT38), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT37), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n338), .B(new_n344), .C1(new_n364), .C2(new_n359), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n371), .A2(KEYINPUT16), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n344), .B1(new_n359), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n377), .A2(new_n378), .A3(new_n652), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n831), .B1(new_n832), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n365), .A2(new_n835), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n832), .A2(new_n838), .A3(new_n831), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(KEYINPUT104), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT104), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n832), .A2(new_n838), .A3(new_n841), .A4(new_n831), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n837), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n652), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n834), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(new_n375), .B2(new_n384), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n830), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(KEYINPUT105), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n840), .A2(new_n842), .ZN(new_n849));
  INV_X1    g0649(.A(new_n837), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n851), .B(KEYINPUT38), .C1(new_n386), .C2(new_n845), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT105), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n853), .B(new_n830), .C1(new_n843), .C2(new_n846), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n848), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT39), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT107), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT39), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT106), .ZN(new_n859));
  INV_X1    g0659(.A(new_n367), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n327), .B1(new_n832), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n327), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n373), .B2(new_n338), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n859), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(KEYINPUT106), .B(new_n366), .C1(new_n374), .C2(new_n327), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n864), .A2(new_n384), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n373), .A2(new_n652), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n832), .A2(new_n838), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT37), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n866), .A2(new_n867), .B1(new_n849), .B2(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n852), .B(new_n858), .C1(new_n870), .C2(KEYINPUT38), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n856), .A2(new_n857), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n857), .B1(new_n856), .B2(new_n871), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n447), .A2(new_n437), .A3(new_n655), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n437), .A2(new_n654), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n877), .B(KEYINPUT102), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n641), .A2(new_n440), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT103), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n448), .A2(KEYINPUT103), .A3(new_n878), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n641), .A2(new_n655), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n789), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n883), .A2(new_n885), .B1(new_n798), .B2(new_n886), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n874), .A2(new_n876), .B1(new_n855), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n385), .A2(new_n652), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n450), .A2(new_n716), .A3(new_n714), .A4(new_n717), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n644), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n890), .B(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n882), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT103), .B1(new_n448), .B2(new_n878), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n885), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n607), .A2(new_n654), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n896), .B(new_n795), .C1(new_n697), .C2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n852), .B1(new_n870), .B2(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT40), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  INV_X1    g0702(.A(new_n855), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n902), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n697), .A2(new_n897), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n451), .A2(new_n906), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n905), .B(new_n907), .Z(new_n908));
  INV_X1    g0708(.A(G330), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n893), .B(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n255), .B2(new_n722), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n211), .B1(new_n458), .B2(KEYINPUT35), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n913), .B(new_n232), .C1(KEYINPUT35), .C2(new_n458), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT36), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n399), .A2(new_n235), .A3(new_n353), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n916), .B(KEYINPUT101), .Z(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n352), .B2(new_n201), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(G1), .A3(new_n646), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n912), .A2(new_n915), .A3(new_n919), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(KEYINPUT108), .Z(G367));
  AND2_X1   g0721(.A1(new_n773), .A2(G137), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n278), .B1(new_n755), .B2(new_n201), .ZN(new_n923));
  INV_X1    g0723(.A(G159), .ZN(new_n924));
  OAI221_X1 g0724(.A(new_n923), .B1(new_n924), .B2(new_n744), .C1(new_n399), .C2(new_n770), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n765), .A2(G68), .ZN(new_n926));
  OAI221_X1 g0726(.A(new_n926), .B1(new_n811), .B2(new_n748), .C1(new_n812), .C2(new_n758), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n922), .B(new_n925), .C1(new_n927), .C2(KEYINPUT110), .ZN(new_n928));
  OAI221_X1 g0728(.A(new_n928), .B1(KEYINPUT110), .B2(new_n927), .C1(new_n209), .C2(new_n768), .ZN(new_n929));
  INV_X1    g0729(.A(new_n768), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT46), .B1(new_n930), .B2(G116), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n930), .A2(KEYINPUT46), .A3(G116), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n802), .B2(new_n744), .ZN(new_n933));
  XOR2_X1   g0733(.A(KEYINPUT109), .B(G311), .Z(new_n934));
  AOI211_X1 g0734(.A(new_n931), .B(new_n933), .C1(new_n749), .C2(new_n934), .ZN(new_n935));
  OAI221_X1 g0735(.A(new_n278), .B1(new_n754), .B2(new_n771), .C1(new_n769), .C2(new_n758), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(G317), .B2(new_n773), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n938), .B1(new_n466), .B2(new_n770), .C1(new_n455), .C2(new_n764), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n929), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT47), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n742), .B1(new_n941), .B2(new_n739), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n245), .A2(new_n729), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n943), .B(new_n740), .C1(new_n227), .C2(new_n394), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n619), .A2(new_n655), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(new_n605), .A3(new_n620), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n706), .B2(new_n945), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n942), .B(new_n944), .C1(new_n786), .C2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n723), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n468), .A2(new_n654), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n499), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n492), .B2(new_n655), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n669), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT45), .Z(new_n954));
  NOR2_X1   g0754(.A1(new_n669), .A2(new_n952), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT44), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n665), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n957), .B(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n666), .B(new_n664), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n660), .B(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n720), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n674), .B(KEYINPUT41), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n949), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n668), .A2(new_n952), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT42), .Z(new_n966));
  OAI21_X1  g0766(.A(new_n492), .B1(new_n951), .B2(new_n537), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n655), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n966), .A2(new_n968), .B1(KEYINPUT43), .B2(new_n947), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n958), .A2(new_n952), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n969), .B(new_n970), .Z(new_n971));
  NOR2_X1   g0771(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n948), .B1(new_n964), .B2(new_n973), .ZN(G387));
  AND2_X1   g0774(.A1(new_n773), .A2(G326), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n749), .A2(G322), .B1(new_n755), .B2(G303), .ZN(new_n976));
  INV_X1    g0776(.A(new_n744), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n934), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n976), .B(new_n978), .C1(new_n745), .C2(new_n758), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT48), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(new_n771), .B2(new_n764), .C1(new_n802), .C2(new_n768), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT49), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n285), .B(new_n975), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n983), .B1(new_n982), .B2(new_n981), .C1(new_n211), .C2(new_n770), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n758), .A2(new_n216), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n930), .A2(new_n221), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n352), .B2(new_n754), .ZN(new_n987));
  XNOR2_X1  g0787(.A(KEYINPUT111), .B(G150), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n987), .B1(new_n773), .B2(new_n988), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n748), .A2(new_n924), .B1(new_n770), .B2(new_n466), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n278), .B(new_n990), .C1(new_n341), .C2(new_n977), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n764), .A2(new_n602), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n989), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n984), .B1(new_n985), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n742), .B1(new_n994), .B2(new_n739), .ZN(new_n995));
  OR3_X1    g0795(.A1(new_n272), .A2(KEYINPUT50), .A3(G50), .ZN(new_n996));
  OAI21_X1  g0796(.A(KEYINPUT50), .B1(new_n272), .B2(G50), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n996), .A2(new_n997), .A3(new_n297), .A4(new_n676), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G68), .B2(G77), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n729), .B1(new_n241), .B2(new_n297), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n285), .B(new_n227), .C1(G116), .C2(new_n592), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n227), .A2(G107), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n740), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n995), .B(new_n1004), .C1(new_n664), .C2(new_n786), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n961), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n674), .B1(new_n720), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n719), .A2(new_n961), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1005), .B1(new_n723), .B2(new_n961), .C1(new_n1007), .C2(new_n1008), .ZN(G393));
  XNOR2_X1  g0809(.A(new_n959), .B(new_n1008), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n674), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n959), .A2(new_n723), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n765), .A2(G77), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n773), .A2(G143), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n977), .A2(new_n201), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n285), .B1(new_n770), .B2(new_n591), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G68), .B2(new_n930), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n748), .A2(new_n812), .B1(new_n758), .B2(new_n924), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT114), .Z(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT113), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT51), .Z(new_n1022));
  AOI211_X1 g0822(.A(new_n1018), .B(new_n1022), .C1(new_n341), .C2(new_n755), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n749), .A2(G317), .B1(new_n759), .B2(G311), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT52), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n278), .B1(new_n754), .B2(new_n802), .C1(new_n455), .C2(new_n770), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G303), .B2(new_n977), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n773), .A2(G322), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(new_n771), .C2(new_n768), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1025), .B(new_n1029), .C1(G116), .C2(new_n765), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n739), .B1(new_n1023), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n729), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n740), .B1(new_n466), .B2(new_n227), .C1(new_n249), .C2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n725), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT112), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1031), .B(new_n1035), .C1(new_n786), .C2(new_n952), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1011), .A2(new_n1012), .A3(new_n1036), .ZN(G390));
  OAI21_X1  g0837(.A(new_n278), .B1(new_n744), .B2(new_n455), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n778), .B(new_n1038), .C1(G283), .C2(new_n749), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n755), .A2(G97), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n758), .A2(new_n211), .B1(new_n770), .B2(new_n352), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G294), .B2(new_n773), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1039), .A2(new_n1013), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n930), .A2(new_n988), .ZN(new_n1044));
  INV_X1    g0844(.A(G128), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n1044), .A2(KEYINPUT53), .B1(new_n1045), .B2(new_n748), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(KEYINPUT53), .B2(new_n1044), .ZN(new_n1047));
  INV_X1    g0847(.A(G132), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n285), .B1(new_n758), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n773), .B2(G125), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n924), .B2(new_n764), .C1(new_n202), .C2(new_n770), .ZN(new_n1052));
  INV_X1    g0852(.A(G137), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(KEYINPUT54), .B(G143), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n744), .A2(new_n1053), .B1(new_n754), .B2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT118), .Z(new_n1056));
  OAI21_X1  g0856(.A(new_n1043), .B1(new_n1052), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n742), .B1(new_n1057), .B2(new_n739), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n341), .B2(new_n827), .C1(new_n874), .C2(new_n737), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n899), .A2(new_n875), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n794), .A2(new_n404), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n655), .B(new_n1061), .C1(new_n703), .C2(new_n710), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n883), .A2(new_n885), .B1(new_n1062), .B2(new_n886), .ZN(new_n1063));
  OAI21_X1  g0863(.A(KEYINPUT115), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1062), .A2(new_n886), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n896), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT115), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1066), .A2(new_n1067), .A3(new_n875), .A4(new_n899), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n872), .A2(new_n873), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT116), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n887), .B2(new_n876), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n798), .A2(new_n886), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n896), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1074), .A2(KEYINPUT116), .A3(new_n875), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1069), .B1(new_n1070), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n896), .ZN(new_n1078));
  NOR4_X1   g0878(.A1(new_n906), .A2(new_n1078), .A3(new_n909), .A4(new_n796), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(KEYINPUT117), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n796), .A2(new_n909), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n701), .A2(new_n896), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1077), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT117), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1086), .A2(new_n872), .A3(new_n873), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1085), .B(new_n1079), .C1(new_n1087), .C2(new_n1069), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1081), .A2(new_n1084), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1059), .B1(new_n1089), .B2(new_n723), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n450), .B(G330), .C1(new_n897), .C2(new_n697), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1091), .A2(new_n891), .A3(new_n644), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n896), .B1(new_n701), .B2(new_n1082), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1073), .B1(new_n1093), .B2(new_n1079), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1065), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n906), .A2(new_n909), .A3(new_n796), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1083), .B(new_n1095), .C1(new_n1096), .C2(new_n896), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1092), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1081), .A2(new_n1084), .A3(new_n1088), .A4(new_n1098), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1099), .A2(new_n674), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1098), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1089), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1090), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(G378));
  XNOR2_X1  g0904(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n324), .A2(KEYINPUT55), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n640), .B1(new_n316), .B2(new_n318), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT55), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n274), .A2(new_n652), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1107), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1112), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1106), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1115), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1117), .A2(new_n1105), .A3(new_n1113), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n736), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n826), .A2(new_n202), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n744), .A2(new_n1048), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n758), .A2(new_n1045), .B1(new_n754), .B2(new_n1053), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1122), .B(new_n1123), .C1(G125), .C2(new_n749), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n1124), .B1(new_n812), .B2(new_n764), .C1(new_n768), .C2(new_n1054), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(KEYINPUT59), .ZN(new_n1126));
  AOI211_X1 g0926(.A(G33), .B(G41), .C1(new_n773), .C2(G124), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1128), .B1(KEYINPUT59), .B2(new_n1125), .C1(new_n924), .C2(new_n770), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n773), .A2(G283), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n672), .A2(new_n285), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n753), .A2(new_n767), .A3(G58), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1130), .A2(new_n986), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT119), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n602), .A2(new_n754), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n758), .A2(new_n455), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT120), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n977), .A2(G97), .ZN(new_n1138));
  AND4_X1   g0938(.A1(new_n926), .A2(new_n1135), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1134), .B(new_n1139), .C1(new_n211), .C2(new_n748), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT58), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1129), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1143), .B1(new_n1141), .B2(new_n1140), .C1(new_n1131), .C2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n742), .B1(new_n1145), .B2(new_n739), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1120), .A2(new_n1121), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1119), .B1(new_n905), .B2(new_n909), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1149), .A2(G330), .A3(new_n904), .A4(new_n901), .ZN(new_n1150));
  AND4_X1   g0950(.A1(new_n889), .A2(new_n1148), .A3(new_n888), .A4(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1150), .A2(new_n1148), .B1(new_n888), .B2(new_n889), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1147), .B1(new_n1153), .B2(new_n723), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT122), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1092), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1099), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1156), .B1(new_n1099), .B2(new_n1157), .ZN(new_n1159));
  NOR3_X1   g0959(.A1(new_n1158), .A2(new_n1159), .A3(new_n1153), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n674), .B1(new_n1160), .B2(KEYINPUT57), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1099), .A2(new_n1157), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(KEYINPUT122), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1099), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT57), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1155), .B1(new_n1161), .B2(new_n1168), .ZN(G375));
  OAI21_X1  g0969(.A(new_n1132), .B1(new_n744), .B2(new_n1054), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n278), .B(new_n1170), .C1(G132), .C2(new_n749), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n768), .A2(new_n924), .B1(new_n754), .B2(new_n812), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G128), .B2(new_n773), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1171), .B(new_n1173), .C1(new_n216), .C2(new_n764), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G137), .B2(new_n759), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n278), .B1(new_n744), .B2(new_n211), .C1(new_n802), .C2(new_n748), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G107), .B2(new_n755), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n758), .A2(new_n771), .B1(new_n770), .B2(new_n206), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G303), .B2(new_n773), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1177), .A2(new_n992), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G97), .B2(new_n930), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n739), .B1(new_n1175), .B2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1182), .B(new_n725), .C1(G68), .C2(new_n827), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT124), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n896), .A2(new_n737), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1186), .B1(new_n1187), .B2(KEYINPUT123), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1185), .B(new_n1188), .C1(KEYINPUT123), .C2(new_n1187), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1189), .B1(new_n1190), .B2(new_n949), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1094), .A2(new_n1097), .A3(new_n1092), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n963), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1191), .B1(new_n1193), .B2(new_n1098), .ZN(G381));
  NOR2_X1   g0994(.A1(G375), .A2(G378), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(G381), .A2(G393), .A3(G396), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(G390), .A2(G387), .A3(G384), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(G407));
  INV_X1    g0998(.A(G213), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n1195), .B2(new_n653), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(G407), .ZN(G409));
  NOR2_X1   g1001(.A1(new_n1199), .A2(G343), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1192), .A2(KEYINPUT125), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n675), .B1(new_n1204), .B2(KEYINPUT60), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1205), .B(new_n1101), .C1(KEYINPUT60), .C2(new_n1204), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n1191), .ZN(new_n1207));
  INV_X1    g1007(.A(G384), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1207), .B(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n675), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1160), .A2(KEYINPUT57), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1103), .B(new_n1154), .C1(new_n1211), .C2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1160), .A2(new_n963), .ZN(new_n1214));
  AOI21_X1  g1014(.A(G378), .B1(new_n1214), .B2(new_n1155), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1203), .B(new_n1210), .C1(new_n1213), .C2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(KEYINPUT62), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT61), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1202), .A2(G2897), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1209), .B(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1154), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1215), .B1(new_n1221), .B2(G378), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1220), .B1(new_n1222), .B2(new_n1202), .ZN(new_n1223));
  OAI211_X1 g1023(.A(G378), .B(new_n1155), .C1(new_n1161), .C2(new_n1168), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1215), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT62), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1226), .A2(new_n1227), .A3(new_n1203), .A4(new_n1210), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1217), .A2(new_n1218), .A3(new_n1223), .A4(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(G387), .A2(KEYINPUT126), .ZN(new_n1230));
  XOR2_X1   g1030(.A(G393), .B(G396), .Z(new_n1231));
  MUX2_X1   g1031(.A(new_n1230), .B(G387), .S(new_n1231), .Z(new_n1232));
  INV_X1    g1032(.A(G390), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1229), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT61), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1226), .A2(KEYINPUT63), .A3(new_n1203), .A4(new_n1210), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT63), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1226), .A2(new_n1203), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1240), .B1(new_n1241), .B2(new_n1220), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1216), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1238), .B(new_n1239), .C1(new_n1242), .C2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1237), .A2(new_n1244), .ZN(G405));
  NAND3_X1  g1045(.A1(G375), .A2(new_n1103), .A3(new_n1210), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1209), .B1(new_n1221), .B2(G378), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1248), .A2(KEYINPUT127), .A3(new_n1224), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1224), .A2(KEYINPUT127), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1246), .A2(new_n1250), .A3(new_n1247), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1249), .A2(new_n1236), .A3(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1236), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(G402));
endmodule


