//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n439, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n579, new_n580, new_n581,
    new_n582, new_n584, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1178, new_n1179,
    new_n1180;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G69), .ZN(new_n439));
  INV_X1    g014(.A(new_n439), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n439), .A2(G57), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(new_n454));
  NAND4_X1  g029(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G2106), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(G137), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT68), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n463), .A2(new_n465), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(new_n472), .A3(G137), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n462), .A2(G2105), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n469), .A2(new_n473), .B1(G101), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n466), .A2(KEYINPUT67), .A3(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n478));
  INV_X1    g053(.A(G125), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n478), .B1(new_n470), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n475), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  NOR2_X1   g059(.A1(new_n470), .A2(new_n467), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n471), .A2(G136), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND2_X1  g066(.A1(G114), .A2(G2104), .ZN(new_n492));
  INV_X1    g067(.A(G126), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n470), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n471), .A2(G138), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n466), .A2(KEYINPUT4), .A3(G138), .ZN(new_n498));
  NAND2_X1  g073(.A1(G102), .A2(G2104), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n496), .A2(new_n497), .B1(new_n467), .B2(new_n500), .ZN(G164));
  NAND2_X1  g076(.A1(G75), .A2(G543), .ZN(new_n502));
  XNOR2_X1  g077(.A(new_n502), .B(KEYINPUT70), .ZN(new_n503));
  INV_X1    g078(.A(G62), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n503), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n505), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n510), .A2(G651), .B1(G50), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  OAI211_X1 g092(.A(new_n506), .B(new_n508), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n511), .A2(new_n512), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT5), .B(G543), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT69), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n514), .B1(new_n515), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(KEYINPUT71), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(KEYINPUT71), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(G166));
  NAND2_X1  g104(.A1(new_n513), .A2(G51), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n522), .A2(G63), .A3(G651), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n520), .A2(G89), .A3(new_n523), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n509), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n540), .A2(G651), .B1(G52), .B2(new_n513), .ZN(new_n541));
  XOR2_X1   g116(.A(KEYINPUT72), .B(G90), .Z(new_n542));
  NAND3_X1  g117(.A1(new_n520), .A2(new_n523), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(G171));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n509), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G651), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n520), .A2(G81), .A3(new_n523), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT73), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n513), .A2(G43), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n551), .B1(new_n550), .B2(new_n552), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n549), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(KEYINPUT74), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT74), .ZN(new_n557));
  OAI211_X1 g132(.A(new_n557), .B(new_n549), .C1(new_n553), .C2(new_n554), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT75), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT76), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n561), .A2(new_n566), .ZN(G188));
  NAND3_X1  g142(.A1(new_n520), .A2(G91), .A3(new_n523), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n509), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G651), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT9), .ZN(new_n573));
  OAI21_X1  g148(.A(G543), .B1(new_n516), .B2(new_n517), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n513), .A2(KEYINPUT9), .A3(G53), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n568), .A2(new_n572), .A3(new_n576), .A4(new_n577), .ZN(G299));
  NAND3_X1  g153(.A1(new_n541), .A2(KEYINPUT77), .A3(new_n543), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(KEYINPUT77), .B1(new_n541), .B2(new_n543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G301));
  INV_X1    g158(.A(new_n528), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n526), .ZN(G303));
  AND2_X1   g160(.A1(new_n520), .A2(new_n523), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT78), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n586), .A2(new_n587), .A3(G87), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n522), .A2(G74), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(new_n513), .B2(G49), .ZN(new_n590));
  INV_X1    g165(.A(G87), .ZN(new_n591));
  OAI21_X1  g166(.A(KEYINPUT78), .B1(new_n524), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n588), .A2(new_n590), .A3(new_n592), .ZN(G288));
  NAND2_X1  g168(.A1(new_n586), .A2(G86), .ZN(new_n594));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G61), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n509), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(G48), .B2(new_n513), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n594), .A2(new_n598), .ZN(G305));
  NAND2_X1  g174(.A1(new_n586), .A2(G85), .ZN(new_n600));
  NAND2_X1  g175(.A1(G72), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G60), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n509), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(G47), .B2(new_n513), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(G290));
  NAND3_X1  g180(.A1(new_n520), .A2(G92), .A3(new_n523), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G66), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n509), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G651), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n513), .A2(KEYINPUT79), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT79), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n574), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n612), .A2(new_n614), .A3(G54), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  NAND4_X1  g191(.A1(new_n520), .A2(new_n523), .A3(new_n616), .A4(G92), .ZN(new_n617));
  NAND4_X1  g192(.A1(new_n607), .A2(new_n611), .A3(new_n615), .A4(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n582), .B2(new_n619), .ZN(G284));
  OAI21_X1  g196(.A(new_n620), .B1(new_n582), .B2(new_n619), .ZN(G321));
  NAND2_X1  g197(.A1(G299), .A2(new_n619), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G168), .B2(new_n619), .ZN(G297));
  XOR2_X1   g199(.A(G297), .B(KEYINPUT80), .Z(G280));
  INV_X1    g200(.A(new_n618), .ZN(new_n626));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G860), .ZN(G148));
  NOR2_X1   g203(.A1(new_n618), .A2(G559), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G868), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n559), .B2(G868), .ZN(G323));
  XNOR2_X1  g207(.A(KEYINPUT81), .B(KEYINPUT11), .ZN(new_n633));
  XNOR2_X1  g208(.A(G323), .B(new_n633), .ZN(G282));
  NAND2_X1  g209(.A1(new_n466), .A2(new_n474), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2100), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n485), .A2(G123), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n471), .A2(G135), .ZN(new_n640));
  OR2_X1    g215(.A1(G99), .A2(G2105), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n641), .B(G2104), .C1(G111), .C2(new_n467), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n638), .A2(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2435), .ZN(new_n647));
  XOR2_X1   g222(.A(G2427), .B(G2438), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT14), .ZN(new_n650));
  XOR2_X1   g225(.A(G2451), .B(G2454), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G1341), .B(G1348), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(G14), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(G401));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  XOR2_X1   g235(.A(G2067), .B(G2678), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n660), .B1(new_n664), .B2(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2096), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2100), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n662), .A2(new_n663), .ZN(new_n669));
  AOI21_X1  g244(.A(KEYINPUT18), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n667), .B(new_n670), .Z(G227));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT82), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1971), .B(G1976), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT20), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n673), .A2(new_n674), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(new_n679), .B2(new_n675), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(KEYINPUT83), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(G1986), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1991), .B(G1996), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT22), .B(G1981), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(G229));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G5), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G171), .B2(new_n693), .ZN(new_n695));
  INV_X1    g270(.A(G1961), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n643), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(G35), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G162), .B2(new_n698), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT29), .Z(new_n702));
  INV_X1    g277(.A(G2090), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT31), .B(G11), .ZN(new_n705));
  OR2_X1    g280(.A1(G29), .A2(G33), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n474), .A2(G103), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT25), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n471), .A2(G139), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n708), .B(new_n709), .C1(new_n467), .C2(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n706), .B1(new_n711), .B2(new_n698), .ZN(new_n712));
  INV_X1    g287(.A(G2072), .ZN(new_n713));
  OR2_X1    g288(.A1(G29), .A2(G32), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n471), .A2(G141), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n485), .A2(G129), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n474), .A2(G105), .ZN(new_n717));
  NAND3_X1  g292(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT26), .Z(new_n719));
  NAND4_X1  g294(.A1(new_n715), .A2(new_n716), .A3(new_n717), .A4(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n714), .B1(new_n720), .B2(new_n698), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT27), .B(G1996), .Z(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n712), .A2(new_n713), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT30), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(G28), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(G28), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n726), .A2(new_n727), .A3(new_n698), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n704), .A2(new_n705), .A3(new_n724), .A4(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n721), .ZN(new_n730));
  AOI211_X1 g305(.A(new_n699), .B(new_n729), .C1(new_n730), .C2(new_n722), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n693), .A2(G21), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G168), .B2(new_n693), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1966), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n626), .A2(G16), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G4), .B2(G16), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT89), .B(G1348), .Z(new_n738));
  AOI21_X1  g313(.A(new_n734), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G160), .A2(new_n698), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT24), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(G34), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(G34), .ZN(new_n743));
  AOI21_X1  g318(.A(G29), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(G2084), .B1(new_n740), .B2(new_n744), .ZN(new_n745));
  AND2_X1   g320(.A1(KEYINPUT85), .A2(G16), .ZN(new_n746));
  NOR2_X1   g321(.A1(KEYINPUT85), .A2(G16), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n749), .A2(KEYINPUT23), .A3(G20), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT23), .ZN(new_n751));
  INV_X1    g326(.A(G20), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n748), .B2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G299), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n750), .B(new_n753), .C1(new_n754), .C2(new_n693), .ZN(new_n755));
  INV_X1    g330(.A(G1956), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n702), .B2(new_n703), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT94), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n731), .A2(new_n739), .A3(new_n745), .A4(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n712), .A2(new_n713), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT92), .Z(new_n762));
  NOR2_X1   g337(.A1(new_n740), .A2(new_n744), .ZN(new_n763));
  INV_X1    g338(.A(G2084), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G27), .ZN(new_n766));
  OAI21_X1  g341(.A(KEYINPUT93), .B1(new_n766), .B2(G29), .ZN(new_n767));
  OR3_X1    g342(.A1(new_n766), .A2(KEYINPUT93), .A3(G29), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n767), .B(new_n768), .C1(G164), .C2(new_n698), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n765), .B1(G2078), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G2078), .B2(new_n769), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n737), .A2(new_n738), .ZN(new_n773));
  NOR4_X1   g348(.A1(new_n760), .A2(new_n762), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n693), .A2(G23), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT87), .ZN(new_n776));
  XNOR2_X1  g351(.A(G288), .B(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n775), .B1(new_n777), .B2(new_n693), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT88), .B(KEYINPUT33), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1976), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n778), .B(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n748), .A2(G22), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G166), .B2(new_n748), .ZN(new_n783));
  INV_X1    g358(.A(G1971), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n693), .A2(G6), .ZN(new_n786));
  INV_X1    g361(.A(G305), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(new_n693), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT32), .B(G1981), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n781), .A2(new_n785), .A3(new_n790), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT34), .Z(new_n792));
  INV_X1    g367(.A(KEYINPUT36), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n749), .A2(G24), .ZN(new_n794));
  INV_X1    g369(.A(G290), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n749), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT86), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1986), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n698), .A2(G25), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n471), .A2(G131), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT84), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n485), .A2(G119), .ZN(new_n802));
  NOR2_X1   g377(.A1(G95), .A2(G2105), .ZN(new_n803));
  OAI21_X1  g378(.A(G2104), .B1(new_n467), .B2(G107), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n799), .B1(new_n806), .B2(new_n698), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT35), .B(G1991), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  NOR3_X1   g385(.A1(new_n798), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n792), .A2(new_n793), .A3(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n793), .B1(new_n792), .B2(new_n811), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n697), .B(new_n774), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n698), .A2(G26), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n471), .A2(G140), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT90), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n485), .A2(G128), .ZN(new_n820));
  OR2_X1    g395(.A1(G104), .A2(G2105), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n821), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n471), .A2(KEYINPUT90), .A3(G140), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n819), .A2(new_n820), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT91), .Z(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n816), .B1(new_n826), .B2(new_n698), .ZN(new_n827));
  MUX2_X1   g402(.A(new_n816), .B(new_n827), .S(KEYINPUT28), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G2067), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n559), .A2(new_n748), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(G19), .B2(new_n748), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(G1341), .Z(new_n832));
  NOR3_X1   g407(.A1(new_n815), .A2(new_n829), .A3(new_n832), .ZN(G311));
  INV_X1    g408(.A(new_n774), .ZN(new_n834));
  INV_X1    g409(.A(new_n814), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(new_n812), .ZN(new_n836));
  INV_X1    g411(.A(new_n829), .ZN(new_n837));
  INV_X1    g412(.A(new_n832), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n836), .A2(new_n837), .A3(new_n838), .A4(new_n697), .ZN(G150));
  NAND3_X1  g414(.A1(new_n520), .A2(G93), .A3(new_n523), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT97), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n513), .A2(G55), .ZN(new_n842));
  AND3_X1   g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n841), .B1(new_n840), .B2(new_n842), .ZN(new_n844));
  NAND2_X1  g419(.A1(G80), .A2(G543), .ZN(new_n845));
  INV_X1    g420(.A(G67), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n509), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(KEYINPUT96), .B1(new_n847), .B2(G651), .ZN(new_n848));
  AND3_X1   g423(.A1(new_n847), .A2(KEYINPUT96), .A3(G651), .ZN(new_n849));
  OAI22_X1  g424(.A1(new_n843), .A2(new_n844), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G860), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT99), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT37), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n559), .A2(new_n850), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n550), .A2(new_n552), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(KEYINPUT73), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n857), .A2(new_n858), .B1(G651), .B2(new_n548), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n855), .B1(new_n859), .B2(new_n850), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n849), .A2(new_n848), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n840), .A2(new_n842), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT97), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n865), .A2(new_n555), .A3(KEYINPUT98), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n860), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n854), .A2(new_n867), .ZN(new_n868));
  XOR2_X1   g443(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n626), .A2(G559), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT39), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n870), .B(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n853), .B1(new_n873), .B2(G860), .ZN(G145));
  XNOR2_X1  g449(.A(new_n806), .B(new_n636), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(new_n711), .Z(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n490), .B(KEYINPUT100), .ZN(new_n878));
  INV_X1    g453(.A(new_n643), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n878), .A2(new_n879), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n483), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NOR3_X1   g458(.A1(new_n880), .A2(new_n881), .A3(new_n483), .ZN(new_n884));
  NOR3_X1   g459(.A1(new_n883), .A2(new_n826), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n826), .B1(new_n883), .B2(new_n884), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n877), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n876), .B1(new_n889), .B2(new_n885), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  AOI22_X1  g466(.A1(G130), .A2(new_n485), .B1(new_n471), .B2(G142), .ZN(new_n892));
  OAI21_X1  g467(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n467), .A2(G118), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT101), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n892), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n720), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(G164), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n891), .B(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G37), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(new_n865), .B2(G868), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n868), .A2(new_n629), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n630), .B1(new_n854), .B2(new_n867), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n618), .A2(new_n754), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n615), .A2(new_n611), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n909), .A2(G299), .A3(new_n607), .A4(new_n617), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT102), .B1(new_n907), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT41), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n914), .B1(new_n911), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n911), .A2(new_n915), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n911), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n908), .A2(KEYINPUT103), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n917), .B1(new_n921), .B2(new_n915), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n916), .B1(new_n922), .B2(new_n914), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n907), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n925), .B(new_n911), .C1(new_n905), .C2(new_n906), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n913), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT42), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n777), .A2(new_n795), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n777), .A2(new_n795), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(G303), .A2(G305), .ZN(new_n932));
  NAND2_X1  g507(.A1(G166), .A2(new_n787), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n932), .A2(new_n933), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n930), .B2(new_n929), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n913), .A2(new_n939), .A3(new_n924), .A4(new_n926), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n928), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n938), .B1(new_n928), .B2(new_n940), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n904), .B1(new_n943), .B2(G868), .ZN(new_n944));
  NOR4_X1   g519(.A1(new_n941), .A2(new_n942), .A3(new_n903), .A4(new_n619), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(G295));
  NOR2_X1   g521(.A1(new_n944), .A2(new_n945), .ZN(G331));
  NAND2_X1  g522(.A1(new_n938), .A2(KEYINPUT109), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n935), .A2(new_n937), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT77), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n544), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(G286), .B1(new_n953), .B2(new_n579), .ZN(new_n954));
  NOR2_X1   g529(.A1(G168), .A2(new_n544), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT107), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(KEYINPUT107), .B2(new_n955), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n865), .A2(KEYINPUT98), .A3(new_n555), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT98), .B1(new_n865), .B2(new_n555), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n865), .B1(new_n556), .B2(new_n558), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n955), .A2(KEYINPUT107), .ZN(new_n964));
  NAND2_X1  g539(.A1(G171), .A2(G286), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(new_n582), .B2(G286), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n964), .B1(new_n966), .B2(KEYINPUT107), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n967), .A2(new_n854), .A3(new_n867), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n962), .A2(new_n963), .A3(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n967), .A2(new_n854), .A3(new_n867), .A4(KEYINPUT108), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n923), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n962), .A2(new_n911), .A3(new_n968), .ZN(new_n972));
  AOI22_X1  g547(.A1(new_n948), .A2(new_n951), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(new_n949), .A3(new_n972), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n900), .ZN(new_n975));
  OR4_X1    g550(.A1(KEYINPUT112), .A2(new_n973), .A3(new_n975), .A4(KEYINPUT43), .ZN(new_n976));
  INV_X1    g551(.A(new_n973), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n974), .A2(new_n900), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT112), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n969), .A2(new_n970), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(new_n983), .B2(new_n911), .ZN(new_n984));
  AOI211_X1 g559(.A(KEYINPUT110), .B(new_n912), .C1(new_n969), .C2(new_n970), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n915), .B1(new_n919), .B2(new_n920), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n911), .A2(KEYINPUT41), .ZN(new_n987));
  AOI211_X1 g562(.A(new_n986), .B(new_n987), .C1(new_n962), .C2(new_n968), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n984), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n948), .A2(new_n951), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n978), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n976), .A2(new_n981), .A3(KEYINPUT44), .A4(new_n992), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n979), .B(new_n978), .C1(new_n989), .C2(new_n990), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT43), .B1(new_n973), .B2(new_n975), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT111), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n1000));
  AOI211_X1 g575(.A(new_n1000), .B(new_n997), .C1(new_n994), .C2(new_n995), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n993), .B1(new_n999), .B2(new_n1001), .ZN(G397));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n1003));
  INV_X1    g578(.A(G40), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1003), .B1(new_n483), .B2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n475), .A2(new_n482), .A3(KEYINPUT113), .A4(G40), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(G164), .B2(G1384), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n825), .B(G2067), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(new_n720), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n1007), .A2(G1996), .A3(new_n1009), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n1013), .A2(KEYINPUT46), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(KEYINPUT46), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT126), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT47), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n720), .B(G1996), .ZN(new_n1019));
  OR2_X1    g594(.A1(new_n1011), .A2(new_n1019), .ZN(new_n1020));
  OR3_X1    g595(.A1(new_n801), .A2(new_n808), .A3(new_n805), .ZN(new_n1021));
  OAI22_X1  g596(.A1(new_n1020), .A2(new_n1021), .B1(G2067), .B2(new_n825), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n1010), .ZN(new_n1023));
  XOR2_X1   g598(.A(new_n806), .B(new_n808), .Z(new_n1024));
  OAI21_X1  g599(.A(new_n1010), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  OR3_X1    g600(.A1(G290), .A2(KEYINPUT114), .A3(G1986), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT114), .B1(G290), .B2(G1986), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1010), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1028), .B(KEYINPUT48), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1018), .A2(new_n1023), .A3(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(G164), .A2(G1384), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1005), .A2(new_n1032), .A3(new_n1006), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(G8), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(G305), .A2(G1981), .ZN(new_n1036));
  XOR2_X1   g611(.A(KEYINPUT119), .B(G86), .Z(new_n1037));
  OAI21_X1  g612(.A(new_n598), .B1(new_n524), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1036), .B1(G1981), .B2(new_n1038), .ZN(new_n1039));
  XOR2_X1   g614(.A(new_n1039), .B(KEYINPUT49), .Z(new_n1040));
  AOI211_X1 g615(.A(G1976), .B(G288), .C1(new_n1040), .C2(new_n1035), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1035), .B1(new_n1041), .B2(new_n1036), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1034), .B1(G1976), .B2(new_n777), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n1044));
  INV_X1    g619(.A(G288), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1043), .B(new_n1044), .C1(G1976), .C2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT118), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1040), .A2(new_n1035), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT118), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1048), .B(new_n1049), .C1(new_n1050), .C2(new_n1046), .ZN(new_n1051));
  INV_X1    g626(.A(G8), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n496), .A2(new_n497), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n500), .A2(new_n467), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G1384), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(KEYINPUT50), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(G164), .B2(G1384), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(new_n1007), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n703), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1055), .A2(KEYINPUT45), .A3(new_n1056), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1005), .A2(new_n1064), .A3(new_n1009), .A4(new_n1006), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n784), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1052), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(G303), .A2(G8), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT117), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1071), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1067), .A2(new_n1073), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n1051), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1005), .A2(new_n1009), .A3(new_n1006), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT120), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1005), .A2(new_n1009), .A3(new_n1078), .A4(new_n1006), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(new_n1079), .A3(new_n1064), .ZN(new_n1080));
  INV_X1    g655(.A(G1966), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1062), .A2(new_n764), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1052), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(G168), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1067), .A2(new_n1073), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1074), .ZN(new_n1087));
  NOR4_X1   g662(.A1(new_n1051), .A2(new_n1085), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT63), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1042), .B(new_n1075), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1084), .A2(G286), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1082), .A2(G168), .A3(new_n1083), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1052), .A2(KEYINPUT124), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1092), .A2(KEYINPUT51), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT51), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1091), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT62), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1080), .A2(new_n1098), .A3(G2078), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n696), .B1(new_n1061), .B2(new_n1007), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1098), .B1(new_n1065), .B2(G2078), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n582), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT62), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1105), .B(new_n1091), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1097), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n756), .B1(new_n1061), .B2(new_n1007), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n1109));
  OAI21_X1  g684(.A(G299), .B1(KEYINPUT121), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(KEYINPUT121), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1110), .B(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT122), .B(G2072), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1113), .B(KEYINPUT56), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1108), .B(new_n1112), .C1(new_n1065), .C2(new_n1115), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n1062), .A2(G1348), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1033), .A2(KEYINPUT123), .ZN(new_n1118));
  INV_X1    g693(.A(G2067), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1005), .A2(new_n1120), .A3(new_n1032), .A4(new_n1006), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1118), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n618), .B1(new_n1117), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1112), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1125));
  AOI21_X1  g700(.A(G1956), .B1(new_n1125), .B2(new_n1060), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1065), .A2(new_n1115), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1124), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1116), .B1(new_n1123), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1122), .B1(G1348), .B2(new_n1062), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n618), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1117), .A2(new_n626), .A3(new_n1122), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1132), .A2(new_n1133), .A3(KEYINPUT60), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT58), .B(G1341), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1135), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1065), .A2(G1996), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n559), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT59), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1140), .B(new_n559), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1134), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1116), .A2(new_n1128), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1144), .B1(new_n1116), .B2(new_n1128), .ZN(new_n1146));
  OAI22_X1  g721(.A1(new_n1145), .A2(new_n1146), .B1(KEYINPUT60), .B2(new_n1133), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1130), .B1(new_n1143), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT54), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1009), .A2(G40), .A3(G160), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT125), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1098), .A2(G2078), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1152), .A2(new_n1064), .A3(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1100), .B(new_n1101), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1103), .B(new_n1149), .C1(new_n582), .C2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1158), .A2(G301), .B1(G171), .B2(new_n1156), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1157), .B1(new_n1159), .B2(new_n1149), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1148), .A2(new_n1160), .A3(new_n1096), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1084), .A2(new_n1089), .A3(G168), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1107), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1051), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1090), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1010), .A2(G1986), .A3(G290), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1028), .A2(new_n1166), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n1167), .B(KEYINPUT115), .Z(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1025), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1169), .B(KEYINPUT116), .Z(new_n1170));
  OAI21_X1  g745(.A(new_n1031), .B1(new_n1165), .B2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g746(.A(G319), .ZN(new_n1173));
  NOR2_X1   g747(.A1(G229), .A2(new_n1173), .ZN(new_n1174));
  OR2_X1    g748(.A1(G401), .A2(G227), .ZN(new_n1175));
  AOI21_X1  g749(.A(new_n1175), .B1(new_n899), .B2(new_n900), .ZN(new_n1176));
  NAND3_X1  g750(.A1(new_n996), .A2(new_n1174), .A3(new_n1176), .ZN(G225));
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n1178));
  NAND2_X1  g752(.A1(G225), .A2(new_n1178), .ZN(new_n1179));
  NAND4_X1  g753(.A1(new_n996), .A2(new_n1174), .A3(new_n1176), .A4(KEYINPUT127), .ZN(new_n1180));
  NAND2_X1  g754(.A1(new_n1179), .A2(new_n1180), .ZN(G308));
endmodule


