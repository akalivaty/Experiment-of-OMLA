//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n495, new_n496, new_n497, new_n498, new_n499, new_n500,
    new_n501, new_n502, new_n503, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n573, new_n575, new_n576, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n632,
    new_n634, new_n635, new_n636, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167, new_n1168;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT66), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT67), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT68), .Z(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT69), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(new_n455), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  AND3_X1   g042(.A1(new_n467), .A2(KEYINPUT72), .A3(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(KEYINPUT72), .B1(new_n467), .B2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT70), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT70), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G137), .ZN(new_n476));
  INV_X1    g051(.A(G101), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n471), .A2(G2104), .ZN(new_n478));
  OAI22_X1  g053(.A1(new_n470), .A2(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT73), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n478), .A2(new_n477), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n467), .A2(G2104), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT72), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n484), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n467), .A2(KEYINPUT72), .A3(G2104), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G137), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n472), .B2(new_n474), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n482), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT73), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n481), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n475), .ZN(new_n493));
  INV_X1    g068(.A(G125), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT71), .B1(new_n495), .B2(new_n483), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n467), .A2(G2104), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n497), .A2(new_n466), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g075(.A1(G113), .A2(G2104), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n493), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n492), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G160));
  NAND2_X1  g079(.A1(new_n487), .A2(new_n471), .ZN(new_n505));
  INV_X1    g080(.A(G136), .ZN(new_n506));
  OR3_X1    g081(.A1(new_n505), .A2(KEYINPUT74), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT74), .B1(new_n505), .B2(new_n506), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n470), .A2(new_n475), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G124), .ZN(new_n510));
  OAI221_X1 g085(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n475), .C2(G112), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n507), .A2(new_n508), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G162));
  INV_X1    g088(.A(new_n478), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G102), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT4), .ZN(new_n517));
  AOI211_X1 g092(.A(new_n517), .B(new_n483), .C1(new_n485), .C2(new_n486), .ZN(new_n518));
  INV_X1    g093(.A(G138), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n519), .B1(new_n472), .B2(new_n474), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n516), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g096(.A(G126), .B(new_n466), .C1(new_n468), .C2(new_n469), .ZN(new_n522));
  NAND2_X1  g097(.A1(G114), .A2(G2104), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G2105), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n497), .A2(new_n466), .A3(new_n498), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n498), .B1(new_n497), .B2(new_n466), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n520), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(new_n517), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n521), .A2(new_n525), .A3(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(G164));
  INV_X1    g106(.A(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT5), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT5), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G543), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n536), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G651), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n536), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n540));
  XOR2_X1   g115(.A(KEYINPUT6), .B(G651), .Z(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(G166));
  NAND3_X1  g118(.A1(new_n536), .A2(G63), .A3(G651), .ZN(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT7), .ZN(new_n546));
  XNOR2_X1  g121(.A(KEYINPUT6), .B(G651), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n536), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(G89), .ZN(new_n549));
  OAI211_X1 g124(.A(new_n544), .B(new_n546), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G51), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n541), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n547), .A2(KEYINPUT75), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n554), .A2(G543), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n551), .B1(new_n552), .B2(new_n556), .ZN(G286));
  INV_X1    g132(.A(G286), .ZN(G168));
  AND3_X1   g133(.A1(new_n554), .A2(G543), .A3(new_n555), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G52), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n536), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(new_n538), .ZN(new_n562));
  INV_X1    g137(.A(G90), .ZN(new_n563));
  OAI211_X1 g138(.A(new_n560), .B(new_n562), .C1(new_n563), .C2(new_n548), .ZN(G301));
  INV_X1    g139(.A(G301), .ZN(G171));
  NAND2_X1  g140(.A1(new_n559), .A2(G43), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n536), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n538), .ZN(new_n568));
  INV_X1    g143(.A(G81), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n566), .B(new_n568), .C1(new_n569), .C2(new_n548), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G860), .ZN(G153));
  AND3_X1   g147(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G36), .ZN(G176));
  NAND2_X1  g149(.A1(G1), .A2(G3), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT8), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n573), .A2(new_n576), .ZN(G188));
  AOI21_X1  g152(.A(KEYINPUT76), .B1(new_n559), .B2(G53), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n548), .ZN(new_n581));
  NAND2_X1  g156(.A1(G78), .A2(G543), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n533), .A2(new_n535), .ZN(new_n583));
  INV_X1    g158(.A(G65), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n581), .A2(G91), .B1(G651), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n580), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n559), .A2(KEYINPUT76), .A3(G53), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(KEYINPUT9), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(new_n578), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n588), .A2(new_n591), .ZN(G299));
  INV_X1    g167(.A(G166), .ZN(G303));
  NAND2_X1  g168(.A1(new_n559), .A2(G49), .ZN(new_n594));
  INV_X1    g169(.A(G74), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n538), .B1(new_n583), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT77), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n581), .A2(G87), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n594), .A2(new_n597), .A3(new_n598), .ZN(G288));
  NAND2_X1  g174(.A1(G73), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G61), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n583), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G651), .ZN(new_n603));
  NAND2_X1  g178(.A1(G48), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G86), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n583), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(new_n547), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(G305));
  NAND2_X1  g183(.A1(new_n559), .A2(G47), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n536), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n610), .A2(new_n538), .ZN(new_n611));
  INV_X1    g186(.A(G85), .ZN(new_n612));
  OAI211_X1 g187(.A(new_n609), .B(new_n611), .C1(new_n612), .C2(new_n548), .ZN(G290));
  NAND2_X1  g188(.A1(G301), .A2(G868), .ZN(new_n614));
  INV_X1    g189(.A(G54), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n536), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n616));
  OAI22_X1  g191(.A1(new_n556), .A2(new_n615), .B1(new_n538), .B2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n581), .A2(G92), .ZN(new_n620));
  XOR2_X1   g195(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT80), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n614), .B1(new_n625), .B2(G868), .ZN(G284));
  OAI21_X1  g201(.A(new_n614), .B1(new_n625), .B2(G868), .ZN(G321));
  NAND2_X1  g202(.A1(G286), .A2(G868), .ZN(new_n628));
  XOR2_X1   g203(.A(G299), .B(KEYINPUT81), .Z(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G868), .ZN(G280));
  XNOR2_X1  g205(.A(G280), .B(KEYINPUT82), .ZN(G297));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n625), .B1(new_n632), .B2(G860), .ZN(G148));
  INV_X1    g208(.A(G868), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n570), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n624), .A2(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(new_n634), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT83), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n496), .A2(new_n499), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(new_n514), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT13), .ZN(new_n644));
  INV_X1    g219(.A(G2100), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n509), .A2(G123), .ZN(new_n647));
  INV_X1    g222(.A(new_n505), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(G135), .ZN(new_n649));
  OAI221_X1 g224(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n475), .C2(G111), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n647), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(G2096), .Z(new_n652));
  NAND2_X1  g227(.A1(new_n646), .A2(new_n652), .ZN(G156));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT85), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2427), .B(G2430), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT14), .ZN(new_n659));
  XOR2_X1   g234(.A(G2451), .B(G2454), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n665), .B(new_n666), .Z(new_n667));
  AND2_X1   g242(.A1(new_n667), .A2(G14), .ZN(G401));
  XOR2_X1   g243(.A(G2067), .B(G2678), .Z(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT87), .Z(new_n670));
  XOR2_X1   g245(.A(G2072), .B(G2078), .Z(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n670), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT18), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n671), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n671), .B(KEYINPUT17), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n676), .B(new_n673), .C1(new_n670), .C2(new_n677), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n670), .A2(new_n677), .A3(new_n672), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G2096), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(new_n645), .ZN(G227));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n683), .A2(new_n684), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT20), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n689), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n686), .A2(new_n688), .A3(new_n690), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n693), .B(new_n694), .C1(new_n692), .C2(new_n691), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT21), .B(G1986), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(G1991), .B(G1996), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT22), .B(G1981), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n699), .B(new_n700), .Z(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(G229));
  OAI21_X1  g277(.A(KEYINPUT92), .B1(G16), .B2(G23), .ZN(new_n703));
  OR3_X1    g278(.A1(KEYINPUT92), .A2(G16), .A3(G23), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n703), .B(new_n704), .C1(G288), .C2(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT33), .B(G1976), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n705), .A2(G22), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G166), .B2(new_n705), .ZN(new_n710));
  INV_X1    g285(.A(G1971), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n705), .A2(G6), .ZN(new_n713));
  INV_X1    g288(.A(G305), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n705), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT32), .B(G1981), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n708), .A2(new_n712), .A3(new_n717), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT91), .Z(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(KEYINPUT34), .ZN(new_n720));
  NAND2_X1  g295(.A1(G290), .A2(G16), .ZN(new_n721));
  INV_X1    g296(.A(G24), .ZN(new_n722));
  OAI21_X1  g297(.A(KEYINPUT90), .B1(new_n722), .B2(G16), .ZN(new_n723));
  OR3_X1    g298(.A1(new_n722), .A2(KEYINPUT90), .A3(G16), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n721), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(G1986), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n719), .A2(KEYINPUT34), .ZN(new_n727));
  NOR2_X1   g302(.A1(G25), .A2(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n648), .A2(G131), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n509), .A2(G119), .ZN(new_n730));
  NOR2_X1   g305(.A1(G95), .A2(G2105), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT88), .Z(new_n732));
  OAI211_X1 g307(.A(new_n732), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n729), .A2(new_n730), .A3(new_n733), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT89), .Z(new_n735));
  AOI21_X1  g310(.A(new_n728), .B1(new_n735), .B2(G29), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT35), .B(G1991), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n720), .A2(new_n726), .A3(new_n727), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT36), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n705), .A2(G21), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G168), .B2(new_n705), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1966), .ZN(new_n743));
  NOR2_X1   g318(.A1(G5), .A2(G16), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G171), .B2(G16), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n743), .B1(G1961), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(G29), .A2(G32), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n648), .A2(G141), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n509), .A2(G129), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n514), .A2(G105), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT26), .Z(new_n752));
  NAND4_X1  g327(.A1(new_n748), .A2(new_n749), .A3(new_n750), .A4(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n747), .B1(new_n754), .B2(G29), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT27), .B(G1996), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G2078), .ZN(new_n758));
  NAND2_X1  g333(.A1(G164), .A2(G29), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G27), .B2(G29), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n757), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n760), .A2(new_n758), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT30), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G28), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT96), .ZN(new_n765));
  INV_X1    g340(.A(G29), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n765), .B(new_n766), .C1(new_n763), .C2(G28), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n746), .A2(new_n761), .A3(new_n762), .A4(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n651), .A2(new_n766), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT31), .B(G11), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n766), .A2(G33), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT25), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n648), .A2(G139), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n640), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n774), .B(new_n775), .C1(new_n475), .C2(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT94), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n771), .B1(new_n778), .B2(new_n766), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G2072), .ZN(new_n780));
  NOR4_X1   g355(.A1(new_n768), .A2(new_n769), .A3(new_n770), .A4(new_n780), .ZN(new_n781));
  AND2_X1   g356(.A1(KEYINPUT24), .A2(G34), .ZN(new_n782));
  NOR2_X1   g357(.A1(KEYINPUT24), .A2(G34), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n782), .A2(new_n783), .A3(G29), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n503), .B2(G29), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT95), .B(G2084), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n781), .B(new_n787), .C1(G1961), .C2(new_n745), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT97), .ZN(new_n789));
  OAI21_X1  g364(.A(KEYINPUT93), .B1(G4), .B2(G16), .ZN(new_n790));
  OR3_X1    g365(.A1(KEYINPUT93), .A2(G4), .A3(G16), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n790), .B(new_n791), .C1(new_n624), .C2(new_n705), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(G1348), .Z(new_n793));
  AND3_X1   g368(.A1(new_n705), .A2(KEYINPUT23), .A3(G20), .ZN(new_n794));
  AOI21_X1  g369(.A(KEYINPUT23), .B1(new_n705), .B2(G20), .ZN(new_n795));
  AOI211_X1 g370(.A(new_n794), .B(new_n795), .C1(G299), .C2(G16), .ZN(new_n796));
  INV_X1    g371(.A(G1956), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n740), .A2(new_n789), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT28), .ZN(new_n801));
  INV_X1    g376(.A(G26), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(G29), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(G29), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n509), .A2(G128), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n648), .A2(G140), .ZN(new_n806));
  OAI221_X1 g381(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n475), .C2(G116), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n804), .B1(new_n808), .B2(G29), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n803), .B1(new_n809), .B2(new_n801), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G2067), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n766), .A2(G35), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G162), .B2(new_n766), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT29), .B(G2090), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n705), .A2(G19), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n571), .B2(new_n705), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(G1341), .Z(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  NOR4_X1   g394(.A1(new_n800), .A2(new_n811), .A3(new_n815), .A4(new_n819), .ZN(G311));
  INV_X1    g395(.A(new_n800), .ZN(new_n821));
  INV_X1    g396(.A(new_n811), .ZN(new_n822));
  INV_X1    g397(.A(new_n815), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n821), .A2(new_n822), .A3(new_n823), .A4(new_n818), .ZN(G150));
  AOI22_X1  g399(.A1(new_n536), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT99), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n826), .A2(new_n538), .ZN(new_n827));
  INV_X1    g402(.A(G55), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT100), .B(G93), .ZN(new_n829));
  OAI22_X1  g404(.A1(new_n556), .A2(new_n828), .B1(new_n548), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G860), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT37), .Z(new_n834));
  NOR2_X1   g409(.A1(new_n624), .A2(new_n632), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT39), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n831), .B(new_n570), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n834), .B1(new_n840), .B2(G860), .ZN(G145));
  INV_X1    g416(.A(KEYINPUT104), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n778), .B(new_n808), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n843), .A2(new_n754), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n754), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(KEYINPUT4), .B1(new_n640), .B2(new_n520), .ZN(new_n847));
  OAI211_X1 g422(.A(KEYINPUT4), .B(new_n466), .C1(new_n468), .C2(new_n469), .ZN(new_n848));
  INV_X1    g423(.A(new_n520), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n515), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(KEYINPUT101), .B1(new_n851), .B2(new_n525), .ZN(new_n852));
  AND4_X1   g427(.A1(KEYINPUT101), .A2(new_n521), .A3(new_n525), .A4(new_n529), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n846), .A2(new_n855), .ZN(new_n856));
  OAI221_X1 g431(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n475), .C2(G118), .ZN(new_n857));
  INV_X1    g432(.A(G142), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n857), .B1(new_n505), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(G130), .B2(new_n509), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n734), .ZN(new_n861));
  XOR2_X1   g436(.A(KEYINPUT102), .B(KEYINPUT103), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(new_n643), .Z(new_n864));
  NAND3_X1  g439(.A1(new_n844), .A2(new_n854), .A3(new_n845), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n856), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n864), .B1(new_n856), .B2(new_n865), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n842), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n867), .A2(new_n842), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n503), .B(new_n512), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n651), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n868), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT105), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n866), .A2(new_n867), .ZN(new_n875));
  AOI21_X1  g450(.A(G37), .B1(new_n875), .B2(new_n871), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT105), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n868), .A2(new_n869), .A3(new_n877), .A4(new_n872), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n874), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(KEYINPUT40), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT40), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n874), .A2(new_n876), .A3(new_n881), .A4(new_n878), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(G395));
  NAND2_X1  g458(.A1(new_n832), .A2(new_n634), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n636), .B(new_n839), .Z(new_n885));
  NAND3_X1  g460(.A1(new_n588), .A2(new_n591), .A3(KEYINPUT106), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT106), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n590), .A2(new_n578), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n887), .B1(new_n888), .B2(new_n587), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n619), .A2(new_n622), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n886), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(G299), .A2(new_n887), .A3(new_n623), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT108), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT41), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(KEYINPUT41), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n891), .A2(new_n897), .A3(new_n892), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(KEYINPUT108), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n885), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n900), .A2(KEYINPUT109), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(KEYINPUT109), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n893), .B(KEYINPUT107), .Z(new_n903));
  OAI211_X1 g478(.A(new_n901), .B(new_n902), .C1(new_n903), .C2(new_n885), .ZN(new_n904));
  XNOR2_X1  g479(.A(G290), .B(G166), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(G288), .ZN(new_n906));
  XOR2_X1   g481(.A(G305), .B(KEYINPUT110), .Z(new_n907));
  XOR2_X1   g482(.A(new_n906), .B(new_n907), .Z(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT42), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n904), .B(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n884), .B1(new_n910), .B2(new_n634), .ZN(G295));
  OAI21_X1  g486(.A(new_n884), .B1(new_n910), .B2(new_n634), .ZN(G331));
  INV_X1    g487(.A(KEYINPUT111), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n899), .A2(new_n895), .ZN(new_n915));
  XNOR2_X1  g490(.A(G168), .B(G301), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n839), .B(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n908), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n917), .B1(new_n892), .B2(new_n891), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n917), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(new_n899), .B2(new_n895), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n908), .B1(new_n924), .B2(new_n920), .ZN(new_n925));
  INV_X1    g500(.A(G37), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n922), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n903), .A2(new_n923), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n917), .A2(new_n896), .A3(new_n898), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n919), .A3(new_n931), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n932), .A2(new_n925), .A3(KEYINPUT43), .A4(new_n926), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n914), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n927), .A2(KEYINPUT43), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n932), .A2(new_n925), .A3(new_n928), .A4(new_n926), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n914), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n913), .B1(new_n935), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT44), .B1(new_n936), .B2(new_n937), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n934), .A2(new_n941), .A3(KEYINPUT111), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n940), .A2(new_n942), .ZN(G397));
  NAND2_X1  g518(.A1(G286), .A2(G8), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n490), .A2(KEYINPUT73), .ZN(new_n945));
  AOI211_X1 g520(.A(new_n480), .B(new_n482), .C1(new_n487), .C2(new_n489), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n502), .B(G40), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n492), .A2(KEYINPUT112), .A3(G40), .A4(new_n502), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT50), .ZN(new_n951));
  INV_X1    g526(.A(G1384), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n530), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n949), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT113), .ZN(new_n955));
  AOI21_X1  g530(.A(G1384), .B1(new_n851), .B2(new_n525), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n955), .B1(new_n956), .B2(new_n951), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n530), .A2(new_n952), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n958), .A2(KEYINPUT113), .A3(KEYINPUT50), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n954), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G2084), .ZN(new_n961));
  INV_X1    g536(.A(G1966), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n958), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n530), .A2(KEYINPUT45), .A3(new_n952), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n964), .A2(new_n949), .A3(new_n950), .A4(new_n965), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n960), .A2(new_n961), .B1(new_n962), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G8), .ZN(new_n968));
  OAI211_X1 g543(.A(KEYINPUT51), .B(new_n944), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n957), .A2(new_n959), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n949), .A2(new_n950), .A3(new_n953), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n961), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n966), .A2(new_n962), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n970), .B(G8), .C1(new_n975), .C2(G286), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n969), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT121), .ZN(new_n978));
  INV_X1    g553(.A(new_n944), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n978), .B1(new_n975), .B2(new_n979), .ZN(new_n980));
  AOI211_X1 g555(.A(KEYINPUT121), .B(new_n944), .C1(new_n973), .C2(new_n974), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT122), .B1(new_n977), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT62), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT121), .B1(new_n967), .B2(new_n944), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n975), .A2(new_n978), .A3(new_n979), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT122), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n987), .A2(new_n988), .A3(new_n976), .A4(new_n969), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n983), .A2(new_n984), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n991));
  NAND3_X1  g566(.A1(G303), .A2(new_n991), .A3(G8), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT55), .B1(G166), .B2(new_n968), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n949), .A2(new_n950), .ZN(new_n995));
  OAI211_X1 g570(.A(KEYINPUT45), .B(new_n952), .C1(new_n852), .C2(new_n853), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n995), .A2(new_n964), .A3(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n956), .A2(new_n951), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n954), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G2090), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n997), .A2(new_n711), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n994), .B1(new_n1001), .B2(new_n968), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n994), .A2(KEYINPUT114), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT114), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n992), .A2(new_n1004), .A3(new_n993), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT113), .B1(new_n958), .B2(KEYINPUT50), .ZN(new_n1008));
  AOI211_X1 g583(.A(new_n955), .B(new_n951), .C1(new_n530), .C2(new_n952), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n1010), .A2(G2090), .A3(new_n954), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n964), .A2(new_n949), .A3(new_n950), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1971), .B1(new_n1012), .B2(new_n996), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1007), .B(G8), .C1(new_n1011), .C2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n949), .A2(new_n950), .A3(new_n956), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1015), .A2(G8), .ZN(new_n1016));
  XNOR2_X1  g591(.A(G305), .B(G1981), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT49), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1976), .ZN(new_n1020));
  OR2_X1    g595(.A1(G288), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1015), .A2(G8), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT52), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT52), .B1(G288), .B2(new_n1020), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1015), .A2(G8), .A3(new_n1021), .A4(new_n1024), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1019), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1002), .A2(new_n1014), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n995), .A2(new_n996), .A3(new_n758), .A4(new_n964), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n971), .A2(new_n972), .ZN(new_n1030));
  INV_X1    g605(.A(G1961), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n1028), .A2(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1028), .A2(G2078), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1012), .A2(new_n965), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(G171), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1027), .A2(new_n1036), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n990), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT125), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n983), .A2(new_n989), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1039), .B1(new_n1040), .B2(KEYINPUT62), .ZN(new_n1041));
  AOI211_X1 g616(.A(KEYINPUT125), .B(new_n984), .C1(new_n983), .C2(new_n989), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1038), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT126), .ZN(new_n1044));
  INV_X1    g619(.A(G1996), .ZN(new_n1045));
  AND4_X1   g620(.A1(new_n1045), .A2(new_n995), .A3(new_n964), .A4(new_n996), .ZN(new_n1046));
  XOR2_X1   g621(.A(KEYINPUT58), .B(G1341), .Z(new_n1047));
  AND2_X1   g622(.A1(new_n1015), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n571), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT59), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1051), .B(new_n571), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1052));
  AOI21_X1  g627(.A(G1348), .B1(new_n971), .B2(new_n972), .ZN(new_n1053));
  INV_X1    g628(.A(G2067), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n949), .A2(new_n950), .A3(new_n1054), .A4(new_n956), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1059));
  NOR4_X1   g634(.A1(new_n1053), .A2(new_n1058), .A3(new_n1059), .A4(KEYINPUT60), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1050), .A2(new_n1052), .B1(new_n1060), .B2(new_n890), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1053), .A2(new_n1059), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n623), .B1(new_n1062), .B2(new_n1057), .ZN(new_n1063));
  NOR4_X1   g638(.A1(new_n1053), .A2(new_n1058), .A3(new_n1059), .A4(new_n890), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT60), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n588), .A2(new_n591), .A3(KEYINPUT57), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n888), .B2(new_n587), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n797), .B1(new_n954), .B2(new_n998), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT56), .B(G2072), .Z(new_n1071));
  OAI211_X1 g646(.A(new_n1069), .B(new_n1070), .C1(new_n997), .C2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT61), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1072), .B(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1061), .A2(new_n1065), .A3(new_n1074), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n997), .A2(new_n1071), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1069), .B1(new_n1076), .B2(new_n1070), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1072), .ZN(new_n1078));
  OAI22_X1  g653(.A1(new_n960), .A2(G1348), .B1(new_n1056), .B2(new_n1055), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n890), .B1(new_n1079), .B2(new_n1058), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1078), .B1(new_n1080), .B2(KEYINPUT119), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1063), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1077), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1075), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1085), .B1(new_n1075), .B2(new_n1084), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1029), .A2(new_n1028), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT123), .ZN(new_n1090));
  INV_X1    g665(.A(new_n947), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT101), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n530), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n851), .A2(KEYINPUT101), .A3(new_n525), .ZN(new_n1094));
  AOI21_X1  g669(.A(G1384), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1091), .B1(new_n1095), .B2(KEYINPUT45), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n996), .A2(new_n1033), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1090), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n952), .B1(new_n852), .B2(new_n853), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n947), .B1(new_n1099), .B2(new_n963), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1033), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1101), .B1(new_n1095), .B2(KEYINPUT45), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1100), .A2(new_n1102), .A3(KEYINPUT123), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1031), .B1(new_n1010), .B2(new_n954), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1089), .A2(new_n1098), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(G171), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1032), .A2(G301), .A3(new_n1034), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(KEYINPUT54), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT124), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT124), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1106), .A2(new_n1110), .A3(KEYINPUT54), .A4(new_n1107), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1027), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1032), .A2(G301), .A3(new_n1098), .A4(new_n1103), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT54), .B1(new_n1036), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(new_n983), .B2(new_n989), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  AOI211_X1 g691(.A(new_n968), .B(G286), .C1(new_n973), .C2(new_n974), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1002), .A2(new_n1014), .A3(new_n1026), .A4(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT116), .B(KEYINPUT63), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT63), .ZN(new_n1121));
  OAI21_X1  g696(.A(G8), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1121), .B1(new_n1122), .B2(new_n994), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1123), .A2(new_n1014), .A3(new_n1026), .A4(new_n1117), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1014), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n1026), .ZN(new_n1127));
  NOR2_X1   g702(.A1(G288), .A2(G1976), .ZN(new_n1128));
  XOR2_X1   g703(.A(new_n1128), .B(KEYINPUT115), .Z(new_n1129));
  OAI22_X1  g704(.A1(new_n1129), .A2(new_n1018), .B1(G1981), .B2(G305), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n1016), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1125), .A2(new_n1127), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(KEYINPUT117), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT117), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1125), .A2(new_n1134), .A3(new_n1127), .A4(new_n1131), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1088), .A2(new_n1116), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1038), .B(new_n1137), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1044), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1095), .A2(KEYINPUT45), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n995), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n753), .B(new_n1045), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n808), .B(new_n1054), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n734), .B(new_n737), .Z(new_n1146));
  OAI21_X1  g721(.A(new_n1142), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(G290), .B(G1986), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1148), .B1(new_n1142), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1139), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1152), .A2(new_n737), .A3(new_n735), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n808), .A2(G2067), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1141), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1142), .A2(KEYINPUT46), .A3(new_n1045), .ZN(new_n1156));
  AOI21_X1  g731(.A(KEYINPUT46), .B1(new_n1142), .B2(new_n1045), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1141), .B1(new_n754), .B2(new_n1144), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT47), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1141), .A2(G1986), .A3(G290), .ZN(new_n1161));
  XNOR2_X1  g736(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1161), .B(new_n1162), .ZN(new_n1163));
  AOI211_X1 g738(.A(new_n1155), .B(new_n1160), .C1(new_n1147), .C2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1151), .A2(new_n1164), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g740(.A1(G401), .A2(G227), .ZN(new_n1167));
  AOI21_X1  g741(.A(new_n463), .B1(new_n936), .B2(new_n937), .ZN(new_n1168));
  NAND4_X1  g742(.A1(new_n879), .A2(new_n701), .A3(new_n1167), .A4(new_n1168), .ZN(G225));
  INV_X1    g743(.A(G225), .ZN(G308));
endmodule


