

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580;

  XNOR2_X1 U321 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U322 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U323 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U324 ( .A(KEYINPUT54), .B(n410), .Z(n289) );
  XNOR2_X1 U325 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n342) );
  XNOR2_X1 U326 ( .A(n343), .B(n342), .ZN(n383) );
  XNOR2_X1 U327 ( .A(n351), .B(KEYINPUT33), .ZN(n352) );
  XNOR2_X1 U328 ( .A(KEYINPUT97), .B(KEYINPUT36), .ZN(n322) );
  XNOR2_X1 U329 ( .A(n353), .B(n352), .ZN(n356) );
  XNOR2_X1 U330 ( .A(n388), .B(n322), .ZN(n577) );
  XNOR2_X1 U331 ( .A(n364), .B(n363), .ZN(n569) );
  NOR2_X1 U332 ( .A1(n524), .A2(n448), .ZN(n558) );
  XOR2_X1 U333 ( .A(n307), .B(n306), .Z(n515) );
  XNOR2_X1 U334 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U335 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XOR2_X1 U336 ( .A(G120GAT), .B(G71GAT), .Z(n360) );
  XOR2_X1 U337 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n291) );
  XNOR2_X1 U338 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n290) );
  XNOR2_X1 U339 ( .A(n291), .B(n290), .ZN(n406) );
  XOR2_X1 U340 ( .A(n360), .B(n406), .Z(n293) );
  XNOR2_X1 U341 ( .A(G43GAT), .B(G190GAT), .ZN(n292) );
  XNOR2_X1 U342 ( .A(n293), .B(n292), .ZN(n299) );
  XOR2_X1 U343 ( .A(G127GAT), .B(KEYINPUT0), .Z(n295) );
  XNOR2_X1 U344 ( .A(G113GAT), .B(G134GAT), .ZN(n294) );
  XNOR2_X1 U345 ( .A(n295), .B(n294), .ZN(n428) );
  XOR2_X1 U346 ( .A(n428), .B(G176GAT), .Z(n297) );
  NAND2_X1 U347 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U349 ( .A(n299), .B(n298), .Z(n307) );
  XOR2_X1 U350 ( .A(KEYINPUT80), .B(KEYINPUT82), .Z(n301) );
  XNOR2_X1 U351 ( .A(G99GAT), .B(KEYINPUT83), .ZN(n300) );
  XNOR2_X1 U352 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U353 ( .A(G183GAT), .B(KEYINPUT20), .Z(n303) );
  XNOR2_X1 U354 ( .A(G15GAT), .B(KEYINPUT81), .ZN(n302) );
  XNOR2_X1 U355 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U356 ( .A(n305), .B(n304), .ZN(n306) );
  INV_X1 U357 ( .A(n515), .ZN(n524) );
  XOR2_X1 U358 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n309) );
  XNOR2_X1 U359 ( .A(G218GAT), .B(KEYINPUT75), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n309), .B(n308), .ZN(n321) );
  XOR2_X1 U361 ( .A(G29GAT), .B(G43GAT), .Z(n311) );
  XNOR2_X1 U362 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n376) );
  XOR2_X1 U364 ( .A(G36GAT), .B(G190GAT), .Z(n399) );
  XNOR2_X1 U365 ( .A(n376), .B(n399), .ZN(n313) );
  AND2_X1 U366 ( .A1(G232GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U367 ( .A(n313), .B(n312), .ZN(n319) );
  XOR2_X1 U368 ( .A(G50GAT), .B(G162GAT), .Z(n431) );
  XOR2_X1 U369 ( .A(G99GAT), .B(G85GAT), .Z(n346) );
  XNOR2_X1 U370 ( .A(n431), .B(n346), .ZN(n317) );
  XOR2_X1 U371 ( .A(KEYINPUT11), .B(G92GAT), .Z(n315) );
  XNOR2_X1 U372 ( .A(G134GAT), .B(G106GAT), .ZN(n314) );
  XOR2_X1 U373 ( .A(n315), .B(n314), .Z(n316) );
  XOR2_X1 U374 ( .A(n321), .B(n320), .Z(n388) );
  XOR2_X1 U375 ( .A(G211GAT), .B(G155GAT), .Z(n324) );
  XNOR2_X1 U376 ( .A(G127GAT), .B(G71GAT), .ZN(n323) );
  XNOR2_X1 U377 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U378 ( .A(G57GAT), .B(KEYINPUT13), .Z(n359) );
  XOR2_X1 U379 ( .A(n325), .B(n359), .Z(n327) );
  XNOR2_X1 U380 ( .A(G22GAT), .B(G78GAT), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n333) );
  XOR2_X1 U382 ( .A(G8GAT), .B(G183GAT), .Z(n398) );
  XOR2_X1 U383 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n329) );
  XNOR2_X1 U384 ( .A(G15GAT), .B(G1GAT), .ZN(n328) );
  XNOR2_X1 U385 ( .A(n329), .B(n328), .ZN(n377) );
  XOR2_X1 U386 ( .A(n398), .B(n377), .Z(n331) );
  NAND2_X1 U387 ( .A1(G231GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U388 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U389 ( .A(n333), .B(n332), .Z(n341) );
  XOR2_X1 U390 ( .A(KEYINPUT14), .B(KEYINPUT79), .Z(n335) );
  XNOR2_X1 U391 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U393 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n337) );
  XNOR2_X1 U394 ( .A(KEYINPUT15), .B(KEYINPUT76), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U397 ( .A(n341), .B(n340), .Z(n573) );
  INV_X1 U398 ( .A(n573), .ZN(n479) );
  NOR2_X1 U399 ( .A1(n577), .A2(n479), .ZN(n343) );
  XNOR2_X1 U400 ( .A(G64GAT), .B(G92GAT), .ZN(n345) );
  XNOR2_X1 U401 ( .A(G176GAT), .B(G204GAT), .ZN(n344) );
  XNOR2_X1 U402 ( .A(n345), .B(n344), .ZN(n347) );
  INV_X1 U403 ( .A(n347), .ZN(n403) );
  NAND2_X1 U404 ( .A1(n346), .A2(n403), .ZN(n350) );
  INV_X1 U405 ( .A(n346), .ZN(n348) );
  NAND2_X1 U406 ( .A1(n348), .A2(n347), .ZN(n349) );
  NAND2_X1 U407 ( .A1(n350), .A2(n349), .ZN(n353) );
  AND2_X1 U408 ( .A1(G230GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U409 ( .A(G106GAT), .B(G78GAT), .ZN(n354) );
  XNOR2_X1 U410 ( .A(n354), .B(G148GAT), .ZN(n432) );
  XOR2_X1 U411 ( .A(n432), .B(KEYINPUT74), .Z(n355) );
  XNOR2_X1 U412 ( .A(n356), .B(n355), .ZN(n364) );
  XOR2_X1 U413 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n358) );
  XNOR2_X1 U414 ( .A(KEYINPUT73), .B(KEYINPUT72), .ZN(n357) );
  XOR2_X1 U415 ( .A(n358), .B(n357), .Z(n362) );
  XNOR2_X1 U416 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U417 ( .A(G141GAT), .B(G22GAT), .Z(n436) );
  XOR2_X1 U418 ( .A(G113GAT), .B(G197GAT), .Z(n366) );
  XNOR2_X1 U419 ( .A(G36GAT), .B(G50GAT), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U421 ( .A(n436), .B(n367), .Z(n369) );
  NAND2_X1 U422 ( .A1(G229GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U423 ( .A(n369), .B(n368), .ZN(n381) );
  XOR2_X1 U424 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n371) );
  XNOR2_X1 U425 ( .A(KEYINPUT68), .B(KEYINPUT66), .ZN(n370) );
  XNOR2_X1 U426 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U427 ( .A(KEYINPUT69), .B(KEYINPUT67), .Z(n373) );
  XNOR2_X1 U428 ( .A(G169GAT), .B(G8GAT), .ZN(n372) );
  XNOR2_X1 U429 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U430 ( .A(n375), .B(n374), .Z(n379) );
  XNOR2_X1 U431 ( .A(n376), .B(n377), .ZN(n378) );
  XNOR2_X1 U432 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U433 ( .A(n381), .B(n380), .Z(n494) );
  AND2_X1 U434 ( .A1(n569), .A2(n494), .ZN(n382) );
  AND2_X1 U435 ( .A1(n383), .A2(n382), .ZN(n384) );
  XNOR2_X1 U436 ( .A(n384), .B(KEYINPUT110), .ZN(n393) );
  INV_X1 U437 ( .A(n494), .ZN(n563) );
  XNOR2_X1 U438 ( .A(KEYINPUT41), .B(n569), .ZN(n555) );
  NAND2_X1 U439 ( .A1(n563), .A2(n555), .ZN(n385) );
  XNOR2_X1 U440 ( .A(KEYINPUT46), .B(n385), .ZN(n386) );
  NAND2_X1 U441 ( .A1(n386), .A2(n479), .ZN(n387) );
  XNOR2_X1 U442 ( .A(KEYINPUT108), .B(n387), .ZN(n389) );
  NOR2_X1 U443 ( .A1(n389), .A2(n388), .ZN(n391) );
  XNOR2_X1 U444 ( .A(KEYINPUT47), .B(KEYINPUT109), .ZN(n390) );
  XNOR2_X1 U445 ( .A(n391), .B(n390), .ZN(n392) );
  NOR2_X1 U446 ( .A1(n393), .A2(n392), .ZN(n394) );
  XNOR2_X1 U447 ( .A(n394), .B(KEYINPUT48), .ZN(n521) );
  XOR2_X1 U448 ( .A(KEYINPUT90), .B(KEYINPUT92), .Z(n396) );
  NAND2_X1 U449 ( .A1(G226GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U450 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U451 ( .A(n397), .B(KEYINPUT91), .Z(n401) );
  XNOR2_X1 U452 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U453 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U454 ( .A(n403), .B(n402), .Z(n408) );
  XOR2_X1 U455 ( .A(G211GAT), .B(KEYINPUT21), .Z(n405) );
  XNOR2_X1 U456 ( .A(G197GAT), .B(G218GAT), .ZN(n404) );
  XNOR2_X1 U457 ( .A(n405), .B(n404), .ZN(n443) );
  XNOR2_X1 U458 ( .A(n406), .B(n443), .ZN(n407) );
  XOR2_X1 U459 ( .A(n408), .B(n407), .Z(n512) );
  INV_X1 U460 ( .A(n512), .ZN(n409) );
  NOR2_X1 U461 ( .A1(n521), .A2(n409), .ZN(n410) );
  XOR2_X1 U462 ( .A(G85GAT), .B(G148GAT), .Z(n412) );
  XNOR2_X1 U463 ( .A(G29GAT), .B(G162GAT), .ZN(n411) );
  XNOR2_X1 U464 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U465 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n414) );
  XNOR2_X1 U466 ( .A(G141GAT), .B(G120GAT), .ZN(n413) );
  XNOR2_X1 U467 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U468 ( .A(n416), .B(n415), .Z(n421) );
  XOR2_X1 U469 ( .A(KEYINPUT87), .B(KEYINPUT4), .Z(n418) );
  NAND2_X1 U470 ( .A1(G225GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U471 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U472 ( .A(KEYINPUT5), .B(n419), .ZN(n420) );
  XNOR2_X1 U473 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U474 ( .A(G57GAT), .B(KEYINPUT1), .Z(n423) );
  XNOR2_X1 U475 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n422) );
  XNOR2_X1 U476 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U477 ( .A(n425), .B(n424), .Z(n430) );
  XOR2_X1 U478 ( .A(G155GAT), .B(KEYINPUT2), .Z(n427) );
  XNOR2_X1 U479 ( .A(KEYINPUT86), .B(KEYINPUT3), .ZN(n426) );
  XNOR2_X1 U480 ( .A(n427), .B(n426), .ZN(n444) );
  XNOR2_X1 U481 ( .A(n428), .B(n444), .ZN(n429) );
  XNOR2_X1 U482 ( .A(n430), .B(n429), .ZN(n510) );
  NOR2_X1 U483 ( .A1(n289), .A2(n510), .ZN(n560) );
  XOR2_X1 U484 ( .A(n432), .B(n431), .Z(n434) );
  NAND2_X1 U485 ( .A1(G228GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U486 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U487 ( .A(n435), .B(G204GAT), .Z(n438) );
  XNOR2_X1 U488 ( .A(n436), .B(KEYINPUT23), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U490 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n440) );
  XNOR2_X1 U491 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U493 ( .A(n442), .B(n441), .Z(n446) );
  XNOR2_X1 U494 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U495 ( .A(n446), .B(n445), .ZN(n462) );
  NAND2_X1 U496 ( .A1(n560), .A2(n462), .ZN(n447) );
  XOR2_X1 U497 ( .A(KEYINPUT55), .B(n447), .Z(n448) );
  NAND2_X1 U498 ( .A1(n558), .A2(n388), .ZN(n452) );
  XOR2_X1 U499 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n450) );
  XNOR2_X1 U500 ( .A(G190GAT), .B(KEYINPUT121), .ZN(n449) );
  XOR2_X1 U501 ( .A(KEYINPUT34), .B(KEYINPUT96), .Z(n471) );
  NAND2_X1 U502 ( .A1(n569), .A2(n563), .ZN(n482) );
  NOR2_X1 U503 ( .A1(n388), .A2(n479), .ZN(n453) );
  XNOR2_X1 U504 ( .A(n453), .B(KEYINPUT16), .ZN(n468) );
  XNOR2_X1 U505 ( .A(n512), .B(KEYINPUT27), .ZN(n464) );
  NOR2_X1 U506 ( .A1(n515), .A2(n462), .ZN(n454) );
  XOR2_X1 U507 ( .A(n454), .B(KEYINPUT26), .Z(n539) );
  INV_X1 U508 ( .A(n539), .ZN(n561) );
  NAND2_X1 U509 ( .A1(n464), .A2(n561), .ZN(n455) );
  XNOR2_X1 U510 ( .A(KEYINPUT93), .B(n455), .ZN(n459) );
  NAND2_X1 U511 ( .A1(n515), .A2(n512), .ZN(n456) );
  NAND2_X1 U512 ( .A1(n462), .A2(n456), .ZN(n457) );
  XNOR2_X1 U513 ( .A(KEYINPUT25), .B(n457), .ZN(n458) );
  NOR2_X1 U514 ( .A1(n459), .A2(n458), .ZN(n460) );
  NOR2_X1 U515 ( .A1(n510), .A2(n460), .ZN(n461) );
  XOR2_X1 U516 ( .A(KEYINPUT94), .B(n461), .Z(n467) );
  XNOR2_X1 U517 ( .A(n462), .B(KEYINPUT65), .ZN(n463) );
  XNOR2_X1 U518 ( .A(n463), .B(KEYINPUT28), .ZN(n527) );
  NAND2_X1 U519 ( .A1(n510), .A2(n464), .ZN(n522) );
  NOR2_X1 U520 ( .A1(n527), .A2(n522), .ZN(n465) );
  NAND2_X1 U521 ( .A1(n524), .A2(n465), .ZN(n466) );
  NAND2_X1 U522 ( .A1(n467), .A2(n466), .ZN(n478) );
  NAND2_X1 U523 ( .A1(n468), .A2(n478), .ZN(n469) );
  XOR2_X1 U524 ( .A(KEYINPUT95), .B(n469), .Z(n496) );
  NOR2_X1 U525 ( .A1(n482), .A2(n496), .ZN(n476) );
  NAND2_X1 U526 ( .A1(n476), .A2(n510), .ZN(n470) );
  XNOR2_X1 U527 ( .A(n471), .B(n470), .ZN(n472) );
  XOR2_X1 U528 ( .A(G1GAT), .B(n472), .Z(G1324GAT) );
  NAND2_X1 U529 ( .A1(n512), .A2(n476), .ZN(n473) );
  XNOR2_X1 U530 ( .A(n473), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U531 ( .A(G15GAT), .B(KEYINPUT35), .Z(n475) );
  NAND2_X1 U532 ( .A1(n476), .A2(n515), .ZN(n474) );
  XNOR2_X1 U533 ( .A(n475), .B(n474), .ZN(G1326GAT) );
  NAND2_X1 U534 ( .A1(n476), .A2(n527), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n477), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U536 ( .A(G29GAT), .B(KEYINPUT39), .Z(n486) );
  NAND2_X1 U537 ( .A1(n479), .A2(n478), .ZN(n480) );
  NOR2_X1 U538 ( .A1(n577), .A2(n480), .ZN(n481) );
  XNOR2_X1 U539 ( .A(KEYINPUT37), .B(n481), .ZN(n508) );
  NOR2_X1 U540 ( .A1(n508), .A2(n482), .ZN(n484) );
  XNOR2_X1 U541 ( .A(KEYINPUT98), .B(KEYINPUT38), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n484), .B(n483), .ZN(n491) );
  NAND2_X1 U543 ( .A1(n491), .A2(n510), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n486), .B(n485), .ZN(G1328GAT) );
  NAND2_X1 U545 ( .A1(n512), .A2(n491), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n487), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT40), .B(KEYINPUT99), .Z(n489) );
  NAND2_X1 U548 ( .A1(n491), .A2(n515), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U550 ( .A(G43GAT), .B(n490), .ZN(G1330GAT) );
  NAND2_X1 U551 ( .A1(n491), .A2(n527), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n492), .B(KEYINPUT100), .ZN(n493) );
  XNOR2_X1 U553 ( .A(G50GAT), .B(n493), .ZN(G1331GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT101), .B(KEYINPUT42), .Z(n498) );
  NAND2_X1 U555 ( .A1(n555), .A2(n494), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n495), .B(KEYINPUT102), .ZN(n509) );
  NOR2_X1 U557 ( .A1(n509), .A2(n496), .ZN(n503) );
  NAND2_X1 U558 ( .A1(n503), .A2(n510), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U560 ( .A(G57GAT), .B(n499), .ZN(G1332GAT) );
  NAND2_X1 U561 ( .A1(n512), .A2(n503), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U563 ( .A(G71GAT), .B(KEYINPUT103), .Z(n502) );
  NAND2_X1 U564 ( .A1(n503), .A2(n515), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n502), .B(n501), .ZN(G1334GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT104), .B(KEYINPUT43), .Z(n505) );
  NAND2_X1 U567 ( .A1(n503), .A2(n527), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(n507) );
  XOR2_X1 U569 ( .A(G78GAT), .B(KEYINPUT105), .Z(n506) );
  XNOR2_X1 U570 ( .A(n507), .B(n506), .ZN(G1335GAT) );
  NOR2_X1 U571 ( .A1(n509), .A2(n508), .ZN(n518) );
  NAND2_X1 U572 ( .A1(n510), .A2(n518), .ZN(n511) );
  XNOR2_X1 U573 ( .A(G85GAT), .B(n511), .ZN(G1336GAT) );
  NAND2_X1 U574 ( .A1(n512), .A2(n518), .ZN(n513) );
  XNOR2_X1 U575 ( .A(n513), .B(KEYINPUT106), .ZN(n514) );
  XNOR2_X1 U576 ( .A(G92GAT), .B(n514), .ZN(G1337GAT) );
  XOR2_X1 U577 ( .A(G99GAT), .B(KEYINPUT107), .Z(n517) );
  NAND2_X1 U578 ( .A1(n518), .A2(n515), .ZN(n516) );
  XNOR2_X1 U579 ( .A(n517), .B(n516), .ZN(G1338GAT) );
  NAND2_X1 U580 ( .A1(n518), .A2(n527), .ZN(n519) );
  XNOR2_X1 U581 ( .A(n519), .B(KEYINPUT44), .ZN(n520) );
  XNOR2_X1 U582 ( .A(G106GAT), .B(n520), .ZN(G1339GAT) );
  NOR2_X1 U583 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U584 ( .A(n523), .B(KEYINPUT111), .ZN(n540) );
  NOR2_X1 U585 ( .A1(n524), .A2(n540), .ZN(n525) );
  XOR2_X1 U586 ( .A(KEYINPUT112), .B(n525), .Z(n526) );
  NOR2_X1 U587 ( .A1(n527), .A2(n526), .ZN(n535) );
  NAND2_X1 U588 ( .A1(n535), .A2(n563), .ZN(n528) );
  XNOR2_X1 U589 ( .A(G113GAT), .B(n528), .ZN(G1340GAT) );
  XOR2_X1 U590 ( .A(G120GAT), .B(KEYINPUT49), .Z(n530) );
  NAND2_X1 U591 ( .A1(n535), .A2(n555), .ZN(n529) );
  XNOR2_X1 U592 ( .A(n530), .B(n529), .ZN(G1341GAT) );
  XNOR2_X1 U593 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n534) );
  XOR2_X1 U594 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n532) );
  NAND2_X1 U595 ( .A1(n535), .A2(n573), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n534), .B(n533), .ZN(G1342GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT51), .B(KEYINPUT115), .Z(n537) );
  NAND2_X1 U599 ( .A1(n535), .A2(n388), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U601 ( .A(G134GAT), .B(n538), .Z(G1343GAT) );
  NOR2_X1 U602 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U603 ( .A(n541), .B(KEYINPUT116), .ZN(n547) );
  NAND2_X1 U604 ( .A1(n547), .A2(n563), .ZN(n542) );
  XNOR2_X1 U605 ( .A(n542), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n544) );
  NAND2_X1 U607 ( .A1(n547), .A2(n555), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(n545), .ZN(G1345GAT) );
  NAND2_X1 U610 ( .A1(n547), .A2(n573), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n546), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U612 ( .A(G162GAT), .B(KEYINPUT117), .Z(n549) );
  NAND2_X1 U613 ( .A1(n388), .A2(n547), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(G1347GAT) );
  NAND2_X1 U615 ( .A1(n563), .A2(n558), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(KEYINPUT118), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G169GAT), .B(n551), .ZN(G1348GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT57), .B(KEYINPUT120), .Z(n553) );
  XNOR2_X1 U619 ( .A(G176GAT), .B(KEYINPUT119), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U621 ( .A(KEYINPUT56), .B(n554), .Z(n557) );
  NAND2_X1 U622 ( .A1(n558), .A2(n555), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1349GAT) );
  NAND2_X1 U624 ( .A1(n573), .A2(n558), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U627 ( .A(n562), .B(KEYINPUT123), .Z(n576) );
  INV_X1 U628 ( .A(n576), .ZN(n572) );
  NAND2_X1 U629 ( .A1(n572), .A2(n563), .ZN(n565) );
  XOR2_X1 U630 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XOR2_X1 U632 ( .A(n566), .B(KEYINPUT124), .Z(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .Z(n571) );
  OR2_X1 U636 ( .A1(n569), .A2(n576), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1353GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(KEYINPUT126), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G211GAT), .B(n575), .ZN(G1354GAT) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n579) );
  XNOR2_X1 U642 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

