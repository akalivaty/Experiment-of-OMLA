//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n450, new_n452, new_n453, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1106,
    new_n1107, new_n1108, new_n1109;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  INV_X1    g026(.A(G2106), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT68), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NOR4_X1   g031(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI22_X1  g035(.A1(new_n456), .A2(new_n452), .B1(new_n460), .B2(new_n457), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT69), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(G125), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n468), .A2(new_n469), .B1(G113), .B2(G2104), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n465), .A2(new_n467), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(KEYINPUT70), .A3(G125), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n463), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n464), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  OAI21_X1  g050(.A(KEYINPUT71), .B1(new_n466), .B2(G2104), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT71), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(new_n464), .A3(KEYINPUT3), .ZN(new_n478));
  NAND4_X1  g053(.A1(new_n476), .A2(new_n478), .A3(new_n463), .A4(new_n467), .ZN(new_n479));
  INV_X1    g054(.A(G137), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n475), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(KEYINPUT72), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT72), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(new_n475), .C1(new_n479), .C2(new_n480), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n473), .B1(new_n482), .B2(new_n484), .ZN(G160));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G112), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n479), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  XOR2_X1   g065(.A(new_n490), .B(KEYINPUT73), .Z(new_n491));
  NAND4_X1  g066(.A1(new_n476), .A2(new_n478), .A3(G2105), .A4(new_n467), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  AOI211_X1 g068(.A(new_n488), .B(new_n491), .C1(G124), .C2(new_n493), .ZN(G162));
  INV_X1    g069(.A(KEYINPUT74), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  AND4_X1   g072(.A1(new_n463), .A2(new_n497), .A3(new_n465), .A4(new_n467), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n466), .A2(KEYINPUT71), .A3(G2104), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n501), .A2(G138), .A3(new_n463), .A4(new_n476), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n498), .B1(new_n502), .B2(KEYINPUT4), .ZN(new_n503));
  INV_X1    g078(.A(G126), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n463), .A2(G114), .ZN(new_n505));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  OAI22_X1  g081(.A1(new_n492), .A2(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n495), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT4), .B1(new_n479), .B2(new_n496), .ZN(new_n509));
  INV_X1    g084(.A(new_n498), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n507), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT74), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(G164));
  XNOR2_X1  g090(.A(KEYINPUT5), .B(G543), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  AND2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n516), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n521), .A2(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n520), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(G166));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n525), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n516), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n524), .A2(G89), .ZN(new_n536));
  NAND2_X1  g111(.A1(G63), .A2(G651), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n534), .A2(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n541), .A2(new_n525), .B1(new_n526), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n518), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n543), .A2(new_n545), .ZN(G171));
  AOI22_X1  g121(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n518), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT75), .ZN(new_n549));
  INV_X1    g124(.A(new_n526), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n522), .A2(new_n523), .ZN(new_n551));
  INV_X1    g126(.A(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n550), .A2(G81), .B1(new_n553), .B2(G43), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(new_n553), .A2(G53), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n535), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(G91), .A2(new_n550), .B1(new_n567), .B2(G651), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n564), .A2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  XOR2_X1   g145(.A(new_n529), .B(KEYINPUT76), .Z(G303));
  NAND2_X1  g146(.A1(new_n550), .A2(G87), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n553), .A2(G49), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  AND2_X1   g150(.A1(new_n516), .A2(G61), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT77), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n579), .B1(new_n576), .B2(KEYINPUT77), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n550), .A2(G86), .B1(new_n553), .B2(G48), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G305));
  INV_X1    g158(.A(G47), .ZN(new_n584));
  INV_X1    g159(.A(G85), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n584), .A2(new_n525), .B1(new_n526), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n518), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n516), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G54), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n518), .A2(new_n592), .B1(new_n525), .B2(new_n593), .ZN(new_n594));
  XOR2_X1   g169(.A(new_n594), .B(KEYINPUT79), .Z(new_n595));
  NAND2_X1  g170(.A1(new_n550), .A2(G92), .ZN(new_n596));
  XOR2_X1   g171(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n591), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n591), .B1(new_n600), .B2(G868), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G299), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G297));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n600), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g187(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n613));
  INV_X1    g188(.A(G111), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n613), .A2(KEYINPUT82), .B1(new_n614), .B2(G2105), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(KEYINPUT82), .B2(new_n613), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n489), .A2(G135), .ZN(new_n617));
  AND2_X1   g192(.A1(new_n493), .A2(G123), .ZN(new_n618));
  AND2_X1   g193(.A1(new_n618), .A2(KEYINPUT81), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n618), .A2(KEYINPUT81), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n616), .B(new_n617), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(KEYINPUT83), .B(G2096), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT80), .B(G2100), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n625), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n623), .A2(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n633), .A2(KEYINPUT14), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT84), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2451), .B(G2454), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n636), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n639), .B(new_n640), .Z(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT85), .ZN(new_n644));
  INV_X1    g219(.A(G14), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n645), .B1(new_n641), .B2(new_n642), .ZN(new_n646));
  AND2_X1   g221(.A1(new_n644), .A2(new_n646), .ZN(G401));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g225(.A1(new_n650), .A2(KEYINPUT17), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n648), .A2(new_n649), .ZN(new_n652));
  AOI21_X1  g227(.A(KEYINPUT18), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2072), .B(G2078), .Z(new_n654));
  AOI21_X1  g229(.A(new_n654), .B1(new_n650), .B2(KEYINPUT18), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n653), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2096), .B(G2100), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1961), .B(G1966), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT86), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1956), .B(G2474), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT20), .Z(new_n667));
  NOR2_X1   g242(.A1(new_n660), .A2(new_n662), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n669), .A2(new_n665), .A3(new_n663), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n667), .B(new_n670), .C1(new_n665), .C2(new_n669), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT87), .ZN(new_n672));
  XOR2_X1   g247(.A(G1981), .B(G1986), .Z(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n672), .B(new_n677), .ZN(G229));
  INV_X1    g253(.A(G29), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n679), .A2(G33), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT97), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT96), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT25), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n683), .A2(KEYINPUT96), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n683), .A2(KEYINPUT96), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n687), .A2(KEYINPUT25), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n471), .A2(G127), .ZN(new_n690));
  INV_X1    g265(.A(G115), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(new_n464), .ZN(new_n692));
  AOI22_X1  g267(.A1(new_n692), .A2(G2105), .B1(G139), .B2(new_n489), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n686), .A2(new_n689), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT98), .Z(new_n695));
  INV_X1    g270(.A(KEYINPUT99), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n680), .B1(new_n697), .B2(G29), .ZN(new_n698));
  INV_X1    g273(.A(G2072), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NOR2_X1   g276(.A1(G168), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(new_n701), .B2(G21), .ZN(new_n703));
  INV_X1    g278(.A(G1966), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n701), .A2(G5), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G171), .B2(new_n701), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n705), .B1(G1961), .B2(new_n707), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n621), .A2(new_n679), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT31), .B(G11), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT30), .B(G28), .Z(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(G29), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n703), .B2(new_n704), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n708), .A2(new_n709), .A3(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT101), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n679), .A2(G32), .ZN(new_n718));
  NAND3_X1  g293(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT26), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n721), .A2(new_n722), .B1(G105), .B2(new_n474), .ZN(new_n723));
  INV_X1    g298(.A(G129), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n492), .B2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G141), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(new_n479), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n718), .B1(new_n729), .B2(new_n679), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT27), .B(G1996), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n707), .A2(G1961), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n716), .A2(new_n717), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(G164), .A2(new_n679), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G27), .B2(new_n679), .ZN(new_n737));
  INV_X1    g312(.A(G2078), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  INV_X1    g315(.A(G34), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n741), .A2(KEYINPUT24), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(KEYINPUT24), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n679), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G160), .B2(new_n679), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT100), .B(G2084), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n739), .A2(new_n740), .A3(new_n747), .ZN(new_n748));
  NOR3_X1   g323(.A1(new_n700), .A2(new_n735), .A3(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT102), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n679), .A2(G35), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G162), .B2(new_n679), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT29), .ZN(new_n754));
  INV_X1    g329(.A(G2090), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n701), .A2(G4), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n600), .B2(new_n701), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT92), .B(G1348), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n701), .A2(G19), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT93), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n556), .B2(new_n701), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1341), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n701), .A2(G20), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT103), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT23), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G299), .B2(G16), .ZN(new_n768));
  INV_X1    g343(.A(G1956), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n764), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n679), .A2(G26), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT28), .Z(new_n773));
  OR2_X1    g348(.A1(G104), .A2(G2105), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n774), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n775));
  INV_X1    g350(.A(G128), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n492), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n489), .B2(G140), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT94), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n773), .B1(new_n779), .B2(G29), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT95), .B(G2067), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n756), .A2(new_n760), .A3(new_n771), .A4(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n749), .B2(new_n750), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n751), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT36), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n701), .A2(G22), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G166), .B2(new_n701), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1971), .ZN(new_n789));
  INV_X1    g364(.A(G305), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n790), .A2(new_n701), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G6), .B2(new_n701), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT32), .B(G1981), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT89), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n789), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n792), .A2(new_n794), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n701), .A2(G23), .ZN(new_n797));
  INV_X1    g372(.A(G288), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(new_n701), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT90), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT33), .B(G1976), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n795), .A2(new_n796), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n803), .A2(KEYINPUT34), .ZN(new_n804));
  NOR2_X1   g379(.A1(G16), .A2(G24), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n589), .B2(G16), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT88), .ZN(new_n807));
  INV_X1    g382(.A(G1986), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n679), .A2(G25), .ZN(new_n810));
  INV_X1    g385(.A(G119), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n463), .A2(G107), .ZN(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n813));
  OAI22_X1  g388(.A1(new_n492), .A2(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n489), .B2(G131), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n810), .B1(new_n815), .B2(new_n679), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT35), .B(G1991), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n809), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n804), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT91), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n803), .A2(KEYINPUT34), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n786), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n821), .A2(new_n786), .A3(new_n822), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n785), .B1(new_n824), .B2(new_n825), .ZN(G311));
  INV_X1    g401(.A(new_n825), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n751), .B(new_n784), .C1(new_n827), .C2(new_n823), .ZN(G150));
  AOI22_X1  g403(.A1(new_n550), .A2(G93), .B1(new_n553), .B2(G55), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n518), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G860), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT105), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT37), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n599), .A2(new_n607), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n555), .B(new_n831), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n841));
  INV_X1    g416(.A(G860), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n840), .B2(KEYINPUT39), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n834), .B1(new_n841), .B2(new_n843), .ZN(G145));
  XNOR2_X1  g419(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n845));
  INV_X1    g420(.A(G37), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n815), .B(KEYINPUT106), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n627), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n489), .A2(G142), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n493), .A2(G130), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n463), .A2(G118), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n849), .B(new_n850), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n848), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n511), .A2(new_n512), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n779), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n728), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n697), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n695), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n854), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT108), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n621), .B(G160), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(G162), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n858), .A2(new_n854), .A3(new_n859), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n866), .B(new_n867), .C1(new_n860), .C2(new_n861), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n846), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n867), .B1(new_n860), .B2(KEYINPUT107), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT107), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n858), .A2(new_n872), .A3(new_n854), .A4(new_n859), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n866), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n845), .B1(new_n870), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n845), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n869), .A2(new_n874), .A3(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n876), .A2(new_n878), .ZN(G395));
  XNOR2_X1  g454(.A(new_n599), .B(G299), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT110), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(KEYINPUT41), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n599), .B(new_n604), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT41), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n882), .B1(new_n885), .B2(KEYINPUT111), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n886), .B1(KEYINPUT111), .B2(new_n885), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n609), .B(new_n838), .Z(new_n888));
  MUX2_X1   g463(.A(new_n881), .B(new_n887), .S(new_n888), .Z(new_n889));
  XNOR2_X1  g464(.A(new_n529), .B(new_n798), .ZN(new_n890));
  XNOR2_X1  g465(.A(G305), .B(G290), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n890), .B(new_n891), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n892), .B(KEYINPUT42), .Z(new_n893));
  XNOR2_X1  g468(.A(new_n889), .B(new_n893), .ZN(new_n894));
  MUX2_X1   g469(.A(new_n831), .B(new_n894), .S(G868), .Z(G295));
  MUX2_X1   g470(.A(new_n831), .B(new_n894), .S(G868), .Z(G331));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n897));
  XNOR2_X1  g472(.A(G171), .B(KEYINPUT112), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n838), .B(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(G286), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n883), .ZN(new_n901));
  INV_X1    g476(.A(new_n892), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n901), .B(new_n902), .C1(new_n887), .C2(new_n900), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n846), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n887), .A2(new_n900), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n902), .B1(new_n905), .B2(new_n901), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n897), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n902), .B1(new_n900), .B2(new_n881), .ZN(new_n908));
  INV_X1    g483(.A(new_n900), .ZN(new_n909));
  INV_X1    g484(.A(new_n882), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n885), .B1(new_n910), .B2(KEYINPUT113), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n880), .A2(KEYINPUT113), .A3(KEYINPUT41), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n908), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n914), .A2(KEYINPUT43), .A3(new_n846), .A4(new_n903), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n907), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT44), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT43), .B1(new_n904), .B2(new_n906), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n914), .A2(new_n897), .A3(new_n846), .A4(new_n903), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n917), .A2(new_n922), .ZN(G397));
  INV_X1    g498(.A(KEYINPUT45), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n924), .B1(new_n925), .B2(G1384), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n482), .A2(new_n484), .ZN(new_n927));
  INV_X1    g502(.A(new_n473), .ZN(new_n928));
  XNOR2_X1  g503(.A(KEYINPUT114), .B(G40), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n926), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G2067), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n779), .B(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G1996), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n728), .B(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n815), .B(new_n817), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n932), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(G290), .A2(G1986), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n932), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(KEYINPUT48), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n934), .A2(new_n729), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT127), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n944), .A2(new_n932), .B1(new_n945), .B2(KEYINPUT46), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(KEYINPUT46), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(new_n932), .B2(new_n935), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n932), .A2(new_n935), .A3(new_n947), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  XOR2_X1   g525(.A(new_n950), .B(KEYINPUT47), .Z(new_n951));
  NAND2_X1  g526(.A1(new_n815), .A2(new_n817), .ZN(new_n952));
  OAI22_X1  g527(.A1(new_n937), .A2(new_n952), .B1(G2067), .B2(new_n779), .ZN(new_n953));
  AOI211_X1 g528(.A(new_n943), .B(new_n951), .C1(new_n932), .C2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G1384), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n855), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n931), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(KEYINPUT116), .B(G8), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OR2_X1    g534(.A1(G305), .A2(G1981), .ZN(new_n960));
  NAND2_X1  g535(.A1(G305), .A2(G1981), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT49), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n960), .A2(KEYINPUT49), .A3(new_n961), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n959), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G1976), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n966), .A2(new_n967), .A3(new_n798), .ZN(new_n968));
  XOR2_X1   g543(.A(new_n960), .B(KEYINPUT117), .Z(new_n969));
  OAI21_X1  g544(.A(new_n959), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(G303), .A2(G8), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT55), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n971), .B(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G8), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(new_n514), .B2(new_n955), .ZN(new_n976));
  OAI211_X1 g551(.A(G160), .B(new_n930), .C1(new_n956), .C2(KEYINPUT50), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n755), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n925), .A2(G1384), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n931), .B1(new_n980), .B2(KEYINPUT45), .ZN(new_n981));
  AOI21_X1  g556(.A(G1384), .B1(new_n508), .B2(new_n513), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n981), .B1(KEYINPUT45), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1971), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n974), .B1(new_n979), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n973), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n959), .B1(new_n967), .B2(G288), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT52), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(new_n798), .B2(G1976), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n966), .B(new_n989), .C1(new_n988), .C2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n970), .B1(new_n987), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n992), .B1(new_n973), .B2(new_n986), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT118), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT45), .B1(new_n855), .B2(new_n955), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n995), .B1(new_n996), .B2(new_n931), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n926), .A2(KEYINPUT118), .A3(G160), .A4(new_n930), .ZN(new_n998));
  INV_X1    g573(.A(new_n513), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT74), .B1(new_n511), .B2(new_n512), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT45), .B(new_n955), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n704), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n925), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1004), .A2(new_n931), .ZN(new_n1005));
  INV_X1    g580(.A(G2084), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1005), .B(new_n1006), .C1(new_n975), .C2(new_n982), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n958), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(G286), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n994), .B(new_n1011), .C1(new_n973), .C2(new_n986), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n993), .B1(new_n1012), .B2(KEYINPUT63), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n1010), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(new_n983), .B2(G2078), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n738), .A2(KEYINPUT53), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT120), .B1(new_n976), .B2(new_n977), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT120), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1005), .B(new_n1019), .C1(new_n975), .C2(new_n982), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  OAI221_X1 g596(.A(new_n1016), .B1(new_n1002), .B2(new_n1017), .C1(new_n1021), .C2(G1961), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(G171), .ZN(new_n1023));
  NOR2_X1   g598(.A1(G168), .A2(new_n958), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(KEYINPUT51), .ZN(new_n1025));
  AOI22_X1  g600(.A1(new_n978), .A2(new_n1006), .B1(new_n1002), .B2(new_n704), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1025), .B1(new_n1026), .B2(new_n958), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1024), .B1(new_n1008), .B2(G8), .ZN(new_n1028));
  XOR2_X1   g603(.A(KEYINPUT126), .B(KEYINPUT51), .Z(new_n1029));
  OAI21_X1  g604(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1008), .A2(new_n1024), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1023), .B1(new_n1032), .B2(KEYINPUT62), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT62), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1030), .A2(new_n1034), .A3(new_n1031), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1014), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n985), .ZN(new_n1037));
  AOI211_X1 g612(.A(KEYINPUT50), .B(G1384), .C1(new_n508), .C2(new_n513), .ZN(new_n1038));
  OAI211_X1 g613(.A(G160), .B(new_n930), .C1(new_n980), .C2(new_n975), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1038), .A2(new_n1039), .A3(G2090), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1009), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n994), .B1(new_n973), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1013), .B1(new_n1036), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1043), .ZN(new_n1045));
  XOR2_X1   g620(.A(G171), .B(KEYINPUT54), .Z(new_n1046));
  NAND2_X1  g621(.A1(new_n1022), .A2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(G160), .A2(KEYINPUT53), .A3(G40), .A4(new_n738), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1048), .B1(KEYINPUT45), .B2(new_n980), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1046), .B1(new_n1049), .B2(new_n926), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1016), .B(new_n1050), .C1(new_n1021), .C2(G1961), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1045), .A2(new_n1032), .A3(new_n1047), .A4(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT57), .B1(new_n564), .B2(KEYINPUT119), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1053), .B(G299), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT56), .B(G2072), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n981), .B(new_n1055), .C1(KEYINPUT45), .C2(new_n982), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n769), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1054), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(new_n1057), .A3(new_n1054), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(KEYINPUT61), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT61), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1060), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1062), .B1(new_n1063), .B2(new_n1058), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n983), .A2(G1996), .ZN(new_n1066));
  XOR2_X1   g641(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n1067));
  XNOR2_X1  g642(.A(new_n1067), .B(G1341), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n931), .B2(new_n956), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1069), .B(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n556), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT123), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT59), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1073), .A3(KEYINPUT59), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1065), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1018), .A2(new_n759), .A3(new_n1020), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n957), .A2(new_n933), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT60), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT124), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1083), .A2(new_n1084), .A3(new_n600), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1081), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT60), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT60), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT124), .B1(new_n1088), .B2(new_n599), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1085), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1087), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1078), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1059), .B1(new_n1086), .B2(new_n599), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1060), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1052), .B1(new_n1095), .B2(KEYINPUT125), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT125), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1092), .A2(new_n1097), .A3(new_n1094), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1044), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n589), .A2(new_n808), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n932), .B1(new_n1100), .B2(new_n940), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1101), .B(KEYINPUT115), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n939), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n954), .B1(new_n1099), .B2(new_n1103), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g679(.A(G319), .ZN(new_n1106));
  OR3_X1    g680(.A1(G229), .A2(new_n1106), .A3(G227), .ZN(new_n1107));
  AOI21_X1  g681(.A(new_n1107), .B1(new_n644), .B2(new_n646), .ZN(new_n1108));
  OAI21_X1  g682(.A(new_n1108), .B1(new_n869), .B2(new_n874), .ZN(new_n1109));
  AOI21_X1  g683(.A(new_n1109), .B1(new_n918), .B2(new_n919), .ZN(G308));
  OAI211_X1 g684(.A(new_n920), .B(new_n1108), .C1(new_n874), .C2(new_n869), .ZN(G225));
endmodule


