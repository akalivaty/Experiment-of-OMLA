//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031;
  NAND2_X1  g000(.A1(KEYINPUT76), .A2(G125), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  NAND3_X1  g003(.A1(KEYINPUT76), .A2(G125), .A3(G140), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(KEYINPUT16), .A3(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G140), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  XNOR2_X1  g010(.A(G125), .B(G140), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  XOR2_X1   g013(.A(KEYINPUT24), .B(G110), .Z(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G119), .ZN(new_n202));
  INV_X1    g016(.A(G119), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT75), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT75), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n200), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n203), .A2(G128), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n210), .B(new_n204), .C1(new_n211), .C2(KEYINPUT23), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G110), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n196), .B(new_n199), .C1(new_n209), .C2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(G110), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n207), .A2(new_n208), .A3(new_n200), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n191), .A2(new_n198), .A3(new_n194), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n198), .B1(new_n191), .B2(new_n194), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT79), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT79), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n214), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT22), .B(G137), .ZN(new_n224));
  INV_X1    g038(.A(G953), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(G221), .A3(G234), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n224), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n227), .B(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n221), .A2(new_n223), .A3(new_n230), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n229), .A2(new_n222), .A3(new_n219), .A4(new_n214), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G902), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(KEYINPUT25), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT80), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT25), .B1(new_n233), .B2(new_n234), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT80), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G234), .ZN(new_n241));
  OAI21_X1  g055(.A(G217), .B1(new_n241), .B2(G902), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n242), .B(KEYINPUT74), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n233), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n242), .A2(new_n234), .ZN(new_n246));
  OAI22_X1  g060(.A1(new_n238), .A2(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT98), .ZN(new_n248));
  INV_X1    g062(.A(G237), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(new_n225), .A3(G214), .ZN(new_n250));
  INV_X1    g064(.A(G143), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n249), .A2(new_n225), .A3(G143), .A4(G214), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XOR2_X1   g068(.A(KEYINPUT65), .B(G131), .Z(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n248), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT17), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n252), .A2(new_n253), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT98), .A3(new_n255), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n254), .A2(new_n256), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n257), .A2(new_n258), .A3(new_n260), .A4(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n260), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT98), .B1(new_n259), .B2(new_n255), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT17), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n217), .A2(new_n218), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n262), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n190), .ZN(new_n268));
  AOI21_X1  g082(.A(G140), .B1(KEYINPUT76), .B2(G125), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT96), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT96), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n189), .A2(new_n271), .A3(new_n190), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n198), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT97), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(KEYINPUT18), .A2(G131), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n259), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n252), .A2(KEYINPUT18), .A3(G131), .A4(new_n253), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n199), .A2(KEYINPUT97), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n275), .B(new_n279), .C1(new_n273), .C2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(G113), .B(G122), .ZN(new_n282));
  INV_X1    g096(.A(G104), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n282), .B(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n284), .B(KEYINPUT100), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n267), .A2(new_n281), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n284), .B1(new_n267), .B2(new_n281), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n234), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT101), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(KEYINPUT101), .B(new_n234), .C1(new_n286), .C2(new_n287), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(G475), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n281), .ZN(new_n293));
  INV_X1    g107(.A(new_n266), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n257), .A2(new_n260), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n294), .B1(new_n295), .B2(KEYINPUT17), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n293), .B1(new_n296), .B2(new_n262), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n257), .A2(new_n260), .A3(new_n261), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n196), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT96), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n271), .B1(new_n189), .B2(new_n190), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT19), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT19), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n197), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(KEYINPUT99), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT99), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n306), .B(KEYINPUT19), .C1(new_n300), .C2(new_n301), .ZN(new_n307));
  AOI21_X1  g121(.A(G146), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n281), .B1(new_n299), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n284), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n297), .A2(new_n285), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(G475), .A2(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT20), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT20), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n309), .A2(new_n310), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n315), .B(new_n312), .C1(new_n316), .C2(new_n286), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G116), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(KEYINPUT14), .A3(G122), .ZN(new_n320));
  XOR2_X1   g134(.A(G116), .B(G122), .Z(new_n321));
  OAI211_X1 g135(.A(G107), .B(new_n320), .C1(new_n321), .C2(KEYINPUT14), .ZN(new_n322));
  OR2_X1    g136(.A1(KEYINPUT82), .A2(G107), .ZN(new_n323));
  NAND2_X1  g137(.A1(KEYINPUT82), .A2(G107), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n251), .A2(G128), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n201), .A2(G143), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G134), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n328), .A2(new_n329), .ZN(new_n331));
  OAI221_X1 g145(.A(new_n322), .B1(new_n325), .B2(new_n321), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n321), .B(new_n325), .ZN(new_n333));
  INV_X1    g147(.A(new_n330), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT13), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n326), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n327), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n326), .A2(new_n335), .ZN(new_n338));
  OAI21_X1  g152(.A(G134), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n333), .A2(new_n334), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n332), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT9), .B(G234), .ZN(new_n342));
  INV_X1    g156(.A(G217), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n342), .A2(new_n343), .A3(G953), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n332), .A2(new_n340), .A3(new_n344), .ZN(new_n347));
  AOI21_X1  g161(.A(G902), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G478), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n349), .A2(KEYINPUT15), .ZN(new_n350));
  OR2_X1    g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n348), .A2(new_n350), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(G234), .A2(G237), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(G952), .A3(new_n225), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT21), .B(G898), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n355), .A2(G902), .A3(G953), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n356), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  XOR2_X1   g174(.A(new_n360), .B(KEYINPUT102), .Z(new_n361));
  NAND4_X1  g175(.A1(new_n292), .A2(new_n318), .A3(new_n354), .A4(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT11), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n329), .B2(G137), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n329), .A2(G137), .ZN(new_n365));
  INV_X1    g179(.A(G137), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(KEYINPUT11), .A3(G134), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n364), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  OR2_X1    g182(.A1(new_n368), .A2(new_n255), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT66), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n364), .A2(new_n367), .A3(KEYINPUT66), .A4(new_n365), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G131), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n369), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT64), .ZN(new_n375));
  XNOR2_X1  g189(.A(G143), .B(G146), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT0), .B(G128), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AND2_X1   g192(.A1(KEYINPUT0), .A2(G128), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n198), .A2(G143), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n251), .A2(G146), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(KEYINPUT0), .A2(G128), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(new_n385), .A3(KEYINPUT64), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n378), .A2(new_n380), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n374), .A2(new_n387), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n251), .A2(KEYINPUT1), .A3(G146), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(new_n383), .B2(new_n201), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(new_n381), .A3(new_n382), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n365), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n329), .A2(G137), .ZN(new_n395));
  OAI21_X1  g209(.A(G131), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n369), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n388), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n203), .A2(G116), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n319), .A2(G119), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT68), .ZN(new_n404));
  NOR2_X1   g218(.A1(KEYINPUT2), .A2(G113), .ZN(new_n405));
  NAND2_X1  g219(.A1(KEYINPUT2), .A2(G113), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT67), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT67), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(KEYINPUT2), .A3(G113), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n405), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  OR2_X1    g224(.A1(new_n404), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n404), .A2(new_n410), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n400), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT69), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n374), .A2(new_n416), .A3(new_n387), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n416), .B1(new_n374), .B2(new_n387), .ZN(new_n418));
  OAI211_X1 g232(.A(KEYINPUT30), .B(new_n397), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT70), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n397), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n368), .A2(new_n255), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n372), .A2(G131), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n368), .A2(new_n370), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n378), .A2(new_n380), .A3(new_n386), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT69), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n374), .A2(new_n416), .A3(new_n387), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n422), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(KEYINPUT70), .B1(new_n430), .B2(KEYINPUT30), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n415), .B1(new_n421), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT71), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n404), .A2(new_n410), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n404), .A2(new_n410), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n411), .A2(KEYINPUT71), .A3(new_n412), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n430), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n249), .A2(new_n225), .A3(G210), .ZN(new_n441));
  XOR2_X1   g255(.A(new_n441), .B(KEYINPUT27), .Z(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT26), .B(G101), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n442), .B(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(KEYINPUT29), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n432), .A2(new_n440), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT29), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n430), .A2(new_n439), .ZN(new_n449));
  AOI211_X1 g263(.A(new_n422), .B(new_n438), .C1(new_n428), .C2(new_n429), .ZN(new_n450));
  OAI21_X1  g264(.A(KEYINPUT28), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n388), .A2(new_n437), .A3(new_n436), .A4(new_n397), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT28), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(KEYINPUT73), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT73), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n456), .B1(new_n452), .B2(new_n453), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n448), .B1(new_n451), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n430), .A2(KEYINPUT28), .A3(new_n439), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n398), .A2(new_n413), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n454), .A3(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n445), .B1(new_n462), .B2(KEYINPUT29), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n447), .B(new_n234), .C1(new_n459), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n419), .A2(new_n420), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n428), .A2(new_n429), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n466), .A2(KEYINPUT70), .A3(KEYINPUT30), .A4(new_n397), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n414), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n445), .A2(KEYINPUT72), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n440), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(KEYINPUT31), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT31), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n440), .A2(new_n472), .A3(new_n469), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n432), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n462), .A2(new_n444), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n471), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(G472), .A2(G902), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT32), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n464), .A2(G472), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n476), .A2(new_n477), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n479), .ZN(new_n483));
  AOI211_X1 g297(.A(new_n247), .B(new_n362), .C1(new_n481), .C2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(G214), .B1(G237), .B2(G902), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n383), .A2(new_n201), .ZN(new_n486));
  INV_X1    g300(.A(new_n389), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n486), .A2(new_n392), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT91), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(new_n489), .A3(new_n193), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT91), .B1(new_n393), .B2(G125), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n490), .B(new_n491), .C1(new_n193), .C2(new_n387), .ZN(new_n492));
  INV_X1    g306(.A(G224), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(G953), .ZN(new_n494));
  XOR2_X1   g308(.A(new_n492), .B(new_n494), .Z(new_n495));
  XNOR2_X1  g309(.A(G110), .B(G122), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT3), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G104), .ZN(new_n499));
  AND2_X1   g313(.A1(KEYINPUT82), .A2(G107), .ZN(new_n500));
  NOR2_X1   g314(.A1(KEYINPUT82), .A2(G107), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(G107), .B1(new_n283), .B2(KEYINPUT3), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n283), .A2(KEYINPUT3), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT83), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT4), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n504), .A2(new_n323), .A3(new_n324), .ZN(new_n508));
  INV_X1    g322(.A(G107), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n509), .B1(new_n498), .B2(G104), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n499), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT83), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n508), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n506), .A2(new_n507), .A3(new_n513), .A4(G101), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n413), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n506), .A2(G101), .A3(new_n513), .ZN(new_n516));
  INV_X1    g330(.A(G101), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n508), .A2(new_n511), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT84), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n507), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n506), .A2(new_n519), .A3(new_n513), .A4(G101), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n515), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(G116), .B(G119), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n410), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n517), .B1(G104), .B2(G107), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n526), .B1(new_n325), .B2(G104), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n518), .A3(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n401), .A2(KEYINPUT5), .ZN(new_n529));
  INV_X1    g343(.A(G113), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n524), .A2(KEYINPUT5), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT88), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n531), .A2(KEYINPUT88), .A3(new_n532), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n528), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n497), .B1(new_n523), .B2(new_n537), .ZN(new_n538));
  XOR2_X1   g352(.A(KEYINPUT90), .B(KEYINPUT6), .Z(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n508), .A2(new_n511), .A3(new_n512), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n512), .B1(new_n508), .B2(new_n511), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n542), .A2(new_n543), .A3(new_n517), .ZN(new_n544));
  INV_X1    g358(.A(new_n520), .ZN(new_n545));
  OAI211_X1 g359(.A(KEYINPUT4), .B(new_n522), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n515), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n537), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT6), .B1(new_n548), .B2(new_n496), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n523), .A2(new_n497), .A3(new_n537), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT89), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n548), .A2(new_n496), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT89), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n552), .A2(new_n538), .A3(new_n553), .A4(KEYINPUT6), .ZN(new_n554));
  AOI211_X1 g368(.A(new_n495), .B(new_n541), .C1(new_n551), .C2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT7), .ZN(new_n556));
  OR3_X1    g370(.A1(new_n492), .A2(new_n556), .A3(new_n494), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n492), .A2(new_n494), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n492), .A2(new_n556), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n535), .A2(new_n536), .B1(new_n410), .B2(new_n524), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n518), .A2(new_n527), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n532), .A2(KEYINPUT93), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n532), .A2(KEYINPUT93), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n563), .A2(new_n531), .A3(new_n564), .ZN(new_n565));
  OAI22_X1  g379(.A1(new_n560), .A2(new_n562), .B1(new_n565), .B2(new_n528), .ZN(new_n566));
  XOR2_X1   g380(.A(KEYINPUT92), .B(KEYINPUT8), .Z(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(new_n496), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n557), .A2(new_n558), .A3(new_n559), .A4(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n234), .B1(new_n570), .B2(new_n550), .ZN(new_n571));
  OAI21_X1  g385(.A(G210), .B1(G237), .B2(G902), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(KEYINPUT94), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n555), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n573), .ZN(new_n575));
  INV_X1    g389(.A(new_n495), .ZN(new_n576));
  INV_X1    g390(.A(new_n541), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT6), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n546), .A2(new_n547), .ZN(new_n579));
  INV_X1    g393(.A(new_n537), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n578), .B1(new_n581), .B2(new_n497), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n553), .B1(new_n582), .B2(new_n552), .ZN(new_n583));
  INV_X1    g397(.A(new_n554), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n576), .B(new_n577), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n571), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n575), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n485), .B1(new_n574), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT95), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(G221), .B1(new_n342), .B2(G902), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(G469), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(new_n234), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n514), .A2(new_n387), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n546), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n392), .A2(KEYINPUT85), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT85), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n376), .A2(new_n599), .A3(new_n391), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n390), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n601), .A2(new_n518), .A3(new_n527), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n562), .A2(KEYINPUT10), .A3(new_n393), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n597), .A2(new_n607), .A3(new_n426), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n595), .B1(new_n521), .B2(new_n522), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n374), .B1(new_n609), .B2(new_n606), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n225), .A2(G227), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT81), .ZN(new_n613));
  XNOR2_X1  g427(.A(G110), .B(G140), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT86), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n609), .A2(new_n374), .A3(new_n606), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n488), .A2(new_n561), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n602), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n621), .A2(KEYINPUT12), .A3(new_n374), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT12), .B1(new_n621), .B2(new_n374), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n618), .B1(new_n619), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n621), .A2(new_n374), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT12), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n621), .A2(KEYINPUT12), .A3(new_n374), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n608), .A2(new_n630), .A3(KEYINPUT86), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n625), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n617), .B1(new_n632), .B2(new_n616), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n594), .B1(new_n633), .B2(G469), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n608), .A2(new_n630), .A3(new_n615), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(KEYINPUT87), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT87), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n608), .A2(new_n630), .A3(new_n637), .A4(new_n615), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n611), .A2(new_n616), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n640), .A2(new_n593), .A3(new_n234), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n592), .B1(new_n634), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n485), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n573), .B1(new_n555), .B2(new_n571), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n585), .A2(new_n586), .A3(new_n575), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT95), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n484), .A2(new_n590), .A3(new_n642), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT103), .B(G101), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G3));
  NAND2_X1  g464(.A1(new_n476), .A2(new_n234), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(G472), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n482), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n619), .A2(new_n624), .A3(new_n618), .ZN(new_n654));
  AOI21_X1  g468(.A(KEYINPUT86), .B1(new_n608), .B2(new_n630), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n616), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n617), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n656), .A2(G469), .A3(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n594), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n641), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n237), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(KEYINPUT80), .A3(new_n235), .ZN(new_n662));
  INV_X1    g476(.A(new_n243), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n663), .B1(new_n237), .B2(new_n239), .ZN(new_n664));
  INV_X1    g478(.A(new_n246), .ZN(new_n665));
  AOI22_X1  g479(.A1(new_n662), .A2(new_n664), .B1(new_n233), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n660), .A2(new_n591), .A3(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n653), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n292), .A2(new_n318), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT104), .B(G478), .ZN(new_n670));
  OAI21_X1  g484(.A(KEYINPUT105), .B1(new_n348), .B2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n347), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n344), .B1(new_n332), .B2(new_n340), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n234), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n675));
  INV_X1    g489(.A(new_n670), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(KEYINPUT33), .B1(new_n672), .B2(new_n673), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT33), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n346), .A2(new_n679), .A3(new_n347), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n349), .A2(G902), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n671), .A2(new_n677), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n669), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n361), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n668), .A2(new_n646), .A3(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT34), .B(G104), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G6));
  NOR2_X1   g504(.A1(new_n354), .A2(new_n643), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n691), .A2(new_n292), .A3(new_n318), .A4(new_n361), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n644), .B2(new_n645), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n668), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT35), .B(G107), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G9));
  NOR2_X1   g510(.A1(new_n229), .A2(KEYINPUT36), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n220), .ZN(new_n698));
  AOI22_X1  g512(.A1(new_n662), .A2(new_n664), .B1(new_n665), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n362), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n700), .A2(new_n482), .A3(new_n652), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n590), .A2(new_n701), .A3(new_n647), .A4(new_n642), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT37), .B(G110), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G12));
  OR2_X1    g518(.A1(new_n359), .A2(G900), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n356), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NOR4_X1   g521(.A1(new_n699), .A2(new_n669), .A3(new_n354), .A4(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n481), .A2(new_n483), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n708), .A2(new_n709), .A3(new_n646), .A4(new_n642), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G128), .ZN(G30));
  NAND2_X1  g525(.A1(new_n660), .A2(new_n591), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n706), .B(KEYINPUT39), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  OR3_X1    g528(.A1(new_n712), .A2(KEYINPUT40), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n445), .B1(new_n468), .B2(new_n450), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n449), .A2(new_n450), .A3(new_n445), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT106), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n716), .A2(new_n721), .A3(new_n718), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n720), .A2(new_n234), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(G472), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n476), .A2(new_n480), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n483), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT40), .B1(new_n712), .B2(new_n714), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n715), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT38), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n729), .B1(new_n574), .B2(new_n587), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n644), .A2(KEYINPUT38), .A3(new_n645), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n669), .A2(new_n691), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n698), .A2(new_n665), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n733), .B1(new_n238), .B2(new_n244), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n730), .A2(new_n731), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n728), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n251), .ZN(G45));
  NAND3_X1  g552(.A1(new_n669), .A2(new_n684), .A3(new_n706), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n699), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n709), .A2(new_n646), .A3(new_n740), .A4(new_n642), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G146), .ZN(G48));
  AOI21_X1  g556(.A(new_n247), .B1(new_n481), .B2(new_n483), .ZN(new_n743));
  INV_X1    g557(.A(new_n641), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n593), .B1(new_n640), .B2(new_n234), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n744), .A2(new_n745), .A3(new_n592), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n743), .A2(new_n646), .A3(new_n687), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(KEYINPUT41), .B(G113), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G15));
  NAND3_X1  g563(.A1(new_n743), .A2(new_n693), .A3(new_n746), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G116), .ZN(G18));
  NAND4_X1  g565(.A1(new_n709), .A2(new_n646), .A3(new_n700), .A4(new_n746), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G119), .ZN(G21));
  AND2_X1   g567(.A1(new_n471), .A2(new_n474), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n445), .B1(new_n451), .B2(new_n458), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n478), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(G472), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n758), .B1(new_n476), .B2(new_n234), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n757), .A2(new_n759), .A3(new_n247), .ZN(new_n760));
  NOR4_X1   g574(.A1(new_n744), .A2(new_n745), .A3(new_n592), .A4(new_n686), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n732), .B1(new_n644), .B2(new_n645), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G122), .ZN(G24));
  AOI211_X1 g578(.A(new_n707), .B(new_n683), .C1(new_n292), .C2(new_n318), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n471), .A2(new_n474), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n477), .B1(new_n766), .B2(new_n755), .ZN(new_n767));
  AND4_X1   g581(.A1(new_n652), .A2(new_n734), .A3(new_n765), .A4(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n646), .A3(new_n746), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G125), .ZN(G27));
  NOR3_X1   g584(.A1(new_n574), .A2(new_n587), .A3(new_n643), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n743), .A2(new_n771), .A3(new_n642), .A4(new_n765), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT42), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n644), .A2(new_n485), .A3(new_n645), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n712), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n776), .A2(KEYINPUT42), .A3(new_n743), .A4(new_n765), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G131), .ZN(G33));
  INV_X1    g593(.A(new_n669), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n353), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n707), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n776), .A2(new_n743), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  NAND2_X1  g598(.A1(new_n633), .A2(KEYINPUT45), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(KEYINPUT107), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT107), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n633), .A2(new_n787), .A3(KEYINPUT45), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(G469), .B1(new_n633), .B2(KEYINPUT45), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(KEYINPUT46), .A3(new_n659), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT46), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n790), .B1(new_n786), .B2(new_n788), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n794), .B1(new_n795), .B2(new_n594), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n793), .A2(new_n641), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n591), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n798), .A2(new_n714), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT43), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n780), .A2(KEYINPUT108), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT108), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n683), .B1(new_n669), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n800), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n669), .A2(KEYINPUT43), .A3(new_n683), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT109), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT109), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n808), .B1(new_n804), .B2(new_n805), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n699), .B1(new_n652), .B2(new_n482), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n807), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT44), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n807), .A2(KEYINPUT44), .A3(new_n809), .A4(new_n810), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n799), .A2(new_n771), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G137), .ZN(G39));
  INV_X1    g630(.A(KEYINPUT47), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n798), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n797), .A2(KEYINPUT47), .A3(new_n591), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n709), .A2(new_n666), .A3(new_n739), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(new_n771), .A3(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G140), .ZN(G42));
  NAND2_X1  g637(.A1(new_n801), .A2(new_n803), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n824), .A2(new_n592), .A3(new_n643), .A4(new_n247), .ZN(new_n825));
  INV_X1    g639(.A(new_n726), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n744), .A2(new_n745), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT49), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n730), .A2(new_n731), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n825), .A2(new_n826), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n778), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n686), .B1(new_n781), .B2(new_n685), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n668), .A2(new_n590), .A3(new_n647), .A4(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n648), .A2(new_n833), .A3(new_n702), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT111), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n642), .A2(new_n485), .A3(new_n644), .A4(new_n645), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n652), .A2(new_n765), .A3(new_n734), .A4(new_n767), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n776), .A2(new_n768), .A3(KEYINPUT111), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n353), .A2(new_n707), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n292), .A3(new_n318), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT110), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT110), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n840), .A2(new_n292), .A3(new_n318), .A4(new_n843), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n842), .A2(new_n734), .A3(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n771), .A2(new_n845), .A3(new_n709), .A4(new_n642), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n838), .A2(new_n839), .A3(new_n783), .A4(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n747), .A2(new_n750), .A3(new_n763), .A4(new_n752), .ZN(new_n848));
  NOR4_X1   g662(.A1(new_n831), .A2(new_n834), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n734), .A2(new_n707), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n726), .A2(new_n642), .A3(new_n762), .A4(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n851), .A2(new_n769), .A3(new_n710), .A4(new_n741), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT52), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n710), .A2(new_n741), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT52), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n854), .A2(new_n855), .A3(new_n769), .A4(new_n851), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT53), .B1(new_n849), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT114), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n848), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n848), .A2(new_n860), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n853), .B(new_n856), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n847), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n648), .A2(new_n833), .A3(new_n702), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n864), .A2(new_n865), .A3(KEYINPUT53), .A4(new_n778), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n859), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n858), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n847), .B1(new_n774), .B2(new_n777), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n834), .A2(new_n848), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n869), .A2(new_n853), .A3(new_n856), .A4(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT112), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT112), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n871), .A2(new_n875), .A3(new_n872), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT113), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n870), .A2(new_n778), .A3(new_n864), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n853), .A2(new_n856), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n877), .B1(new_n880), .B2(KEYINPUT53), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n871), .A2(KEYINPUT113), .A3(new_n872), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n874), .B(new_n876), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n868), .B1(new_n883), .B2(KEYINPUT54), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n827), .A2(new_n591), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(new_n775), .ZN(new_n886));
  INV_X1    g700(.A(new_n356), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n806), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n743), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT48), .Z(new_n891));
  NAND3_X1  g705(.A1(new_n806), .A2(new_n887), .A3(new_n760), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n892), .A2(new_n588), .A3(new_n885), .ZN(new_n893));
  INV_X1    g707(.A(G952), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n893), .A2(new_n894), .A3(G953), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n247), .A2(new_n356), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n826), .A2(new_n886), .A3(new_n896), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n891), .B(new_n895), .C1(new_n685), .C2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n827), .A2(new_n592), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n818), .A2(new_n819), .A3(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n806), .A2(new_n887), .A3(new_n760), .A4(new_n771), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT115), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n780), .A2(new_n683), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n652), .A2(new_n734), .A3(new_n767), .ZN(new_n906));
  OAI22_X1  g720(.A1(new_n897), .A2(new_n905), .B1(new_n888), .B2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT50), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n746), .A2(new_n643), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT117), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n909), .A2(KEYINPUT117), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n912), .A2(new_n913), .A3(new_n829), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n908), .B1(new_n914), .B2(new_n892), .ZN(new_n915));
  INV_X1    g729(.A(new_n892), .ZN(new_n916));
  AOI22_X1  g730(.A1(new_n910), .A2(new_n911), .B1(new_n731), .B2(new_n730), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n916), .A2(KEYINPUT50), .A3(new_n917), .A4(new_n913), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n907), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT51), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n899), .B1(new_n904), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n901), .A2(new_n903), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n922), .A2(KEYINPUT118), .A3(KEYINPUT51), .A4(new_n919), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n898), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT51), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT116), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n919), .B1(new_n904), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n922), .A2(KEYINPUT116), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n884), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(G952), .A2(G953), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n830), .B1(new_n931), .B2(new_n932), .ZN(G75));
  NOR2_X1   g747(.A1(new_n225), .A2(G952), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n863), .ZN(new_n936));
  INV_X1    g750(.A(new_n866), .ZN(new_n937));
  AOI22_X1  g751(.A1(new_n936), .A2(new_n937), .B1(new_n871), .B2(new_n872), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n938), .A2(new_n234), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT56), .B1(new_n939), .B2(new_n573), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n577), .B1(new_n583), .B2(new_n584), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(new_n576), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT55), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n935), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n940), .B2(new_n943), .ZN(G51));
  OAI21_X1  g759(.A(KEYINPUT119), .B1(new_n858), .B2(new_n867), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n831), .A2(new_n872), .A3(new_n834), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n848), .B(new_n860), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n857), .A2(new_n947), .A3(new_n864), .A4(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT119), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n873), .A2(new_n949), .A3(new_n950), .A4(new_n859), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n946), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT120), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n938), .B2(new_n859), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n873), .A2(new_n949), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n955), .A2(KEYINPUT120), .A3(KEYINPUT54), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n952), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n594), .B(KEYINPUT57), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n640), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n939), .A2(new_n795), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n934), .B1(new_n960), .B2(new_n961), .ZN(G54));
  NAND4_X1  g776(.A1(new_n955), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n963));
  OR3_X1    g777(.A1(new_n963), .A2(KEYINPUT121), .A3(new_n311), .ZN(new_n964));
  OAI21_X1  g778(.A(KEYINPUT121), .B1(new_n963), .B2(new_n311), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n934), .B1(new_n963), .B2(new_n311), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(G60));
  INV_X1    g781(.A(new_n681), .ZN(new_n968));
  XNOR2_X1  g782(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n349), .A2(new_n234), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n968), .B1(new_n884), .B2(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n968), .A2(new_n971), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n934), .B1(new_n957), .B2(new_n973), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n972), .A2(new_n974), .ZN(G63));
  OR3_X1    g789(.A1(new_n343), .A2(new_n234), .A3(KEYINPUT60), .ZN(new_n976));
  OAI21_X1  g790(.A(KEYINPUT60), .B1(new_n343), .B2(new_n234), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n245), .B1(new_n938), .B2(new_n978), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n955), .A2(new_n698), .A3(new_n976), .A4(new_n977), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n979), .A2(new_n980), .A3(new_n935), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g796(.A(G953), .B1(new_n357), .B2(new_n493), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(new_n870), .B2(G953), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n941), .B1(G898), .B2(new_n225), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT123), .Z(new_n986));
  XNOR2_X1  g800(.A(new_n984), .B(new_n986), .ZN(G69));
  NAND2_X1  g801(.A1(new_n854), .A2(new_n769), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n989), .B(KEYINPUT62), .C1(new_n736), .C2(new_n728), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT62), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n991), .B1(new_n988), .B2(new_n737), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n822), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n781), .A2(new_n685), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n995), .A2(new_n642), .A3(new_n713), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n996), .A2(new_n775), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n815), .B1(new_n889), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n225), .B1(new_n994), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n400), .B1(new_n421), .B2(new_n431), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n305), .A2(new_n307), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n225), .B1(G227), .B2(G900), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  AND2_X1   g819(.A1(new_n743), .A2(new_n762), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n797), .A2(new_n591), .A3(new_n713), .A4(new_n1006), .ZN(new_n1007));
  AND4_X1   g821(.A1(new_n778), .A2(new_n989), .A3(new_n783), .A4(new_n1007), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n822), .A2(new_n1008), .A3(new_n225), .A4(new_n815), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1002), .B1(G900), .B2(G953), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1003), .A2(new_n1005), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(KEYINPUT124), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT124), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1009), .A2(new_n1014), .A3(new_n1010), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1003), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT125), .ZN(new_n1017));
  AND3_X1   g831(.A1(new_n1016), .A2(new_n1017), .A3(new_n1004), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1017), .B1(new_n1016), .B2(new_n1004), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1012), .B1(new_n1018), .B2(new_n1019), .ZN(G72));
  NAND3_X1  g834(.A1(new_n432), .A2(new_n444), .A3(new_n440), .ZN(new_n1021));
  XNOR2_X1  g835(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n758), .A2(new_n234), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  AND4_X1   g838(.A1(new_n716), .A2(new_n883), .A3(new_n1021), .A4(new_n1024), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n994), .A2(new_n998), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(new_n870), .ZN(new_n1027));
  XOR2_X1   g841(.A(new_n1024), .B(KEYINPUT127), .Z(new_n1028));
  AOI21_X1  g842(.A(new_n716), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n822), .A2(new_n1008), .A3(new_n815), .A4(new_n870), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1021), .B1(new_n1030), .B2(new_n1028), .ZN(new_n1031));
  NOR4_X1   g845(.A1(new_n1025), .A2(new_n1029), .A3(new_n934), .A4(new_n1031), .ZN(G57));
endmodule


