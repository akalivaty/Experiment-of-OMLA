

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U552 ( .A(n747), .B(KEYINPUT93), .ZN(n714) );
  NAND2_X1 U553 ( .A1(n716), .A2(n715), .ZN(n718) );
  NOR2_X1 U554 ( .A1(n626), .A2(n533), .ZN(n644) );
  INV_X1 U555 ( .A(KEYINPUT96), .ZN(n717) );
  XNOR2_X1 U556 ( .A(n718), .B(n717), .ZN(n728) );
  XNOR2_X1 U557 ( .A(KEYINPUT29), .B(KEYINPUT97), .ZN(n736) );
  XOR2_X1 U558 ( .A(n678), .B(KEYINPUT89), .Z(n704) );
  NOR2_X1 U559 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  NOR2_X1 U560 ( .A1(G651), .A2(n626), .ZN(n641) );
  AND2_X2 U561 ( .A1(n524), .A2(G2104), .ZN(n874) );
  NOR2_X1 U562 ( .A1(G651), .A2(G543), .ZN(n648) );
  INV_X1 U563 ( .A(G2105), .ZN(n524) );
  NAND2_X1 U564 ( .A1(G101), .A2(n874), .ZN(n518) );
  XNOR2_X1 U565 ( .A(n518), .B(KEYINPUT23), .ZN(n519) );
  XNOR2_X1 U566 ( .A(n519), .B(KEYINPUT65), .ZN(n522) );
  NAND2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  XOR2_X1 U568 ( .A(KEYINPUT66), .B(n520), .Z(n879) );
  NAND2_X1 U569 ( .A1(G113), .A2(n879), .ZN(n521) );
  NAND2_X1 U570 ( .A1(n522), .A2(n521), .ZN(n528) );
  XOR2_X1 U571 ( .A(KEYINPUT17), .B(n523), .Z(n872) );
  NAND2_X1 U572 ( .A1(G137), .A2(n872), .ZN(n526) );
  NOR2_X1 U573 ( .A1(G2104), .A2(n524), .ZN(n878) );
  NAND2_X1 U574 ( .A1(G125), .A2(n878), .ZN(n525) );
  NAND2_X1 U575 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U576 ( .A1(n528), .A2(n527), .ZN(G160) );
  XNOR2_X1 U577 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  INV_X1 U578 ( .A(G651), .ZN(n533) );
  NOR2_X1 U579 ( .A1(G543), .A2(n533), .ZN(n530) );
  XNOR2_X1 U580 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n529) );
  XNOR2_X1 U581 ( .A(n530), .B(n529), .ZN(n640) );
  NAND2_X1 U582 ( .A1(G64), .A2(n640), .ZN(n532) );
  XOR2_X1 U583 ( .A(KEYINPUT0), .B(G543), .Z(n626) );
  NAND2_X1 U584 ( .A1(G52), .A2(n641), .ZN(n531) );
  NAND2_X1 U585 ( .A1(n532), .A2(n531), .ZN(n538) );
  NAND2_X1 U586 ( .A1(G90), .A2(n648), .ZN(n535) );
  NAND2_X1 U587 ( .A1(G77), .A2(n644), .ZN(n534) );
  NAND2_X1 U588 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U589 ( .A(KEYINPUT9), .B(n536), .Z(n537) );
  NOR2_X1 U590 ( .A1(n538), .A2(n537), .ZN(G171) );
  AND2_X1 U591 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U592 ( .A1(n878), .A2(G123), .ZN(n540) );
  XNOR2_X1 U593 ( .A(KEYINPUT76), .B(KEYINPUT18), .ZN(n539) );
  XNOR2_X1 U594 ( .A(n540), .B(n539), .ZN(n547) );
  NAND2_X1 U595 ( .A1(G99), .A2(n874), .ZN(n542) );
  NAND2_X1 U596 ( .A1(G111), .A2(n879), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n542), .A2(n541), .ZN(n545) );
  NAND2_X1 U598 ( .A1(G135), .A2(n872), .ZN(n543) );
  XNOR2_X1 U599 ( .A(KEYINPUT77), .B(n543), .ZN(n544) );
  NOR2_X1 U600 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n547), .A2(n546), .ZN(n935) );
  XNOR2_X1 U602 ( .A(G2096), .B(n935), .ZN(n548) );
  OR2_X1 U603 ( .A1(G2100), .A2(n548), .ZN(G156) );
  INV_X1 U604 ( .A(G132), .ZN(G219) );
  INV_X1 U605 ( .A(G82), .ZN(G220) );
  INV_X1 U606 ( .A(G57), .ZN(G237) );
  NAND2_X1 U607 ( .A1(G102), .A2(n874), .ZN(n549) );
  XNOR2_X1 U608 ( .A(n549), .B(KEYINPUT86), .ZN(n552) );
  NAND2_X1 U609 ( .A1(n872), .A2(G138), .ZN(n550) );
  XOR2_X1 U610 ( .A(KEYINPUT87), .B(n550), .Z(n551) );
  NAND2_X1 U611 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U612 ( .A1(G126), .A2(n878), .ZN(n554) );
  NAND2_X1 U613 ( .A1(G114), .A2(n879), .ZN(n553) );
  NAND2_X1 U614 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U615 ( .A1(n556), .A2(n555), .ZN(G164) );
  NAND2_X1 U616 ( .A1(n648), .A2(G89), .ZN(n557) );
  XNOR2_X1 U617 ( .A(n557), .B(KEYINPUT4), .ZN(n559) );
  NAND2_X1 U618 ( .A1(G76), .A2(n644), .ZN(n558) );
  NAND2_X1 U619 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U620 ( .A(n560), .B(KEYINPUT5), .ZN(n566) );
  XNOR2_X1 U621 ( .A(KEYINPUT6), .B(KEYINPUT73), .ZN(n564) );
  NAND2_X1 U622 ( .A1(G63), .A2(n640), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G51), .A2(n641), .ZN(n561) );
  NAND2_X1 U624 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U625 ( .A(n564), .B(n563), .ZN(n565) );
  NAND2_X1 U626 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U627 ( .A(KEYINPUT7), .B(n567), .ZN(G168) );
  XOR2_X1 U628 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U629 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U630 ( .A(n568), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U631 ( .A(G223), .ZN(n817) );
  NAND2_X1 U632 ( .A1(n817), .A2(G567), .ZN(n569) );
  XNOR2_X1 U633 ( .A(n569), .B(KEYINPUT11), .ZN(n570) );
  XNOR2_X1 U634 ( .A(KEYINPUT69), .B(n570), .ZN(G234) );
  NAND2_X1 U635 ( .A1(n640), .A2(G56), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(KEYINPUT14), .ZN(n573) );
  NAND2_X1 U637 ( .A1(G43), .A2(n641), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n581) );
  NAND2_X1 U639 ( .A1(G81), .A2(n648), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(KEYINPUT12), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(KEYINPUT70), .ZN(n577) );
  NAND2_X1 U642 ( .A1(G68), .A2(n644), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(KEYINPUT13), .B(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(KEYINPUT71), .B(n579), .ZN(n580) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n967) );
  NAND2_X1 U647 ( .A1(n967), .A2(G860), .ZN(G153) );
  INV_X1 U648 ( .A(G171), .ZN(G301) );
  NAND2_X1 U649 ( .A1(G868), .A2(G301), .ZN(n591) );
  NAND2_X1 U650 ( .A1(G79), .A2(n644), .ZN(n588) );
  NAND2_X1 U651 ( .A1(G66), .A2(n640), .ZN(n583) );
  NAND2_X1 U652 ( .A1(G54), .A2(n641), .ZN(n582) );
  NAND2_X1 U653 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n648), .A2(G92), .ZN(n584) );
  XOR2_X1 U655 ( .A(KEYINPUT72), .B(n584), .Z(n585) );
  NOR2_X1 U656 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U657 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U658 ( .A(n589), .B(KEYINPUT15), .ZN(n966) );
  OR2_X1 U659 ( .A1(n966), .A2(G868), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n591), .A2(n590), .ZN(G284) );
  NAND2_X1 U661 ( .A1(G65), .A2(n640), .ZN(n593) );
  NAND2_X1 U662 ( .A1(G53), .A2(n641), .ZN(n592) );
  NAND2_X1 U663 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U664 ( .A1(G91), .A2(n648), .ZN(n595) );
  NAND2_X1 U665 ( .A1(G78), .A2(n644), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U667 ( .A1(n597), .A2(n596), .ZN(n972) );
  INV_X1 U668 ( .A(n972), .ZN(G299) );
  INV_X1 U669 ( .A(G868), .ZN(n651) );
  NOR2_X1 U670 ( .A1(G286), .A2(n651), .ZN(n598) );
  XNOR2_X1 U671 ( .A(n598), .B(KEYINPUT74), .ZN(n600) );
  NOR2_X1 U672 ( .A1(G299), .A2(G868), .ZN(n599) );
  NOR2_X1 U673 ( .A1(n600), .A2(n599), .ZN(G297) );
  INV_X1 U674 ( .A(G860), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n601), .A2(G559), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n602), .A2(n966), .ZN(n603) );
  XNOR2_X1 U677 ( .A(n603), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U678 ( .A1(n967), .A2(n651), .ZN(n604) );
  XNOR2_X1 U679 ( .A(KEYINPUT75), .B(n604), .ZN(n607) );
  NAND2_X1 U680 ( .A1(G868), .A2(n966), .ZN(n605) );
  NOR2_X1 U681 ( .A1(G559), .A2(n605), .ZN(n606) );
  NOR2_X1 U682 ( .A1(n607), .A2(n606), .ZN(G282) );
  NAND2_X1 U683 ( .A1(G67), .A2(n640), .ZN(n609) );
  NAND2_X1 U684 ( .A1(G55), .A2(n641), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U686 ( .A1(G93), .A2(n648), .ZN(n610) );
  XNOR2_X1 U687 ( .A(KEYINPUT79), .B(n610), .ZN(n611) );
  NOR2_X1 U688 ( .A1(n612), .A2(n611), .ZN(n614) );
  NAND2_X1 U689 ( .A1(n644), .A2(G80), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n653) );
  NAND2_X1 U691 ( .A1(G559), .A2(n966), .ZN(n615) );
  XOR2_X1 U692 ( .A(n967), .B(n615), .Z(n659) );
  NOR2_X1 U693 ( .A1(G860), .A2(n659), .ZN(n617) );
  XNOR2_X1 U694 ( .A(KEYINPUT78), .B(KEYINPUT80), .ZN(n616) );
  XNOR2_X1 U695 ( .A(n617), .B(n616), .ZN(n618) );
  XOR2_X1 U696 ( .A(n653), .B(n618), .Z(G145) );
  NAND2_X1 U697 ( .A1(G62), .A2(n640), .ZN(n620) );
  NAND2_X1 U698 ( .A1(G50), .A2(n641), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n623) );
  NAND2_X1 U700 ( .A1(n648), .A2(G88), .ZN(n621) );
  XOR2_X1 U701 ( .A(KEYINPUT82), .B(n621), .Z(n622) );
  NOR2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n644), .A2(G75), .ZN(n624) );
  NAND2_X1 U704 ( .A1(n625), .A2(n624), .ZN(G303) );
  INV_X1 U705 ( .A(G303), .ZN(G166) );
  NAND2_X1 U706 ( .A1(n626), .A2(G87), .ZN(n631) );
  NAND2_X1 U707 ( .A1(G49), .A2(n641), .ZN(n628) );
  NAND2_X1 U708 ( .A1(G74), .A2(G651), .ZN(n627) );
  NAND2_X1 U709 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U710 ( .A1(n640), .A2(n629), .ZN(n630) );
  NAND2_X1 U711 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U712 ( .A(KEYINPUT81), .B(n632), .Z(G288) );
  NAND2_X1 U713 ( .A1(n648), .A2(G85), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n640), .A2(G60), .ZN(n633) );
  NAND2_X1 U715 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U716 ( .A1(G47), .A2(n641), .ZN(n636) );
  NAND2_X1 U717 ( .A1(G72), .A2(n644), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U720 ( .A(KEYINPUT68), .B(n639), .Z(G290) );
  NAND2_X1 U721 ( .A1(G61), .A2(n640), .ZN(n643) );
  NAND2_X1 U722 ( .A1(G48), .A2(n641), .ZN(n642) );
  NAND2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U724 ( .A1(n644), .A2(G73), .ZN(n645) );
  XOR2_X1 U725 ( .A(KEYINPUT2), .B(n645), .Z(n646) );
  NOR2_X1 U726 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U727 ( .A1(n648), .A2(G86), .ZN(n649) );
  NAND2_X1 U728 ( .A1(n650), .A2(n649), .ZN(G305) );
  AND2_X1 U729 ( .A1(n651), .A2(n653), .ZN(n652) );
  XNOR2_X1 U730 ( .A(n652), .B(KEYINPUT83), .ZN(n662) );
  XNOR2_X1 U731 ( .A(G166), .B(KEYINPUT19), .ZN(n658) );
  XNOR2_X1 U732 ( .A(n972), .B(n653), .ZN(n656) );
  XOR2_X1 U733 ( .A(G290), .B(G305), .Z(n654) );
  XNOR2_X1 U734 ( .A(G288), .B(n654), .ZN(n655) );
  XNOR2_X1 U735 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U736 ( .A(n658), .B(n657), .ZN(n843) );
  XNOR2_X1 U737 ( .A(n843), .B(n659), .ZN(n660) );
  NAND2_X1 U738 ( .A1(G868), .A2(n660), .ZN(n661) );
  NAND2_X1 U739 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U740 ( .A1(G2078), .A2(G2084), .ZN(n663) );
  XOR2_X1 U741 ( .A(KEYINPUT20), .B(n663), .Z(n664) );
  NAND2_X1 U742 ( .A1(G2090), .A2(n664), .ZN(n665) );
  XNOR2_X1 U743 ( .A(KEYINPUT21), .B(n665), .ZN(n666) );
  NAND2_X1 U744 ( .A1(n666), .A2(G2072), .ZN(n667) );
  XNOR2_X1 U745 ( .A(KEYINPUT84), .B(n667), .ZN(G158) );
  NAND2_X1 U746 ( .A1(G69), .A2(G120), .ZN(n668) );
  NOR2_X1 U747 ( .A1(G237), .A2(n668), .ZN(n669) );
  NAND2_X1 U748 ( .A1(G108), .A2(n669), .ZN(n906) );
  NAND2_X1 U749 ( .A1(G567), .A2(n906), .ZN(n670) );
  XNOR2_X1 U750 ( .A(n670), .B(KEYINPUT85), .ZN(n675) );
  NOR2_X1 U751 ( .A1(G220), .A2(G219), .ZN(n671) );
  XNOR2_X1 U752 ( .A(KEYINPUT22), .B(n671), .ZN(n672) );
  NAND2_X1 U753 ( .A1(n672), .A2(G96), .ZN(n673) );
  OR2_X1 U754 ( .A1(G218), .A2(n673), .ZN(n907) );
  AND2_X1 U755 ( .A1(G2106), .A2(n907), .ZN(n674) );
  NOR2_X1 U756 ( .A1(n675), .A2(n674), .ZN(G319) );
  INV_X1 U757 ( .A(G319), .ZN(n677) );
  NAND2_X1 U758 ( .A1(G661), .A2(G483), .ZN(n676) );
  NOR2_X1 U759 ( .A1(n677), .A2(n676), .ZN(n819) );
  NAND2_X1 U760 ( .A1(n819), .A2(G36), .ZN(G176) );
  NAND2_X1 U761 ( .A1(G160), .A2(G40), .ZN(n678) );
  NOR2_X1 U762 ( .A1(G164), .A2(G1384), .ZN(n705) );
  NOR2_X1 U763 ( .A1(n704), .A2(n705), .ZN(n813) );
  NAND2_X1 U764 ( .A1(G128), .A2(n878), .ZN(n680) );
  NAND2_X1 U765 ( .A1(G116), .A2(n879), .ZN(n679) );
  NAND2_X1 U766 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U767 ( .A(n681), .B(KEYINPUT35), .ZN(n686) );
  NAND2_X1 U768 ( .A1(G104), .A2(n874), .ZN(n683) );
  NAND2_X1 U769 ( .A1(G140), .A2(n872), .ZN(n682) );
  NAND2_X1 U770 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U771 ( .A(KEYINPUT34), .B(n684), .Z(n685) );
  NAND2_X1 U772 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U773 ( .A(n687), .B(KEYINPUT36), .Z(n887) );
  XNOR2_X1 U774 ( .A(G2067), .B(KEYINPUT37), .ZN(n808) );
  NOR2_X1 U775 ( .A1(n887), .A2(n808), .ZN(n955) );
  NAND2_X1 U776 ( .A1(n813), .A2(n955), .ZN(n806) );
  NAND2_X1 U777 ( .A1(G95), .A2(n874), .ZN(n689) );
  NAND2_X1 U778 ( .A1(G131), .A2(n872), .ZN(n688) );
  NAND2_X1 U779 ( .A1(n689), .A2(n688), .ZN(n693) );
  NAND2_X1 U780 ( .A1(G119), .A2(n878), .ZN(n691) );
  NAND2_X1 U781 ( .A1(G107), .A2(n879), .ZN(n690) );
  NAND2_X1 U782 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U783 ( .A1(n693), .A2(n692), .ZN(n868) );
  INV_X1 U784 ( .A(G1991), .ZN(n1000) );
  NOR2_X1 U785 ( .A1(n868), .A2(n1000), .ZN(n702) );
  NAND2_X1 U786 ( .A1(G129), .A2(n878), .ZN(n695) );
  NAND2_X1 U787 ( .A1(G117), .A2(n879), .ZN(n694) );
  NAND2_X1 U788 ( .A1(n695), .A2(n694), .ZN(n698) );
  NAND2_X1 U789 ( .A1(n874), .A2(G105), .ZN(n696) );
  XOR2_X1 U790 ( .A(KEYINPUT38), .B(n696), .Z(n697) );
  NOR2_X1 U791 ( .A1(n698), .A2(n697), .ZN(n700) );
  NAND2_X1 U792 ( .A1(n872), .A2(G141), .ZN(n699) );
  NAND2_X1 U793 ( .A1(n700), .A2(n699), .ZN(n855) );
  AND2_X1 U794 ( .A1(G1996), .A2(n855), .ZN(n701) );
  NOR2_X1 U795 ( .A1(n702), .A2(n701), .ZN(n940) );
  INV_X1 U796 ( .A(n813), .ZN(n796) );
  NOR2_X1 U797 ( .A1(n940), .A2(n796), .ZN(n803) );
  INV_X1 U798 ( .A(n803), .ZN(n703) );
  NAND2_X1 U799 ( .A1(n806), .A2(n703), .ZN(n793) );
  INV_X1 U800 ( .A(G1961), .ZN(n968) );
  XNOR2_X1 U801 ( .A(KEYINPUT91), .B(n704), .ZN(n706) );
  NAND2_X2 U802 ( .A1(n706), .A2(n705), .ZN(n747) );
  NAND2_X1 U803 ( .A1(n968), .A2(n747), .ZN(n708) );
  XNOR2_X1 U804 ( .A(KEYINPUT25), .B(G2078), .ZN(n1008) );
  NAND2_X1 U805 ( .A1(n714), .A2(n1008), .ZN(n707) );
  NAND2_X1 U806 ( .A1(n708), .A2(n707), .ZN(n743) );
  AND2_X1 U807 ( .A1(n743), .A2(G171), .ZN(n709) );
  XOR2_X1 U808 ( .A(KEYINPUT94), .B(n709), .Z(n739) );
  NAND2_X1 U809 ( .A1(n714), .A2(G2072), .ZN(n710) );
  XNOR2_X1 U810 ( .A(n710), .B(KEYINPUT27), .ZN(n712) );
  INV_X1 U811 ( .A(G1956), .ZN(n913) );
  NOR2_X1 U812 ( .A1(n913), .A2(n714), .ZN(n711) );
  NOR2_X1 U813 ( .A1(n712), .A2(n711), .ZN(n731) );
  NOR2_X1 U814 ( .A1(n731), .A2(n972), .ZN(n713) );
  XOR2_X1 U815 ( .A(n713), .B(KEYINPUT28), .Z(n735) );
  NAND2_X1 U816 ( .A1(G2067), .A2(n714), .ZN(n716) );
  NAND2_X1 U817 ( .A1(G1348), .A2(n747), .ZN(n715) );
  NAND2_X1 U818 ( .A1(n728), .A2(n966), .ZN(n727) );
  NAND2_X1 U819 ( .A1(n747), .A2(G1341), .ZN(n719) );
  XNOR2_X1 U820 ( .A(n719), .B(KEYINPUT95), .ZN(n724) );
  XNOR2_X1 U821 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n722) );
  INV_X1 U822 ( .A(n747), .ZN(n720) );
  NAND2_X1 U823 ( .A1(G1996), .A2(n720), .ZN(n721) );
  XOR2_X1 U824 ( .A(n722), .B(n721), .Z(n723) );
  NOR2_X1 U825 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U826 ( .A1(n967), .A2(n725), .ZN(n726) );
  NAND2_X1 U827 ( .A1(n727), .A2(n726), .ZN(n730) );
  OR2_X1 U828 ( .A1(n966), .A2(n728), .ZN(n729) );
  NAND2_X1 U829 ( .A1(n730), .A2(n729), .ZN(n733) );
  NAND2_X1 U830 ( .A1(n731), .A2(n972), .ZN(n732) );
  NAND2_X1 U831 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U832 ( .A1(n735), .A2(n734), .ZN(n737) );
  XNOR2_X1 U833 ( .A(n737), .B(n736), .ZN(n738) );
  NAND2_X1 U834 ( .A1(n739), .A2(n738), .ZN(n759) );
  NAND2_X1 U835 ( .A1(G8), .A2(n747), .ZN(n789) );
  NOR2_X1 U836 ( .A1(G1966), .A2(n789), .ZN(n762) );
  NOR2_X1 U837 ( .A1(G2084), .A2(n747), .ZN(n758) );
  NOR2_X1 U838 ( .A1(n762), .A2(n758), .ZN(n740) );
  NAND2_X1 U839 ( .A1(G8), .A2(n740), .ZN(n741) );
  XNOR2_X1 U840 ( .A(KEYINPUT30), .B(n741), .ZN(n742) );
  NOR2_X1 U841 ( .A1(G168), .A2(n742), .ZN(n745) );
  NOR2_X1 U842 ( .A1(G171), .A2(n743), .ZN(n744) );
  NOR2_X1 U843 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U844 ( .A(KEYINPUT31), .B(n746), .Z(n760) );
  NOR2_X1 U845 ( .A1(G1971), .A2(n789), .ZN(n749) );
  NOR2_X1 U846 ( .A1(G2090), .A2(n747), .ZN(n748) );
  NOR2_X1 U847 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U848 ( .A1(n750), .A2(G303), .ZN(n752) );
  AND2_X1 U849 ( .A1(n760), .A2(n752), .ZN(n751) );
  NAND2_X1 U850 ( .A1(n759), .A2(n751), .ZN(n756) );
  INV_X1 U851 ( .A(n752), .ZN(n753) );
  OR2_X1 U852 ( .A1(n753), .A2(G286), .ZN(n754) );
  AND2_X1 U853 ( .A1(G8), .A2(n754), .ZN(n755) );
  NAND2_X1 U854 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U855 ( .A(n757), .B(KEYINPUT32), .ZN(n766) );
  NAND2_X1 U856 ( .A1(G8), .A2(n758), .ZN(n764) );
  AND2_X1 U857 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U858 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U859 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U860 ( .A1(n766), .A2(n765), .ZN(n773) );
  NOR2_X1 U861 ( .A1(G2090), .A2(G303), .ZN(n767) );
  NAND2_X1 U862 ( .A1(G8), .A2(n767), .ZN(n768) );
  NAND2_X1 U863 ( .A1(n773), .A2(n768), .ZN(n769) );
  NAND2_X1 U864 ( .A1(n769), .A2(n789), .ZN(n785) );
  NOR2_X1 U865 ( .A1(G1976), .A2(G288), .ZN(n776) );
  NOR2_X1 U866 ( .A1(G1971), .A2(G303), .ZN(n770) );
  NOR2_X1 U867 ( .A1(n776), .A2(n770), .ZN(n982) );
  INV_X1 U868 ( .A(KEYINPUT33), .ZN(n771) );
  AND2_X1 U869 ( .A1(n982), .A2(n771), .ZN(n772) );
  NAND2_X1 U870 ( .A1(n773), .A2(n772), .ZN(n783) );
  NAND2_X1 U871 ( .A1(G1976), .A2(G288), .ZN(n981) );
  INV_X1 U872 ( .A(n981), .ZN(n774) );
  NOR2_X1 U873 ( .A1(n789), .A2(n774), .ZN(n775) );
  NOR2_X1 U874 ( .A1(KEYINPUT33), .A2(n775), .ZN(n781) );
  XOR2_X1 U875 ( .A(G1981), .B(G305), .Z(n978) );
  INV_X1 U876 ( .A(n978), .ZN(n779) );
  NAND2_X1 U877 ( .A1(n776), .A2(KEYINPUT33), .ZN(n777) );
  NOR2_X1 U878 ( .A1(n789), .A2(n777), .ZN(n778) );
  OR2_X1 U879 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U880 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U881 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U882 ( .A1(n785), .A2(n784), .ZN(n791) );
  NOR2_X1 U883 ( .A1(G1981), .A2(G305), .ZN(n786) );
  XOR2_X1 U884 ( .A(n786), .B(KEYINPUT24), .Z(n787) );
  XNOR2_X1 U885 ( .A(KEYINPUT92), .B(n787), .ZN(n788) );
  NOR2_X1 U886 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U887 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U888 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U889 ( .A(n794), .B(KEYINPUT98), .ZN(n799) );
  XOR2_X1 U890 ( .A(G1986), .B(G290), .Z(n795) );
  XNOR2_X1 U891 ( .A(KEYINPUT88), .B(n795), .ZN(n991) );
  NOR2_X1 U892 ( .A1(n796), .A2(n991), .ZN(n797) );
  XOR2_X1 U893 ( .A(KEYINPUT90), .B(n797), .Z(n798) );
  NAND2_X1 U894 ( .A1(n799), .A2(n798), .ZN(n815) );
  NOR2_X1 U895 ( .A1(G1996), .A2(n855), .ZN(n953) );
  NOR2_X1 U896 ( .A1(G1986), .A2(G290), .ZN(n801) );
  AND2_X1 U897 ( .A1(n1000), .A2(n868), .ZN(n800) );
  XOR2_X1 U898 ( .A(KEYINPUT99), .B(n800), .Z(n938) );
  NOR2_X1 U899 ( .A1(n801), .A2(n938), .ZN(n802) );
  NOR2_X1 U900 ( .A1(n803), .A2(n802), .ZN(n804) );
  NOR2_X1 U901 ( .A1(n953), .A2(n804), .ZN(n805) );
  XNOR2_X1 U902 ( .A(KEYINPUT39), .B(n805), .ZN(n807) );
  NAND2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n810) );
  AND2_X1 U904 ( .A1(n887), .A2(n808), .ZN(n809) );
  XOR2_X1 U905 ( .A(KEYINPUT100), .B(n809), .Z(n947) );
  NAND2_X1 U906 ( .A1(n810), .A2(n947), .ZN(n811) );
  XOR2_X1 U907 ( .A(KEYINPUT101), .B(n811), .Z(n812) );
  NAND2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U910 ( .A(n816), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n817), .ZN(G217) );
  AND2_X1 U912 ( .A1(G15), .A2(G2), .ZN(n818) );
  NAND2_X1 U913 ( .A1(G661), .A2(n818), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n820) );
  NAND2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n821) );
  XOR2_X1 U916 ( .A(KEYINPUT103), .B(n821), .Z(G188) );
  XOR2_X1 U917 ( .A(G96), .B(KEYINPUT104), .Z(G221) );
  XOR2_X1 U918 ( .A(KEYINPUT105), .B(G2084), .Z(n823) );
  XNOR2_X1 U919 ( .A(G2067), .B(G2078), .ZN(n822) );
  XNOR2_X1 U920 ( .A(n823), .B(n822), .ZN(n824) );
  XOR2_X1 U921 ( .A(n824), .B(G2100), .Z(n826) );
  XNOR2_X1 U922 ( .A(G2072), .B(G2090), .ZN(n825) );
  XNOR2_X1 U923 ( .A(n826), .B(n825), .ZN(n830) );
  XOR2_X1 U924 ( .A(G2096), .B(KEYINPUT43), .Z(n828) );
  XNOR2_X1 U925 ( .A(G2678), .B(KEYINPUT42), .ZN(n827) );
  XNOR2_X1 U926 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U927 ( .A(n830), .B(n829), .Z(G227) );
  XOR2_X1 U928 ( .A(G1976), .B(G1971), .Z(n832) );
  XNOR2_X1 U929 ( .A(G1966), .B(G1956), .ZN(n831) );
  XNOR2_X1 U930 ( .A(n832), .B(n831), .ZN(n842) );
  XOR2_X1 U931 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n834) );
  XNOR2_X1 U932 ( .A(G1996), .B(KEYINPUT41), .ZN(n833) );
  XNOR2_X1 U933 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U934 ( .A(G1981), .B(G1961), .Z(n836) );
  XNOR2_X1 U935 ( .A(G1991), .B(G1986), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U937 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U938 ( .A(KEYINPUT106), .B(G2474), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(G229) );
  XOR2_X1 U941 ( .A(n843), .B(G286), .Z(n845) );
  XNOR2_X1 U942 ( .A(n966), .B(G171), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U944 ( .A(n967), .B(n846), .Z(n847) );
  NOR2_X1 U945 ( .A1(G37), .A2(n847), .ZN(G397) );
  NAND2_X1 U946 ( .A1(G124), .A2(n878), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n848), .B(KEYINPUT44), .ZN(n850) );
  NAND2_X1 U948 ( .A1(n874), .A2(G100), .ZN(n849) );
  NAND2_X1 U949 ( .A1(n850), .A2(n849), .ZN(n854) );
  NAND2_X1 U950 ( .A1(G136), .A2(n872), .ZN(n852) );
  NAND2_X1 U951 ( .A1(G112), .A2(n879), .ZN(n851) );
  NAND2_X1 U952 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U953 ( .A1(n854), .A2(n853), .ZN(G162) );
  XOR2_X1 U954 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n857) );
  XOR2_X1 U955 ( .A(n855), .B(KEYINPUT111), .Z(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n935), .B(n858), .ZN(n860) );
  XNOR2_X1 U958 ( .A(G164), .B(G160), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n871) );
  NAND2_X1 U960 ( .A1(G130), .A2(n878), .ZN(n862) );
  NAND2_X1 U961 ( .A1(G118), .A2(n879), .ZN(n861) );
  NAND2_X1 U962 ( .A1(n862), .A2(n861), .ZN(n867) );
  NAND2_X1 U963 ( .A1(G106), .A2(n874), .ZN(n864) );
  NAND2_X1 U964 ( .A1(G142), .A2(n872), .ZN(n863) );
  NAND2_X1 U965 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U966 ( .A(n865), .B(KEYINPUT45), .Z(n866) );
  NOR2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n869) );
  XOR2_X1 U968 ( .A(n869), .B(n868), .Z(n870) );
  XOR2_X1 U969 ( .A(n871), .B(n870), .Z(n886) );
  NAND2_X1 U970 ( .A1(n872), .A2(G139), .ZN(n873) );
  XOR2_X1 U971 ( .A(KEYINPUT109), .B(n873), .Z(n876) );
  NAND2_X1 U972 ( .A1(n874), .A2(G103), .ZN(n875) );
  NAND2_X1 U973 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U974 ( .A(KEYINPUT110), .B(n877), .ZN(n884) );
  NAND2_X1 U975 ( .A1(G127), .A2(n878), .ZN(n881) );
  NAND2_X1 U976 ( .A1(G115), .A2(n879), .ZN(n880) );
  NAND2_X1 U977 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U978 ( .A(KEYINPUT47), .B(n882), .Z(n883) );
  NOR2_X1 U979 ( .A1(n884), .A2(n883), .ZN(n941) );
  XNOR2_X1 U980 ( .A(n941), .B(G162), .ZN(n885) );
  XNOR2_X1 U981 ( .A(n886), .B(n885), .ZN(n888) );
  XOR2_X1 U982 ( .A(n888), .B(n887), .Z(n889) );
  NOR2_X1 U983 ( .A1(G37), .A2(n889), .ZN(n890) );
  XNOR2_X1 U984 ( .A(KEYINPUT112), .B(n890), .ZN(G395) );
  XOR2_X1 U985 ( .A(KEYINPUT102), .B(G2446), .Z(n892) );
  XNOR2_X1 U986 ( .A(G2443), .B(G2454), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U988 ( .A(n893), .B(G2451), .Z(n895) );
  XNOR2_X1 U989 ( .A(G1341), .B(G1348), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n895), .B(n894), .ZN(n899) );
  XOR2_X1 U991 ( .A(G2435), .B(G2427), .Z(n897) );
  XNOR2_X1 U992 ( .A(G2430), .B(G2438), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U994 ( .A(n899), .B(n898), .Z(n900) );
  NAND2_X1 U995 ( .A1(G14), .A2(n900), .ZN(n908) );
  NAND2_X1 U996 ( .A1(G319), .A2(n908), .ZN(n903) );
  NOR2_X1 U997 ( .A1(G227), .A2(G229), .ZN(n901) );
  XNOR2_X1 U998 ( .A(KEYINPUT49), .B(n901), .ZN(n902) );
  NOR2_X1 U999 ( .A1(n903), .A2(n902), .ZN(n905) );
  NOR2_X1 U1000 ( .A1(G397), .A2(G395), .ZN(n904) );
  NAND2_X1 U1001 ( .A1(n905), .A2(n904), .ZN(G225) );
  XNOR2_X1 U1002 ( .A(KEYINPUT113), .B(G225), .ZN(G308) );
  INV_X1 U1004 ( .A(G120), .ZN(G236) );
  INV_X1 U1005 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1006 ( .A1(n907), .A2(n906), .ZN(G325) );
  INV_X1 U1007 ( .A(G325), .ZN(G261) );
  INV_X1 U1008 ( .A(G108), .ZN(G238) );
  INV_X1 U1009 ( .A(n908), .ZN(G401) );
  XNOR2_X1 U1010 ( .A(G1966), .B(G21), .ZN(n910) );
  XNOR2_X1 U1011 ( .A(G1961), .B(G5), .ZN(n909) );
  NOR2_X1 U1012 ( .A1(n910), .A2(n909), .ZN(n922) );
  XOR2_X1 U1013 ( .A(KEYINPUT126), .B(G4), .Z(n912) );
  XNOR2_X1 U1014 ( .A(G1348), .B(KEYINPUT59), .ZN(n911) );
  XNOR2_X1 U1015 ( .A(n912), .B(n911), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(G20), .B(n913), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(G1341), .B(G19), .ZN(n915) );
  XNOR2_X1 U1018 ( .A(G6), .B(G1981), .ZN(n914) );
  NOR2_X1 U1019 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1020 ( .A1(n917), .A2(n916), .ZN(n918) );
  NOR2_X1 U1021 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1022 ( .A(n920), .B(KEYINPUT60), .ZN(n921) );
  NAND2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n930) );
  XNOR2_X1 U1024 ( .A(G1971), .B(G22), .ZN(n924) );
  XNOR2_X1 U1025 ( .A(G23), .B(G1976), .ZN(n923) );
  NOR2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n927) );
  XNOR2_X1 U1027 ( .A(G1986), .B(KEYINPUT127), .ZN(n925) );
  XNOR2_X1 U1028 ( .A(n925), .B(G24), .ZN(n926) );
  NAND2_X1 U1029 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1030 ( .A(KEYINPUT58), .B(n928), .ZN(n929) );
  NOR2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1032 ( .A(KEYINPUT61), .B(n931), .ZN(n933) );
  INV_X1 U1033 ( .A(G16), .ZN(n932) );
  NAND2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1035 ( .A1(n934), .A2(G11), .ZN(n965) );
  XNOR2_X1 U1036 ( .A(G160), .B(G2084), .ZN(n936) );
  NAND2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n950) );
  XOR2_X1 U1040 ( .A(G2072), .B(n941), .Z(n943) );
  XOR2_X1 U1041 ( .A(G164), .B(G2078), .Z(n942) );
  NOR2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n946) );
  XOR2_X1 U1043 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n944) );
  XNOR2_X1 U1044 ( .A(KEYINPUT50), .B(n944), .ZN(n945) );
  XNOR2_X1 U1045 ( .A(n946), .B(n945), .ZN(n948) );
  NAND2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n958) );
  XOR2_X1 U1048 ( .A(G2090), .B(G162), .Z(n951) );
  XNOR2_X1 U1049 ( .A(KEYINPUT114), .B(n951), .ZN(n952) );
  NOR2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(KEYINPUT51), .B(n954), .ZN(n956) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(KEYINPUT52), .B(n959), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(KEYINPUT117), .B(n960), .ZN(n961) );
  XOR2_X1 U1056 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n1018) );
  NAND2_X1 U1057 ( .A1(n961), .A2(n1018), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(G29), .A2(n962), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(KEYINPUT119), .B(n963), .ZN(n964) );
  NOR2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n996) );
  XNOR2_X1 U1061 ( .A(KEYINPUT56), .B(G16), .ZN(n994) );
  XNOR2_X1 U1062 ( .A(n966), .B(G1348), .ZN(n977) );
  XNOR2_X1 U1063 ( .A(n967), .B(G1341), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(G171), .B(KEYINPUT123), .ZN(n969) );
  XNOR2_X1 U1065 ( .A(n969), .B(n968), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n975) );
  XOR2_X1 U1067 ( .A(G1956), .B(n972), .Z(n973) );
  XNOR2_X1 U1068 ( .A(KEYINPUT124), .B(n973), .ZN(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n990) );
  XNOR2_X1 U1071 ( .A(G1966), .B(G168), .ZN(n979) );
  NAND2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(n980), .B(KEYINPUT57), .ZN(n988) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n985) );
  INV_X1 U1075 ( .A(G1971), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(G166), .A2(n983), .ZN(n984) );
  NOR2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1078 ( .A(KEYINPUT125), .B(n986), .Z(n987) );
  NAND2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n1021) );
  XNOR2_X1 U1084 ( .A(G2084), .B(G34), .ZN(n997) );
  XNOR2_X1 U1085 ( .A(n997), .B(KEYINPUT54), .ZN(n1016) );
  XNOR2_X1 U1086 ( .A(G2090), .B(G35), .ZN(n1013) );
  XNOR2_X1 U1087 ( .A(G1996), .B(G32), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(G33), .B(G2072), .ZN(n998) );
  NOR2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1007) );
  XNOR2_X1 U1090 ( .A(n1000), .B(G25), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(G28), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(n1002), .B(KEYINPUT120), .ZN(n1005) );
  XOR2_X1 U1093 ( .A(G2067), .B(KEYINPUT121), .Z(n1003) );
  XNOR2_X1 U1094 ( .A(G26), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1010) );
  XOR2_X1 U1097 ( .A(G27), .B(n1008), .Z(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(KEYINPUT53), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1101 ( .A(KEYINPUT122), .B(n1014), .Z(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(n1018), .B(n1017), .ZN(n1019) );
  NOR2_X1 U1104 ( .A1(G29), .A2(n1019), .ZN(n1020) );
  NOR2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1106 ( .A(n1022), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

