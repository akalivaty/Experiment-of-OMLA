//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n554, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n617, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1226, new_n1227,
    new_n1228;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT64), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT66), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI21_X1  g033(.A(KEYINPUT67), .B1(new_n453), .B2(G2106), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(G567), .B2(new_n456), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n453), .A2(KEYINPUT67), .A3(G2106), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(G137), .A3(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT68), .ZN(G160));
  NOR2_X1   g056(.A1(new_n476), .A2(new_n465), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n476), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(G162));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n465), .B2(G114), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n491), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G102), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(new_n465), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n490), .A2(new_n492), .A3(G2104), .A4(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n473), .A2(new_n475), .A3(G126), .A4(G2105), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n473), .A2(new_n475), .A3(G138), .A4(new_n465), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n464), .A2(new_n500), .A3(G138), .A4(new_n465), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n497), .B1(new_n499), .B2(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT70), .A3(G543), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n505), .A2(new_n507), .B1(KEYINPUT5), .B2(new_n504), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n512), .A2(G543), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n511), .A2(new_n517), .ZN(G166));
  INV_X1    g093(.A(new_n516), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G51), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n508), .A2(G89), .A3(new_n512), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n520), .A2(new_n521), .A3(new_n522), .A4(new_n524), .ZN(G286));
  INV_X1    g100(.A(G286), .ZN(G168));
  NAND2_X1  g101(.A1(new_n508), .A2(G64), .ZN(new_n527));
  NAND2_X1  g102(.A1(G77), .A2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n508), .A2(G90), .A3(new_n512), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n512), .A2(G52), .A3(G543), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n530), .A2(new_n533), .ZN(G301));
  INV_X1    g109(.A(G301), .ZN(G171));
  NAND2_X1  g110(.A1(G68), .A2(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n505), .A2(new_n507), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G56), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n536), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G651), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n537), .A2(G81), .A3(new_n538), .A4(new_n512), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT71), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n512), .A2(G43), .A3(G543), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n544), .B1(new_n543), .B2(new_n545), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n542), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(KEYINPUT72), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT72), .ZN(new_n550));
  OAI211_X1 g125(.A(new_n542), .B(new_n550), .C1(new_n546), .C2(new_n547), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(G188));
  INV_X1    g133(.A(KEYINPUT73), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT6), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n560), .A2(new_n562), .A3(G53), .A4(G543), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n508), .A2(G91), .A3(new_n512), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n508), .A2(G65), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n510), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n559), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n568), .B1(new_n539), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G651), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n573), .A2(KEYINPUT73), .A3(new_n565), .A4(new_n564), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n570), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G166), .ZN(G303));
  NAND2_X1  g151(.A1(new_n519), .A2(G49), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n578));
  INV_X1    g153(.A(G87), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n577), .B(new_n578), .C1(new_n579), .C2(new_n513), .ZN(G288));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  INV_X1    g156(.A(G48), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n513), .A2(new_n581), .B1(new_n582), .B2(new_n516), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n508), .A2(G61), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n510), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G305));
  INV_X1    g163(.A(G85), .ZN(new_n589));
  INV_X1    g164(.A(G47), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n513), .A2(new_n589), .B1(new_n590), .B2(new_n516), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT74), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(new_n510), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n508), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G54), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n598), .A2(new_n510), .B1(new_n599), .B2(new_n516), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI221_X1 g177(.A(KEYINPUT75), .B1(new_n599), .B2(new_n516), .C1(new_n598), .C2(new_n510), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n513), .B2(new_n605), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n508), .A2(new_n512), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n607), .A2(KEYINPUT10), .A3(G92), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n602), .A2(new_n603), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n597), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n597), .B1(new_n609), .B2(G868), .ZN(G321));
  NAND2_X1  g186(.A1(G286), .A2(G868), .ZN(new_n612));
  INV_X1    g187(.A(G299), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(G297));
  OAI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(G280));
  XOR2_X1   g190(.A(KEYINPUT76), .B(G559), .Z(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n609), .B1(G860), .B2(new_n617), .ZN(G148));
  NAND2_X1  g193(.A1(new_n609), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n482), .A2(G123), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n484), .A2(G135), .ZN(new_n624));
  OR2_X1    g199(.A1(G99), .A2(G2105), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n625), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n464), .A2(new_n468), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT77), .B(KEYINPUT12), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT13), .B(G2100), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n628), .A2(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(G2427), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT79), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2438), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(G2438), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n636), .A2(new_n640), .A3(new_n639), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(G14), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n650), .B2(new_n651), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n652), .A2(new_n654), .ZN(G401));
  XOR2_X1   g230(.A(G2067), .B(G2678), .Z(new_n656));
  XNOR2_X1  g231(.A(G2084), .B(G2090), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT80), .B(KEYINPUT18), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2072), .B(G2078), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(G2100), .Z(new_n663));
  NAND2_X1  g238(.A1(new_n656), .A2(new_n657), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n658), .A2(new_n664), .A3(KEYINPUT17), .ZN(new_n665));
  INV_X1    g240(.A(new_n659), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT81), .B(G2096), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n663), .B(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1981), .B(G1986), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  OR2_X1    g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT19), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n674), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n676), .A2(new_n677), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT83), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(new_n675), .B2(new_n679), .ZN(new_n689));
  NAND4_X1  g264(.A1(new_n682), .A2(new_n676), .A3(new_n677), .A4(new_n687), .ZN(new_n690));
  NAND4_X1  g265(.A1(new_n685), .A2(new_n686), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  NAND4_X1  g266(.A1(new_n689), .A2(new_n690), .A3(new_n684), .A4(new_n680), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(KEYINPUT83), .ZN(new_n693));
  INV_X1    g268(.A(G1991), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n694), .B1(new_n691), .B2(new_n693), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n673), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n697), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n699), .A2(G1996), .A3(new_n695), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n672), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n698), .A2(new_n700), .A3(new_n672), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n703), .ZN(new_n706));
  INV_X1    g281(.A(new_n704), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(new_n701), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n705), .A2(new_n708), .ZN(G229));
  NAND2_X1  g284(.A1(G162), .A2(G29), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G29), .B2(G35), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G2090), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT94), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n716), .A2(G26), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT91), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n465), .A2(G116), .ZN(new_n719));
  OAI21_X1  g294(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OR3_X1    g296(.A1(new_n719), .A2(new_n720), .A3(new_n718), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n721), .A2(new_n722), .B1(new_n482), .B2(G128), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n464), .A2(new_n465), .ZN(new_n724));
  INV_X1    g299(.A(G140), .ZN(new_n725));
  OR3_X1    g300(.A1(new_n724), .A2(KEYINPUT90), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(KEYINPUT90), .B1(new_n724), .B2(new_n725), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n723), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n717), .B1(new_n728), .B2(G29), .ZN(new_n729));
  MUX2_X1   g304(.A(new_n717), .B(new_n729), .S(KEYINPUT28), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G2067), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n715), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n716), .A2(G33), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n468), .A2(G103), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT25), .Z(new_n735));
  INV_X1    g310(.A(G139), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(new_n724), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(new_n465), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n733), .B1(new_n740), .B2(new_n716), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n482), .A2(G129), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n484), .A2(G141), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n468), .A2(G105), .ZN(new_n744));
  NAND3_X1  g319(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT26), .Z(new_n746));
  NAND4_X1  g321(.A1(new_n742), .A2(new_n743), .A3(new_n744), .A4(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G29), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G29), .B2(G32), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G1996), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n741), .A2(G2072), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n750), .B2(new_n751), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT31), .B(G11), .Z(new_n754));
  NOR2_X1   g329(.A1(new_n627), .A2(new_n716), .ZN(new_n755));
  INV_X1    g330(.A(G28), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(KEYINPUT30), .ZN(new_n757));
  AOI21_X1  g332(.A(G29), .B1(new_n756), .B2(KEYINPUT30), .ZN(new_n758));
  AOI211_X1 g333(.A(new_n754), .B(new_n755), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(G168), .A2(G16), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G16), .B2(G21), .ZN(new_n761));
  INV_X1    g336(.A(G1966), .ZN(new_n762));
  OAI221_X1 g337(.A(new_n759), .B1(new_n761), .B2(new_n762), .C1(G2072), .C2(new_n741), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n753), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n713), .ZN(new_n765));
  INV_X1    g340(.A(G2090), .ZN(new_n766));
  INV_X1    g341(.A(G2084), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT68), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n480), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(KEYINPUT24), .A2(G34), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT24), .ZN(new_n771));
  INV_X1    g346(.A(G34), .ZN(new_n772));
  AOI21_X1  g347(.A(G29), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n769), .A2(G29), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n765), .A2(new_n766), .B1(new_n767), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n761), .A2(new_n762), .ZN(new_n776));
  NOR2_X1   g351(.A1(G27), .A2(G29), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G164), .B2(G29), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n776), .B1(G2078), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G2078), .B2(new_n778), .ZN(new_n780));
  NOR2_X1   g355(.A1(G5), .A2(G16), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G171), .B2(G16), .ZN(new_n782));
  INV_X1    g357(.A(G1961), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n764), .A2(new_n775), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(G16), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(G4), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n609), .B2(new_n786), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1348), .ZN(new_n789));
  NOR3_X1   g364(.A1(new_n732), .A2(new_n785), .A3(new_n789), .ZN(new_n790));
  AND2_X1   g365(.A1(KEYINPUT85), .A2(G16), .ZN(new_n791));
  NOR2_X1   g366(.A1(KEYINPUT85), .A2(G16), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(G19), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n552), .B2(new_n793), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G1341), .Z(new_n796));
  NOR2_X1   g371(.A1(new_n774), .A2(new_n767), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT92), .Z(new_n798));
  INV_X1    g373(.A(new_n793), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G20), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT23), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n613), .B2(new_n786), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT95), .B(G1956), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n798), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n790), .A2(new_n796), .A3(new_n805), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(KEYINPUT96), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(KEYINPUT96), .ZN(new_n808));
  MUX2_X1   g383(.A(G23), .B(G288), .S(G16), .Z(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT33), .B(G1976), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT88), .B(KEYINPUT89), .Z(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n811), .A2(new_n813), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n799), .A2(G22), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G166), .B2(new_n799), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(G1971), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n786), .A2(G6), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n587), .B2(new_n786), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT32), .B(G1981), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT87), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n814), .A2(new_n815), .A3(new_n818), .A4(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT34), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n799), .A2(G24), .ZN(new_n826));
  INV_X1    g401(.A(G290), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(new_n799), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT86), .ZN(new_n829));
  INV_X1    g404(.A(G1986), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n830), .ZN(new_n832));
  NOR2_X1   g407(.A1(G25), .A2(G29), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n482), .A2(G119), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n484), .A2(G131), .ZN(new_n835));
  OR2_X1    g410(.A1(G95), .A2(G2105), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n836), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n833), .B1(new_n839), .B2(G29), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT35), .B(G1991), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT84), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n840), .B(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n831), .A2(new_n832), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(KEYINPUT36), .B1(new_n825), .B2(new_n844), .ZN(new_n845));
  OR3_X1    g420(.A1(new_n825), .A2(new_n844), .A3(KEYINPUT36), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n807), .A2(new_n808), .B1(new_n845), .B2(new_n846), .ZN(G311));
  XNOR2_X1  g422(.A(new_n806), .B(KEYINPUT96), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n845), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(G150));
  XNOR2_X1  g425(.A(KEYINPUT99), .B(G860), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n852), .A2(new_n510), .ZN(new_n853));
  INV_X1    g428(.A(G93), .ZN(new_n854));
  XNOR2_X1  g429(.A(KEYINPUT97), .B(G55), .ZN(new_n855));
  OAI22_X1  g430(.A1(new_n513), .A2(new_n854), .B1(new_n516), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n548), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n857), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n858), .B1(new_n552), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n609), .A2(G559), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT39), .ZN(new_n863));
  XNOR2_X1  g438(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n851), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(new_n864), .B2(new_n863), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n859), .A2(new_n851), .ZN(new_n867));
  XOR2_X1   g442(.A(KEYINPUT100), .B(KEYINPUT37), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n866), .A2(new_n869), .ZN(G145));
  NAND2_X1  g445(.A1(new_n769), .A2(new_n627), .ZN(new_n871));
  INV_X1    g446(.A(new_n627), .ZN(new_n872));
  NAND2_X1  g447(.A1(G160), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(G162), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n871), .A2(new_n873), .A3(G162), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n740), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n499), .A2(new_n501), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n495), .A2(new_n496), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n728), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n728), .A2(new_n882), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n883), .A2(new_n747), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n747), .B1(new_n883), .B2(new_n884), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n879), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n883), .A2(new_n884), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n748), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n890), .A2(new_n740), .A3(new_n885), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n482), .A2(G130), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n484), .A2(G142), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n465), .A2(G118), .ZN(new_n895));
  OAI21_X1  g470(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n893), .B(new_n894), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(new_n838), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(new_n631), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n878), .B1(new_n892), .B2(new_n901), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n888), .A2(new_n891), .A3(new_n900), .A4(new_n899), .ZN(new_n903));
  AOI21_X1  g478(.A(G37), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n886), .A2(new_n879), .A3(new_n887), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n740), .B1(new_n890), .B2(new_n885), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n899), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n899), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(new_n888), .A3(new_n891), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n909), .A3(new_n878), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT101), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT101), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n907), .A2(new_n912), .A3(new_n909), .A4(new_n878), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n904), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n914), .B(KEYINPUT40), .Z(G395));
  INV_X1    g490(.A(G868), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n859), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n613), .A2(new_n609), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n602), .A2(new_n603), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n608), .A2(new_n606), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(G299), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT41), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n918), .A2(new_n922), .A3(KEYINPUT41), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n860), .B(new_n619), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n609), .B(G299), .ZN(new_n930));
  AOI22_X1  g505(.A1(new_n929), .A2(KEYINPUT103), .B1(new_n930), .B2(new_n928), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(KEYINPUT103), .B2(new_n929), .ZN(new_n932));
  XNOR2_X1  g507(.A(G290), .B(G288), .ZN(new_n933));
  XNOR2_X1  g508(.A(G166), .B(new_n587), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n933), .B(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT42), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n932), .B(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n917), .B1(new_n937), .B2(new_n916), .ZN(G295));
  OAI21_X1  g513(.A(new_n917), .B1(new_n937), .B2(new_n916), .ZN(G331));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n530), .A2(new_n533), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n510), .B1(new_n527), .B2(new_n528), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n531), .A2(new_n532), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT104), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n941), .A2(G168), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n940), .B1(new_n530), .B2(new_n533), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n942), .A2(new_n943), .A3(KEYINPUT104), .ZN(new_n947));
  OAI21_X1  g522(.A(G286), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n857), .B1(new_n549), .B2(new_n551), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n945), .B(new_n948), .C1(new_n949), .C2(new_n858), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n945), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n860), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n951), .B1(new_n860), .B2(new_n952), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n930), .B(new_n950), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n547), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n550), .B1(new_n958), .B2(new_n542), .ZN(new_n959));
  INV_X1    g534(.A(new_n551), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n859), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n858), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(new_n952), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n950), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(new_n925), .A3(new_n926), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n935), .A2(new_n955), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G37), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n935), .B1(new_n965), .B2(new_n955), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT43), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n935), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n963), .A2(KEYINPUT105), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n860), .A2(new_n951), .A3(new_n952), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n927), .B1(new_n974), .B2(new_n950), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n950), .A2(new_n930), .A3(new_n963), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT106), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n950), .A2(new_n930), .A3(new_n963), .A4(KEYINPUT106), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n971), .B1(new_n975), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT43), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n981), .A2(new_n982), .A3(new_n967), .A4(new_n966), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n970), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n982), .B1(new_n968), .B2(new_n969), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n981), .A2(new_n967), .A3(new_n966), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n985), .B1(new_n986), .B2(new_n982), .ZN(new_n987));
  MUX2_X1   g562(.A(new_n984), .B(new_n987), .S(KEYINPUT44), .Z(G397));
  NAND3_X1  g563(.A1(new_n471), .A2(G40), .A3(new_n479), .ZN(new_n989));
  AOI21_X1  g564(.A(G1384), .B1(new_n880), .B2(new_n881), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n989), .A2(new_n990), .A3(KEYINPUT45), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n827), .A2(new_n830), .ZN(new_n992));
  XOR2_X1   g567(.A(new_n992), .B(KEYINPUT107), .Z(new_n993));
  XOR2_X1   g568(.A(new_n728), .B(G2067), .Z(new_n994));
  XNOR2_X1  g569(.A(new_n747), .B(new_n673), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n841), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n838), .B(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n997), .B(new_n999), .C1(new_n830), .C2(new_n827), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n991), .B1(new_n993), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(G303), .A2(G8), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1002), .B(KEYINPUT55), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  XOR2_X1   g579(.A(KEYINPUT109), .B(G1971), .Z(new_n1005));
  NAND2_X1  g580(.A1(new_n464), .A2(G125), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n465), .B1(new_n1006), .B2(new_n472), .ZN(new_n1007));
  INV_X1    g582(.A(G40), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1007), .A2(new_n470), .A3(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n990), .B2(KEYINPUT45), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT108), .B1(new_n990), .B2(KEYINPUT45), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n990), .A2(KEYINPUT108), .A3(KEYINPUT45), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1005), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT110), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n1016));
  INV_X1    g591(.A(G1384), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n882), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n882), .A2(new_n1017), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1023), .A2(new_n1019), .A3(KEYINPUT50), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1022), .A2(new_n1009), .A3(new_n1024), .ZN(new_n1025));
  OAI22_X1  g600(.A1(new_n1014), .A2(new_n1015), .B1(new_n1025), .B2(G2090), .ZN(new_n1026));
  AOI211_X1 g601(.A(KEYINPUT110), .B(new_n1005), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1004), .B(G8), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1009), .A2(new_n990), .ZN(new_n1029));
  INV_X1    g604(.A(G1976), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1029), .B(G8), .C1(new_n1030), .C2(G288), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT52), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1032), .B(KEYINPUT112), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1023), .A2(new_n989), .ZN(new_n1034));
  INV_X1    g609(.A(G8), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT52), .B1(G288), .B2(new_n1030), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1036), .B(new_n1037), .C1(new_n1030), .C2(G288), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n607), .A2(G86), .B1(G48), .B2(new_n519), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n584), .A2(new_n585), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(G651), .ZN(new_n1041));
  INV_X1    g616(.A(G1981), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1039), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(G1981), .B1(new_n583), .B2(new_n586), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(new_n1044), .A3(KEYINPUT49), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT49), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1036), .B(new_n1045), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1038), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1033), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1021), .A2(new_n1009), .A3(new_n1018), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(G2090), .ZN(new_n1053));
  OAI21_X1  g628(.A(G8), .B1(new_n1014), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n1003), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1028), .A2(new_n1051), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1025), .A2(new_n783), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1011), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT45), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n989), .B1(new_n1023), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G2078), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .A4(new_n1013), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n990), .A2(KEYINPUT45), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1060), .A2(KEYINPUT53), .A3(new_n1061), .A4(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1057), .A2(new_n1064), .A3(G301), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT54), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1025), .A2(new_n783), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1069));
  OR2_X1    g644(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1070));
  AOI21_X1  g645(.A(G301), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1056), .A2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1022), .A2(new_n767), .A3(new_n1009), .A4(new_n1024), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1060), .A2(new_n1065), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n762), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(G286), .A2(G8), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1074), .A2(KEYINPUT121), .A3(new_n1076), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n1085), .B2(G168), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1077), .A2(G8), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1081), .A2(KEYINPUT51), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(KEYINPUT122), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1035), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1088), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1090), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1083), .B1(new_n1086), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1069), .A2(G301), .A3(new_n1070), .ZN(new_n1097));
  AOI21_X1  g672(.A(G301), .B1(new_n1069), .B2(new_n1066), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT123), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT123), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1101), .B(new_n1096), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1073), .A2(new_n1095), .A3(new_n1100), .A4(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n573), .A2(new_n565), .A3(new_n564), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1104), .A2(KEYINPUT116), .A3(KEYINPUT57), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT57), .B1(new_n1104), .B2(KEYINPUT116), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT56), .B(G2072), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1058), .A2(new_n1060), .A3(new_n1013), .A4(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT115), .ZN(new_n1110));
  INV_X1    g685(.A(G1956), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1009), .B1(new_n990), .B2(new_n1016), .ZN(new_n1112));
  NOR3_X1   g687(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1110), .B(new_n1111), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1110), .B1(new_n1052), .B2(new_n1111), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1107), .B(new_n1109), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1109), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1107), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT115), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n1114), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT117), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(new_n1125), .A3(new_n1107), .A4(new_n1109), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1118), .A2(new_n1121), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1117), .A2(KEYINPUT61), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1119), .A2(new_n1131), .A3(new_n1120), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1131), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1130), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1058), .A2(new_n1060), .A3(new_n1013), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT58), .B(G1341), .ZN(new_n1136));
  OAI22_X1  g711(.A1(new_n1135), .A2(G1996), .B1(new_n1034), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n552), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(KEYINPUT59), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1129), .A2(new_n1134), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT118), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n989), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1142));
  AOI21_X1  g717(.A(G1348), .B1(new_n1142), .B2(new_n1024), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1029), .A2(G2067), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1141), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1144), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT111), .B1(new_n990), .B2(new_n1016), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n990), .A2(new_n1016), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1009), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1024), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI211_X1 g726(.A(KEYINPUT118), .B(new_n1146), .C1(new_n1151), .C2(G1348), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1145), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT60), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT60), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1145), .A2(new_n1155), .A3(new_n1152), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1156), .A2(new_n1157), .A3(new_n609), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1157), .B1(new_n1156), .B2(new_n609), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1154), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1156), .A2(new_n609), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT120), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1154), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1156), .A2(new_n1157), .A3(new_n609), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1140), .A2(new_n1160), .A3(new_n1165), .ZN(new_n1166));
  OAI22_X1  g741(.A1(new_n1132), .A2(new_n1133), .B1(new_n1153), .B2(new_n921), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1167), .A2(new_n1118), .A3(new_n1126), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1103), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1051), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1043), .B(KEYINPUT114), .ZN(new_n1171));
  OR2_X1    g746(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1172));
  NOR2_X1   g747(.A1(G288), .A2(G1976), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1036), .ZN(new_n1175));
  OAI22_X1  g750(.A1(new_n1170), .A2(new_n1028), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT63), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1091), .A2(G168), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1177), .B1(new_n1056), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(G8), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n1003), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1178), .A2(new_n1177), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1181), .A2(new_n1028), .A3(new_n1051), .A4(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1176), .B1(new_n1179), .B2(new_n1183), .ZN(new_n1184));
  AND4_X1   g759(.A1(new_n1055), .A2(new_n1028), .A3(new_n1051), .A4(new_n1098), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1083), .ZN(new_n1186));
  AOI21_X1  g761(.A(KEYINPUT122), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1091), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AND3_X1   g764(.A1(new_n1074), .A2(KEYINPUT121), .A3(new_n1076), .ZN(new_n1190));
  AOI21_X1  g765(.A(KEYINPUT121), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1191));
  OAI21_X1  g766(.A(G168), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1192), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1186), .B1(new_n1189), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT62), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1185), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  OAI211_X1 g771(.A(new_n1083), .B(new_n1195), .C1(new_n1086), .C2(new_n1094), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1197), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1184), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1001), .B1(new_n1169), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n993), .A2(new_n991), .ZN(new_n1201));
  XNOR2_X1  g776(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1202));
  OR2_X1    g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1204));
  INV_X1    g779(.A(new_n991), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1205), .B1(new_n997), .B2(new_n999), .ZN(new_n1206));
  XOR2_X1   g781(.A(new_n1206), .B(KEYINPUT125), .Z(new_n1207));
  NAND3_X1  g782(.A1(new_n1203), .A2(new_n1204), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1205), .B1(new_n994), .B2(new_n748), .ZN(new_n1209));
  AND3_X1   g784(.A1(new_n991), .A2(KEYINPUT46), .A3(new_n673), .ZN(new_n1210));
  AOI21_X1  g785(.A(KEYINPUT46), .B1(new_n991), .B2(new_n673), .ZN(new_n1211));
  NOR3_X1   g786(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  XOR2_X1   g787(.A(new_n1212), .B(KEYINPUT47), .Z(new_n1213));
  NAND2_X1  g788(.A1(new_n839), .A2(new_n998), .ZN(new_n1214));
  OAI22_X1  g789(.A1(new_n996), .A2(new_n1214), .B1(G2067), .B2(new_n728), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1215), .A2(new_n991), .ZN(new_n1216));
  XNOR2_X1  g791(.A(new_n1216), .B(KEYINPUT124), .ZN(new_n1217));
  AND3_X1   g792(.A1(new_n1208), .A2(new_n1213), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1200), .A2(new_n1218), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g794(.A1(new_n652), .A2(new_n654), .ZN(new_n1221));
  NOR2_X1   g795(.A1(G227), .A2(new_n462), .ZN(new_n1222));
  NAND4_X1  g796(.A1(new_n705), .A2(new_n708), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  NOR2_X1   g797(.A1(new_n914), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n1224), .ZN(G225));
  NAND2_X1  g799(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1226));
  INV_X1    g800(.A(KEYINPUT127), .ZN(new_n1227));
  NAND3_X1  g801(.A1(new_n984), .A2(new_n1224), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g802(.A1(new_n1226), .A2(new_n1228), .ZN(G308));
endmodule


