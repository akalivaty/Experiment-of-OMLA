//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1332, new_n1333;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n203), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT66), .Z(new_n223));
  NAND2_X1  g0023(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT65), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n221), .A2(new_n223), .A3(new_n224), .A4(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(new_n209), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n212), .B(new_n217), .C1(new_n228), .C2(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT67), .B(G50), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(KEYINPUT3), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G1698), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n251), .A2(G232), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(G238), .A3(G1698), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G107), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n253), .A2(new_n254), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G274), .ZN(new_n263));
  INV_X1    g0063(.A(new_n215), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT68), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n206), .B(KEYINPUT68), .C1(G41), .C2(G45), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n266), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT69), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n264), .A2(new_n265), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n206), .B(KEYINPUT69), .C1(G41), .C2(G45), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n273), .A2(new_n274), .A3(G244), .A4(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(G200), .B1(new_n262), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n206), .A2(G20), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT72), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n206), .A2(KEYINPUT72), .A3(G13), .A4(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n215), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(KEYINPUT73), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT73), .ZN(new_n289));
  AOI211_X1 g0089(.A(new_n289), .B(new_n286), .C1(new_n282), .C2(new_n283), .ZN(new_n290));
  OAI211_X1 g0090(.A(G77), .B(new_n279), .C1(new_n288), .C2(new_n290), .ZN(new_n291));
  XOR2_X1   g0091(.A(KEYINPUT15), .B(G87), .Z(new_n292));
  NAND2_X1  g0092(.A1(new_n207), .A2(G33), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n292), .A2(new_n294), .B1(G20), .B2(G77), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n207), .A2(new_n248), .A3(KEYINPUT71), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT71), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(G20), .B2(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT8), .B(G58), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n295), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G77), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n282), .A2(new_n283), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n302), .A2(new_n286), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n277), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n261), .A2(new_n306), .A3(G190), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n278), .A2(new_n291), .A3(new_n305), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n291), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(new_n262), .B2(new_n277), .ZN(new_n311));
  INV_X1    g0111(.A(G179), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n261), .A2(new_n306), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n309), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT74), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n316), .A2(KEYINPUT10), .ZN(new_n317));
  INV_X1    g0117(.A(G150), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n300), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(new_n293), .B2(new_n301), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n286), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n280), .A2(new_n215), .A3(new_n285), .ZN(new_n323));
  INV_X1    g0123(.A(G50), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n324), .B1(new_n206), .B2(G20), .ZN(new_n325));
  INV_X1    g0125(.A(new_n280), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n323), .A2(new_n325), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT9), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n322), .A2(KEYINPUT9), .A3(new_n327), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n316), .A2(KEYINPUT10), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n273), .A2(new_n274), .A3(G226), .A4(new_n275), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n271), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n257), .A2(new_n303), .ZN(new_n337));
  NOR2_X1   g0137(.A1(G222), .A2(G1698), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT70), .B(G223), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(G1698), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n260), .B(new_n337), .C1(new_n340), .C2(new_n257), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G200), .ZN(new_n343));
  INV_X1    g0143(.A(G190), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n343), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n317), .B1(new_n333), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G200), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(new_n336), .B2(new_n341), .ZN(new_n348));
  INV_X1    g0148(.A(new_n342), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n348), .B1(new_n349), .B2(G190), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n328), .A2(new_n329), .B1(new_n316), .B2(KEYINPUT10), .ZN(new_n351));
  INV_X1    g0151(.A(new_n317), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n350), .A2(new_n331), .A3(new_n351), .A4(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n349), .A2(new_n312), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n342), .A2(new_n310), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(new_n355), .A3(new_n328), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n315), .A2(new_n346), .A3(new_n353), .A4(new_n356), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n273), .A2(new_n274), .A3(G232), .A4(new_n275), .ZN(new_n358));
  NOR2_X1   g0158(.A1(G223), .A2(G1698), .ZN(new_n359));
  INV_X1    g0159(.A(G226), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n359), .B1(new_n360), .B2(G1698), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n361), .A2(new_n251), .B1(G33), .B2(G87), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n271), .B(new_n358), .C1(new_n362), .C2(new_n274), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n347), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT78), .B1(new_n362), .B2(new_n274), .ZN(new_n365));
  OR2_X1    g0165(.A1(G223), .A2(G1698), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n360), .A2(G1698), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n366), .B(new_n367), .C1(new_n255), .C2(new_n256), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G33), .A2(G87), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT78), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n371), .A3(new_n260), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n365), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n271), .A2(new_n358), .A3(new_n344), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n364), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n249), .A2(new_n207), .A3(new_n250), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT7), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT7), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n249), .A2(new_n378), .A3(new_n207), .A4(new_n250), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(G68), .A3(new_n379), .ZN(new_n380));
  XNOR2_X1  g0180(.A(G58), .B(G68), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n299), .A2(G159), .B1(new_n381), .B2(G20), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT16), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n380), .A2(KEYINPUT16), .A3(new_n382), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n286), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n301), .B1(new_n206), .B2(G20), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n388), .A2(new_n323), .B1(new_n326), .B2(new_n301), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n375), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT17), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n387), .A2(new_n389), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n271), .A2(new_n358), .A3(new_n312), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n394), .A2(new_n365), .A3(new_n372), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n363), .A2(new_n310), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT18), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n393), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n389), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n287), .B1(new_n383), .B2(new_n384), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n401), .B1(new_n402), .B2(new_n386), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT18), .B1(new_n403), .B2(new_n397), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(KEYINPUT17), .A3(new_n375), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n392), .A2(new_n400), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n357), .A2(new_n406), .ZN(new_n407));
  OAI211_X1 g0207(.A(G226), .B(new_n252), .C1(new_n255), .C2(new_n256), .ZN(new_n408));
  OAI211_X1 g0208(.A(G232), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G97), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT75), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n408), .A2(new_n409), .A3(KEYINPUT75), .A4(new_n410), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n414), .A3(new_n260), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n273), .A2(new_n274), .A3(G238), .A4(new_n275), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n271), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT13), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT13), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n415), .A2(new_n420), .A3(new_n417), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(KEYINPUT76), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT76), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n415), .A2(new_n423), .A3(new_n420), .A4(new_n417), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n422), .A2(G200), .A3(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n300), .A2(new_n324), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n293), .A2(new_n303), .B1(new_n207), .B2(G68), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n286), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n428), .B(KEYINPUT11), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n289), .B1(new_n304), .B2(new_n286), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n284), .A2(KEYINPUT73), .A3(new_n287), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(G68), .A3(new_n279), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT12), .B1(new_n284), .B2(G68), .ZN(new_n434));
  INV_X1    g0234(.A(G13), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(G1), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT12), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(G20), .A4(new_n202), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n429), .A2(new_n433), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n419), .A2(G190), .A3(new_n421), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n425), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n419), .A2(G179), .A3(new_n421), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n310), .B1(KEYINPUT77), .B2(KEYINPUT14), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n422), .A2(new_n424), .A3(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(KEYINPUT77), .A2(KEYINPUT14), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n448), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n422), .A2(new_n424), .A3(new_n446), .A4(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n445), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n407), .B(new_n443), .C1(new_n452), .C2(new_n441), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT84), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G283), .ZN(new_n456));
  OAI211_X1 g0256(.A(G250), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n457));
  OAI211_X1 g0257(.A(G244), .B(new_n252), .C1(new_n255), .C2(new_n256), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT4), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n456), .B(new_n457), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(G1698), .B1(new_n249), .B2(new_n250), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT4), .B1(new_n461), .B2(G244), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n260), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT80), .ZN(new_n464));
  INV_X1    g0264(.A(G41), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT5), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT5), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(KEYINPUT80), .B2(G41), .ZN(new_n468));
  INV_X1    g0268(.A(G45), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G1), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n266), .A2(new_n466), .A3(new_n468), .A4(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n466), .A2(new_n468), .A3(new_n470), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(G257), .A3(new_n274), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(G169), .B1(new_n463), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n471), .A2(new_n473), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n461), .A2(KEYINPUT4), .A3(G244), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n458), .A2(new_n459), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n478), .A2(new_n479), .A3(new_n456), .A4(new_n457), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n477), .B1(new_n480), .B2(new_n260), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n312), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT6), .ZN(new_n483));
  AND2_X1   g0283(.A1(G97), .A2(G107), .ZN(new_n484));
  NOR2_X1   g0284(.A1(G97), .A2(G107), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G107), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(KEYINPUT6), .A3(G97), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n489), .A2(G20), .B1(G77), .B2(new_n299), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n377), .A2(KEYINPUT79), .A3(G107), .A4(new_n379), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n377), .A2(G107), .A3(new_n379), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT79), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n287), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G97), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n326), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n206), .A2(G33), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n280), .A2(new_n499), .A3(new_n215), .A4(new_n285), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n498), .B1(new_n500), .B2(new_n497), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n476), .B(new_n482), .C1(new_n496), .C2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n495), .A2(new_n491), .A3(new_n490), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n501), .B1(new_n503), .B2(new_n286), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n463), .A2(new_n474), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G200), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n481), .A2(G190), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n206), .A2(G45), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G250), .ZN(new_n511));
  OAI22_X1  g0311(.A1(new_n260), .A2(new_n511), .B1(new_n263), .B2(new_n510), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT81), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(G116), .ZN(new_n514));
  INV_X1    g0314(.A(G116), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(KEYINPUT81), .ZN(new_n516));
  OAI21_X1  g0316(.A(G33), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(G244), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n518));
  OAI211_X1 g0318(.A(G238), .B(new_n252), .C1(new_n255), .C2(new_n256), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n512), .B1(new_n520), .B2(new_n260), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G190), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT83), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n520), .A2(new_n260), .ZN(new_n524));
  INV_X1    g0324(.A(new_n512), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G200), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT19), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n207), .B1(new_n410), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(G87), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n485), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n207), .B(G68), .C1(new_n255), .C2(new_n256), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n528), .B1(new_n293), .B2(new_n497), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n286), .ZN(new_n536));
  XNOR2_X1  g0336(.A(KEYINPUT15), .B(G87), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n304), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n323), .A2(G87), .A3(new_n499), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT83), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n521), .A2(new_n542), .A3(G190), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n523), .A2(new_n527), .A3(new_n541), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n526), .A2(new_n310), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n323), .A2(KEYINPUT82), .A3(new_n292), .A4(new_n499), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT82), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n500), .B2(new_n537), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n535), .A2(new_n286), .B1(new_n304), .B2(new_n537), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n521), .A2(new_n312), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n545), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n544), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n455), .B1(new_n509), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n554), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n556), .A2(KEYINPUT84), .A3(new_n502), .A4(new_n508), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT85), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(KEYINPUT21), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n515), .A2(KEYINPUT81), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n513), .A2(G116), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n563), .A2(new_n282), .A3(new_n283), .ZN(new_n564));
  AOI21_X1  g0364(.A(G20), .B1(G33), .B2(G283), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n248), .A2(G97), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n565), .A2(new_n566), .B1(new_n285), .B2(new_n215), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n560), .A2(new_n561), .A3(G20), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n567), .A2(KEYINPUT20), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT20), .B1(new_n567), .B2(new_n568), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n564), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n515), .B1(new_n206), .B2(G33), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n571), .B1(new_n432), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(G264), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n574));
  OAI211_X1 g0374(.A(G257), .B(new_n252), .C1(new_n255), .C2(new_n256), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n249), .A2(G303), .A3(new_n250), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n260), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n472), .A2(G270), .A3(new_n274), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(new_n471), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G169), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n559), .B1(new_n573), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n572), .B1(new_n288), .B2(new_n290), .ZN(new_n583));
  OR2_X1    g0383(.A1(new_n569), .A2(new_n570), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(new_n584), .A3(new_n564), .ZN(new_n585));
  INV_X1    g0385(.A(new_n559), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n471), .A2(new_n579), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n310), .B1(new_n587), .B2(new_n578), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n580), .A2(new_n312), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n582), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n207), .B(G87), .C1(new_n255), .C2(new_n256), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT22), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT22), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n251), .A2(new_n595), .A3(new_n207), .A4(G87), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT24), .ZN(new_n598));
  OAI21_X1  g0398(.A(KEYINPUT86), .B1(new_n207), .B2(G107), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT23), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT23), .ZN(new_n601));
  OAI211_X1 g0401(.A(KEYINPUT86), .B(new_n601), .C1(new_n207), .C2(G107), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n600), .A2(new_n602), .B1(new_n562), .B2(new_n294), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n597), .A2(new_n598), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n598), .B1(new_n597), .B2(new_n603), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n286), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n280), .A2(G107), .ZN(new_n607));
  XNOR2_X1  g0407(.A(KEYINPUT87), .B(KEYINPUT25), .ZN(new_n608));
  XNOR2_X1  g0408(.A(new_n607), .B(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n500), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n609), .B1(G107), .B2(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(G257), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n612));
  OAI211_X1 g0412(.A(G250), .B(new_n252), .C1(new_n255), .C2(new_n256), .ZN(new_n613));
  INV_X1    g0413(.A(G294), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n612), .B(new_n613), .C1(new_n248), .C2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n260), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n472), .A2(G264), .A3(new_n274), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n616), .A2(G190), .A3(new_n471), .A4(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n471), .A3(new_n617), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(G200), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n606), .A2(new_n611), .A3(new_n618), .A4(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n578), .A2(new_n471), .A3(new_n579), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(G190), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n580), .A2(G200), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(new_n573), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n619), .A2(new_n310), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n616), .A2(new_n312), .A3(new_n471), .A4(new_n617), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n606), .B2(new_n611), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n592), .A2(new_n626), .A3(new_n630), .ZN(new_n631));
  AND4_X1   g0431(.A1(new_n454), .A2(new_n555), .A3(new_n557), .A4(new_n631), .ZN(G372));
  NAND2_X1  g0432(.A1(new_n400), .A2(new_n404), .ZN(new_n633));
  INV_X1    g0433(.A(new_n314), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n443), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n452), .B2(new_n441), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n392), .A2(new_n405), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n633), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n346), .A2(new_n353), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n356), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n592), .A2(new_n630), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n540), .B1(G200), .B2(new_n526), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n549), .A2(new_n550), .B1(new_n521), .B2(new_n312), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n645), .A2(new_n522), .B1(new_n646), .B2(new_n545), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n502), .A2(new_n647), .A3(new_n508), .A4(new_n621), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT26), .B1(new_n554), .B2(new_n502), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n463), .A2(new_n312), .A3(new_n474), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n504), .A2(new_n651), .A3(new_n475), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT26), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(new_n653), .A3(new_n647), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n650), .A2(new_n553), .A3(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n643), .B1(new_n453), .B2(new_n656), .ZN(G369));
  NAND2_X1  g0457(.A1(new_n606), .A2(new_n611), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n436), .A2(new_n207), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G213), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G343), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n630), .B1(new_n665), .B2(new_n621), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n627), .A2(new_n628), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n658), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(new_n664), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n664), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(new_n592), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n669), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n674), .A2(KEYINPUT88), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(KEYINPUT88), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n573), .A2(new_n671), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n592), .B(new_n678), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n679), .A2(new_n625), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n680), .A2(G330), .A3(new_n670), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n677), .A2(new_n681), .ZN(G399));
  NAND2_X1  g0482(.A1(new_n210), .A2(new_n465), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n531), .A2(G116), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G1), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n213), .B2(new_n683), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT28), .ZN(new_n687));
  INV_X1    g0487(.A(G330), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT30), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n521), .A2(KEYINPUT89), .A3(new_n616), .A4(new_n617), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n690), .A2(new_n481), .A3(new_n622), .A4(G179), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n616), .A2(new_n617), .ZN(new_n692));
  AOI21_X1  g0492(.A(KEYINPUT89), .B1(new_n692), .B2(new_n521), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n689), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n505), .A2(new_n312), .A3(new_n580), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT89), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n616), .A2(new_n617), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n696), .B1(new_n697), .B2(new_n526), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n695), .A2(KEYINPUT30), .A3(new_n698), .A4(new_n690), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n521), .A2(G179), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n700), .A2(new_n505), .A3(new_n619), .A4(new_n580), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n694), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n702), .A2(KEYINPUT31), .A3(new_n664), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT31), .B1(new_n702), .B2(new_n664), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n631), .A2(new_n557), .A3(new_n555), .A4(new_n671), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n688), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT29), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n656), .B2(new_n664), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT91), .B1(new_n592), .B2(new_n630), .ZN(new_n710));
  AND4_X1   g0510(.A1(new_n502), .A2(new_n647), .A3(new_n508), .A4(new_n621), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n585), .A2(new_n588), .ZN(new_n712));
  AOI22_X1  g0512(.A1(new_n712), .A2(new_n559), .B1(new_n585), .B2(new_n590), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT91), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n713), .A2(new_n668), .A3(new_n714), .A4(new_n589), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n710), .A2(new_n711), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT90), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n651), .A2(new_n475), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n493), .A2(new_n494), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n490), .A2(new_n491), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n286), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n501), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n527), .A2(new_n541), .A3(new_n522), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n718), .A2(new_n723), .A3(new_n553), .A4(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n717), .B1(new_n725), .B2(new_n653), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n653), .B1(new_n554), .B2(new_n502), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n652), .A2(new_n647), .A3(KEYINPUT90), .A4(KEYINPUT26), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n716), .A2(new_n729), .A3(new_n553), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(KEYINPUT29), .A3(new_n671), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n707), .B1(new_n709), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n687), .B1(new_n732), .B2(G1), .ZN(G364));
  INV_X1    g0533(.A(new_n683), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n435), .A2(new_n469), .A3(G20), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n735), .A2(KEYINPUT92), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(KEYINPUT92), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n736), .A2(G1), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n210), .A2(new_n251), .ZN(new_n740));
  INV_X1    g0540(.A(G355), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n740), .A2(new_n741), .B1(G116), .B2(new_n210), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n242), .A2(G45), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n210), .A2(new_n257), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(new_n469), .B2(new_n214), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n742), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n264), .B1(new_n207), .B2(G169), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n747), .A2(KEYINPUT93), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(KEYINPUT93), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n739), .B1(new_n746), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n207), .A2(new_n344), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n347), .A2(G179), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n530), .ZN(new_n760));
  INV_X1    g0560(.A(new_n757), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n761), .A2(new_n312), .A3(G200), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n312), .A2(new_n347), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n757), .A2(new_n764), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n763), .A2(new_n201), .B1(new_n765), .B2(new_n324), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n207), .A2(G190), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n760), .B(new_n766), .C1(G68), .C2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G179), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G190), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n497), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n767), .A2(new_n758), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n487), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n775), .A2(new_n257), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n767), .A2(new_n771), .ZN(new_n779));
  INV_X1    g0579(.A(G159), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT32), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n767), .A2(G179), .A3(new_n347), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n784), .A2(KEYINPUT94), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(KEYINPUT94), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G77), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n770), .A2(new_n778), .A3(new_n782), .A4(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G317), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n791), .A2(KEYINPUT33), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(KEYINPUT33), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n768), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G322), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n763), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n779), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n794), .B(new_n796), .C1(G329), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n773), .A2(G294), .ZN(new_n799));
  INV_X1    g0599(.A(G311), .ZN(new_n800));
  INV_X1    g0600(.A(G303), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n800), .A2(new_n783), .B1(new_n759), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n776), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n251), .B(new_n802), .C1(G283), .C2(new_n803), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n765), .B(KEYINPUT95), .Z(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G326), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n798), .A2(new_n799), .A3(new_n804), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n790), .A2(new_n808), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n809), .A2(KEYINPUT96), .ZN(new_n810));
  INV_X1    g0610(.A(new_n750), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(new_n809), .B2(KEYINPUT96), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n756), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n753), .B(KEYINPUT97), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n680), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n680), .A2(G330), .ZN(new_n816));
  INV_X1    g0616(.A(new_n739), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n680), .A2(G330), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n815), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT98), .Z(G396));
  NOR2_X1   g0621(.A1(new_n750), .A2(new_n751), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n739), .B1(new_n823), .B2(G77), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n763), .A2(new_n614), .B1(new_n765), .B2(new_n801), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n251), .B(new_n825), .C1(G283), .C2(new_n769), .ZN(new_n826));
  INV_X1    g0626(.A(new_n775), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n788), .A2(new_n562), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n759), .A2(new_n487), .B1(new_n779), .B2(new_n800), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(G87), .B2(new_n803), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n826), .A2(new_n827), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n759), .A2(new_n324), .B1(new_n776), .B2(new_n202), .ZN(new_n832));
  INV_X1    g0632(.A(G132), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n251), .B1(new_n779), .B2(new_n833), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT99), .Z(new_n835));
  AOI211_X1 g0635(.A(new_n832), .B(new_n835), .C1(G58), .C2(new_n773), .ZN(new_n836));
  INV_X1    g0636(.A(new_n765), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n762), .A2(G143), .B1(new_n837), .B2(G137), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n838), .B1(new_n318), .B2(new_n768), .C1(new_n787), .C2(new_n780), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n836), .B1(new_n840), .B2(KEYINPUT34), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT34), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n831), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n824), .B1(new_n844), .B2(new_n750), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n671), .B1(new_n291), .B2(new_n305), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n308), .B1(new_n846), .B2(KEYINPUT100), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n846), .A2(KEYINPUT100), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n314), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n634), .A2(new_n671), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n845), .B1(new_n852), .B2(new_n752), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n851), .B1(new_n656), .B2(new_n664), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n852), .B(new_n671), .C1(new_n649), .C2(new_n655), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n707), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n855), .A2(new_n856), .ZN(new_n858));
  INV_X1    g0658(.A(new_n707), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n739), .B(new_n857), .C1(KEYINPUT101), .C2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(KEYINPUT101), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n854), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(G384));
  AOI21_X1  g0665(.A(new_n206), .B1(G13), .B2(new_n207), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n393), .A2(new_n398), .ZN(new_n867));
  INV_X1    g0667(.A(new_n662), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n393), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n867), .A2(new_n869), .A3(new_n390), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT37), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n867), .A2(new_n869), .A3(new_n872), .A4(new_n390), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n871), .A2(KEYINPUT103), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n869), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n406), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT103), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n870), .A2(new_n877), .A3(KEYINPUT37), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n874), .A2(KEYINPUT38), .A3(new_n876), .A4(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT104), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n375), .A2(new_n387), .A3(new_n389), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n397), .B1(new_n387), .B2(new_n389), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n872), .B1(new_n884), .B2(new_n869), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n885), .A2(new_n877), .B1(new_n406), .B2(new_n875), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n886), .B2(new_n874), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n881), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n874), .A2(new_n876), .A3(new_n878), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n889), .A2(KEYINPUT104), .A3(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT39), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT106), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n871), .A2(new_n873), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n876), .ZN(new_n896));
  XNOR2_X1  g0696(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n879), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT39), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n893), .A2(new_n894), .A3(new_n901), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n871), .A2(KEYINPUT103), .A3(new_n873), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n876), .A2(new_n878), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n890), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(new_n880), .A3(new_n879), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n900), .B1(new_n906), .B2(new_n891), .ZN(new_n907));
  INV_X1    g0707(.A(new_n901), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT106), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n449), .A2(new_n451), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n444), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(new_n440), .A3(new_n671), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n902), .A2(new_n909), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n856), .A2(new_n850), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n440), .A2(new_n664), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n443), .B(new_n916), .C1(new_n452), .C2(new_n441), .ZN(new_n917));
  INV_X1    g0717(.A(new_n916), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n911), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n921), .A2(new_n888), .A3(new_n892), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(new_n633), .B2(new_n662), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n914), .A2(new_n923), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n454), .A2(new_n731), .A3(new_n709), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n925), .A2(new_n642), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n924), .B(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n851), .B1(new_n917), .B2(new_n919), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n705), .A2(new_n706), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n928), .A2(new_n929), .A3(new_n899), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT40), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n928), .A2(new_n929), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT40), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n906), .A2(new_n933), .A3(new_n891), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n931), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n453), .B1(new_n706), .B2(new_n705), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n935), .A2(new_n936), .ZN(new_n939));
  NOR3_X1   g0739(.A1(new_n938), .A2(new_n939), .A3(new_n688), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n866), .B1(new_n927), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n927), .B2(new_n941), .ZN(new_n943));
  OAI211_X1 g0743(.A(G116), .B(new_n216), .C1(new_n489), .C2(KEYINPUT35), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT102), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n945), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n489), .A2(KEYINPUT35), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT36), .ZN(new_n950));
  OAI21_X1  g0750(.A(G77), .B1(new_n201), .B2(new_n202), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n213), .A2(new_n951), .B1(G50), .B2(new_n202), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n952), .A2(G1), .A3(new_n435), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n943), .A2(new_n950), .A3(new_n953), .ZN(G367));
  AOI21_X1  g0754(.A(new_n509), .B1(new_n723), .B2(new_n664), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT109), .Z(new_n956));
  NAND2_X1  g0756(.A1(new_n652), .A2(new_n664), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OR3_X1    g0758(.A1(new_n958), .A2(KEYINPUT42), .A3(new_n672), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n502), .B1(new_n956), .B2(new_n668), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n671), .ZN(new_n961));
  OAI21_X1  g0761(.A(KEYINPUT42), .B1(new_n958), .B2(new_n672), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n664), .A2(new_n540), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT107), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n647), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n967), .A2(KEYINPUT108), .B1(new_n553), .B2(new_n966), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(KEYINPUT108), .B2(new_n967), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT43), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n963), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n969), .A2(new_n970), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n963), .A2(new_n970), .A3(new_n969), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n958), .ZN(new_n977));
  INV_X1    g0777(.A(new_n681), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT110), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n976), .B(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(KEYINPUT111), .B(KEYINPUT41), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n683), .B(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n677), .A2(new_n977), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT45), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n675), .A2(new_n958), .A3(new_n676), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT44), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n978), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT45), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n985), .B(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT44), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n987), .B(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n991), .A2(new_n681), .A3(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n670), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n592), .A2(new_n671), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n672), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(new_n816), .Z(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n732), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n989), .A2(new_n994), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n984), .B1(new_n1002), .B2(new_n732), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n981), .B1(new_n1003), .B2(new_n738), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n814), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n969), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n754), .B1(new_n210), .B2(new_n537), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n237), .A2(new_n744), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n739), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(G294), .A2(new_n769), .B1(new_n797), .B2(G317), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n759), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1011), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1010), .B(new_n1012), .C1(new_n801), .C2(new_n763), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n805), .A2(new_n800), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(G283), .C2(new_n788), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n257), .B1(new_n776), .B2(new_n497), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(KEYINPUT112), .B(KEYINPUT46), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n1011), .B2(new_n562), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1016), .B(new_n1018), .C1(G107), .C2(new_n773), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n763), .A2(new_n318), .B1(new_n768), .B2(new_n780), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n251), .B1(new_n759), .B2(new_n201), .C1(new_n774), .C2(new_n202), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n803), .A2(G77), .ZN(new_n1022));
  INV_X1    g0822(.A(G137), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1022), .B1(new_n1023), .B2(new_n779), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1020), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n788), .A2(G50), .B1(new_n806), .B2(G143), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n1015), .A2(new_n1019), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1027), .A2(KEYINPUT47), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n811), .B1(new_n1027), .B2(KEYINPUT47), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1009), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1006), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1004), .A2(new_n1031), .ZN(G387));
  OAI22_X1  g0832(.A1(new_n740), .A2(new_n684), .B1(G107), .B2(new_n210), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n234), .A2(new_n469), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n684), .ZN(new_n1035));
  AOI211_X1 g0835(.A(G45), .B(new_n1035), .C1(G68), .C2(G77), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n301), .A2(G50), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT50), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n744), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1033), .B1(new_n1034), .B2(new_n1039), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n784), .A2(G68), .B1(new_n797), .B2(G150), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n301), .B2(new_n768), .C1(new_n324), .C2(new_n763), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n774), .A2(new_n537), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n251), .B1(new_n776), .B2(new_n497), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n765), .A2(new_n780), .B1(new_n759), .B2(new_n303), .ZN(new_n1045));
  NOR4_X1   g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(G283), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n774), .A2(new_n1047), .B1(new_n759), .B2(new_n614), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT113), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n762), .A2(G317), .B1(G311), .B2(new_n769), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n805), .B2(new_n795), .C1(new_n787), .C2(new_n801), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT48), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n1052), .B2(new_n1051), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1054), .A2(KEYINPUT49), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n251), .B1(new_n797), .B2(G326), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n563), .B2(new_n776), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n1054), .B2(KEYINPUT49), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1046), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n739), .B1(new_n755), .B2(new_n1040), .C1(new_n1059), .C2(new_n811), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n995), .B2(new_n1005), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n999), .B2(new_n738), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1000), .A2(new_n734), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n999), .A2(new_n732), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(G393));
  NOR3_X1   g0865(.A1(new_n986), .A2(new_n978), .A3(new_n988), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n681), .B1(new_n991), .B2(new_n993), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n958), .A2(new_n753), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n754), .B1(new_n497), .B2(new_n210), .ZN(new_n1070));
  AND3_X1   g0870(.A1(new_n245), .A2(new_n210), .A3(new_n257), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n739), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n774), .A2(new_n303), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n257), .B(new_n1073), .C1(G87), .C2(new_n803), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n324), .A2(new_n768), .B1(new_n759), .B2(new_n202), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(G143), .B2(new_n797), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1074), .B(new_n1076), .C1(new_n301), .C2(new_n787), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n762), .A2(G159), .B1(new_n837), .B2(G150), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT51), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n762), .A2(G311), .B1(new_n837), .B2(G317), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT52), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n251), .B(new_n777), .C1(new_n562), .C2(new_n773), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n784), .A2(G294), .B1(new_n769), .B2(G303), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(G283), .A2(new_n1011), .B1(new_n797), .B2(G322), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n1077), .A2(new_n1079), .B1(new_n1081), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1072), .B1(new_n1086), .B2(new_n750), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1068), .A2(new_n738), .B1(new_n1069), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1000), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1089), .A2(new_n734), .A3(new_n1002), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1088), .A2(new_n1090), .ZN(G390));
  NAND2_X1  g0891(.A1(new_n921), .A2(new_n912), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n894), .B1(new_n893), .B2(new_n901), .ZN(new_n1093));
  NOR3_X1   g0893(.A1(new_n907), .A2(new_n908), .A3(KEYINPUT106), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1092), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n920), .A2(new_n707), .A3(new_n852), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n730), .A2(new_n671), .A3(new_n849), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n1097), .A2(new_n850), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n917), .A2(new_n919), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n899), .A2(new_n912), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1095), .A2(new_n1096), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1096), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1092), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n902), .B2(new_n909), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1105), .B1(new_n1107), .B2(new_n1102), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1104), .A2(new_n1108), .A3(new_n738), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n751), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n837), .A2(G283), .B1(new_n797), .B2(G294), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n487), .B2(new_n768), .C1(new_n787), .C2(new_n497), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n760), .A2(new_n251), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1113), .B1(new_n202), .B2(new_n776), .C1(new_n763), .C2(new_n515), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n1112), .A2(new_n1073), .A3(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT117), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n759), .A2(new_n318), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT53), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT54), .B(G143), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT115), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1118), .B1(new_n787), .B2(new_n1120), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n762), .A2(G132), .B1(new_n837), .B2(G128), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G137), .A2(new_n769), .B1(new_n797), .B2(G125), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n251), .B1(new_n776), .B2(new_n324), .C1(new_n774), .C2(new_n780), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n1121), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT116), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n811), .B1(new_n1116), .B2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n817), .B(new_n1128), .C1(new_n301), .C2(new_n822), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1110), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1109), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n911), .A2(new_n440), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n637), .B1(new_n1133), .B2(new_n635), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n640), .B1(new_n1134), .B2(new_n633), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n454), .A2(new_n731), .A3(new_n709), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n454), .A2(new_n707), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1135), .A2(new_n356), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT114), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AND4_X1   g0940(.A1(new_n555), .A2(new_n631), .A3(new_n557), .A4(new_n671), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n702), .A2(new_n664), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT31), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n702), .A2(KEYINPUT31), .A3(new_n664), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g0946(.A(G330), .B(new_n852), .C1(new_n1141), .C2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1099), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1148), .A2(new_n1098), .A3(new_n1096), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1099), .A2(new_n1147), .B1(new_n928), .B2(new_n707), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n856), .A2(new_n850), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n643), .A2(KEYINPUT114), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1140), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n683), .B1(new_n1132), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1154), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1104), .A2(new_n1108), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1131), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(G378));
  NAND2_X1  g0959(.A1(new_n640), .A2(new_n356), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1160), .A2(new_n328), .A3(new_n868), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n328), .A2(new_n868), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n640), .A2(new_n356), .A3(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n1161), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1164), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n751), .ZN(new_n1168));
  AOI21_X1  g0968(.A(G50), .B1(new_n250), .B2(new_n465), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n776), .A2(new_n201), .B1(new_n779), .B2(new_n1047), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n465), .B(new_n257), .C1(new_n759), .C2(new_n303), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(G68), .C2(new_n773), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n837), .A2(G116), .B1(new_n784), .B2(new_n292), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n762), .A2(G107), .B1(G97), .B2(new_n769), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT58), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1169), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1120), .A2(new_n759), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n762), .A2(G128), .B1(new_n837), .B2(G125), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n784), .A2(G137), .B1(new_n769), .B2(G132), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1178), .B(new_n1181), .C1(G150), .C2(new_n773), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT59), .Z(new_n1183));
  AOI211_X1 g0983(.A(G33), .B(G41), .C1(new_n803), .C2(G159), .ZN(new_n1184));
  INV_X1    g0984(.A(G124), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1184), .B1(new_n1185), .B2(new_n779), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1177), .B1(new_n1176), .B2(new_n1175), .C1(new_n1183), .C2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n750), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n822), .A2(new_n324), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1168), .A2(new_n739), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n906), .A2(new_n933), .A3(new_n891), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n932), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1192), .A2(new_n1193), .B1(KEYINPUT40), .B2(new_n930), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1167), .B1(new_n1194), .B2(new_n688), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1167), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n935), .A2(G330), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n914), .A2(new_n923), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1195), .A2(new_n914), .A3(new_n923), .A4(new_n1197), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1191), .B1(new_n1202), .B2(new_n738), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1140), .A2(new_n1153), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT118), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1204), .B(new_n1205), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1157), .A2(new_n1206), .B1(new_n1201), .B2(new_n1200), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n734), .B1(new_n1207), .B2(KEYINPUT57), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT119), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n924), .A2(new_n1209), .A3(new_n1195), .A4(new_n1197), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1201), .A2(KEYINPUT119), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1210), .A2(new_n1211), .A3(new_n1200), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1157), .A2(new_n1206), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1212), .A2(KEYINPUT57), .A3(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1203), .B1(new_n1208), .B2(new_n1214), .ZN(G375));
  AOI21_X1  g1015(.A(new_n1152), .B1(new_n1140), .B2(new_n1153), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1156), .A2(new_n1216), .A3(new_n984), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT120), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1152), .A2(new_n738), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n739), .B1(new_n823), .B2(G68), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n251), .B1(new_n776), .B2(new_n201), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT121), .Z(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n768), .B2(new_n1120), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n784), .A2(G150), .B1(new_n1011), .B2(G159), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n837), .A2(G132), .B1(new_n797), .B2(G128), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n762), .A2(G137), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n773), .A2(G50), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G97), .A2(new_n1011), .B1(new_n797), .B2(G303), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1229), .B1(new_n563), .B2(new_n768), .C1(new_n787), .C2(new_n487), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n762), .A2(G283), .B1(new_n837), .B2(G294), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1043), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1231), .A2(new_n1232), .A3(new_n257), .A4(new_n1022), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1223), .A2(new_n1228), .B1(new_n1230), .B2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1220), .B1(new_n1234), .B2(new_n750), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n920), .B2(new_n752), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1219), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1218), .A2(new_n1238), .ZN(G381));
  OR3_X1    g1039(.A1(G384), .A2(G393), .A3(G396), .ZN(new_n1240));
  NOR4_X1   g1040(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1240), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(KEYINPUT122), .Z(new_n1242));
  INV_X1    g1042(.A(G375), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1158), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1245), .ZN(G407));
  OAI211_X1 g1046(.A(G407), .B(G213), .C1(G343), .C2(new_n1244), .ZN(G409));
  XOR2_X1   g1047(.A(G393), .B(G396), .Z(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1004), .A2(G390), .A3(new_n1031), .ZN(new_n1250));
  AOI21_X1  g1050(.A(G390), .B1(new_n1004), .B2(new_n1031), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1249), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(G390), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G387), .A2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1004), .A2(G390), .A3(new_n1031), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n1248), .A3(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT61), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1252), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n1258), .A2(KEYINPUT125), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1258), .A2(KEYINPUT125), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G375), .A2(G378), .ZN(new_n1262));
  INV_X1    g1062(.A(G213), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1263), .A2(G343), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1096), .B1(new_n1095), .B2(new_n1103), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1107), .A2(new_n1105), .A3(new_n1102), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1154), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(new_n734), .A3(new_n1157), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1109), .A2(new_n1130), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n1269), .A3(new_n1190), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1213), .A2(new_n983), .A3(new_n1202), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1212), .A2(new_n738), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1264), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT123), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n734), .B(new_n1154), .C1(new_n1216), .C2(KEYINPUT60), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1151), .B1(new_n1148), .B2(new_n1096), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n1098), .B2(new_n1150), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT114), .B1(new_n926), .B2(new_n1137), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1278), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT60), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1275), .B1(new_n1276), .B2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1154), .A2(new_n734), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1216), .A2(KEYINPUT60), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1285), .A2(new_n1286), .A3(KEYINPUT123), .A4(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1284), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(G384), .B1(new_n1289), .B2(new_n1238), .ZN(new_n1290));
  AOI211_X1 g1090(.A(new_n864), .B(new_n1237), .C1(new_n1284), .C2(new_n1288), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1262), .A2(new_n1274), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1289), .A2(new_n1238), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n864), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT124), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1289), .A2(G384), .A3(new_n1238), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1295), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(KEYINPUT124), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1264), .A2(G2897), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1300), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1292), .A2(new_n1296), .A3(new_n1302), .ZN(new_n1303));
  AOI22_X1  g1103(.A1(new_n1301), .A2(new_n1303), .B1(new_n1262), .B2(new_n1274), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT63), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1293), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1261), .B(new_n1306), .C1(new_n1305), .C2(new_n1293), .ZN(new_n1307));
  NOR4_X1   g1107(.A1(new_n1290), .A2(new_n1291), .A3(KEYINPUT124), .A4(new_n1300), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1302), .B1(new_n1292), .B2(new_n1296), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1308), .B1(new_n1309), .B2(new_n1299), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1212), .A2(KEYINPUT57), .A3(new_n1213), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1311), .B(new_n734), .C1(KEYINPUT57), .C2(new_n1207), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1158), .B1(new_n1312), .B2(new_n1203), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1207), .A2(new_n983), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1158), .A2(new_n1314), .A3(new_n1190), .A4(new_n1273), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1263), .B2(G343), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1313), .A2(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1257), .B1(new_n1310), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT62), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1293), .A2(new_n1319), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1262), .A2(new_n1274), .A3(KEYINPUT62), .A4(new_n1292), .ZN(new_n1321));
  AOI22_X1  g1121(.A1(new_n1318), .A2(KEYINPUT126), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT126), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n1323), .B(new_n1257), .C1(new_n1310), .C2(new_n1317), .ZN(new_n1324));
  AOI21_X1  g1124(.A(KEYINPUT127), .B1(new_n1322), .B2(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(KEYINPUT126), .B1(new_n1304), .B2(KEYINPUT61), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1326), .A2(new_n1324), .A3(KEYINPUT127), .A4(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1252), .A2(new_n1256), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1307), .B1(new_n1325), .B2(new_n1330), .ZN(G405));
  NAND2_X1  g1131(.A1(new_n1244), .A2(new_n1262), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(new_n1332), .B(new_n1292), .ZN(new_n1333));
  XOR2_X1   g1133(.A(new_n1333), .B(new_n1329), .Z(G402));
endmodule


