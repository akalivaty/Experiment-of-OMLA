//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 1 0 0 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1221, new_n1222, new_n1223, new_n1224, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1298, new_n1299;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n207));
  INV_X1    g0007(.A(G226), .ZN(new_n208));
  INV_X1    g0008(.A(G116), .ZN(new_n209));
  INV_X1    g0009(.A(G270), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n207), .B1(new_n202), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G58), .ZN(new_n213));
  INV_X1    g0013(.A(G232), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n206), .B1(new_n211), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  AND3_X1   g0019(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n220));
  AOI21_X1  g0020(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n206), .A2(G13), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT0), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n219), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n218), .ZN(G361));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT65), .B(KEYINPUT66), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n214), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT67), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n246), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G274), .ZN(new_n252));
  AND2_X1   g0052(.A1(G1), .A2(G13), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n254), .A2(G1), .A3(G13), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n257), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n259), .B1(new_n208), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G222), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G77), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n263), .A2(G1698), .ZN(new_n267));
  INV_X1    g0067(.A(G223), .ZN(new_n268));
  OAI221_X1 g0068(.A(new_n265), .B1(new_n266), .B2(new_n263), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n254), .B1(new_n220), .B2(new_n221), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n262), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n203), .A2(G20), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G150), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n223), .A2(G33), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n273), .B(new_n275), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n222), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n278), .A2(new_n280), .B1(new_n202), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G1), .A2(G13), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT64), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n286), .A2(new_n281), .A3(new_n287), .A4(new_n279), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n256), .A2(G20), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(G50), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n283), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT9), .ZN(new_n293));
  AOI22_X1  g0093(.A1(G190), .A2(new_n272), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n283), .A2(KEYINPUT9), .A3(new_n291), .ZN(new_n295));
  INV_X1    g0095(.A(new_n272), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G200), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n294), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT10), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n294), .A2(new_n297), .A3(new_n295), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n292), .B1(new_n272), .B2(G169), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT68), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n304), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n305), .B(new_n306), .C1(G179), .C2(new_n296), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n263), .A2(G232), .A3(new_n264), .ZN(new_n308));
  INV_X1    g0108(.A(G107), .ZN(new_n309));
  INV_X1    g0109(.A(G238), .ZN(new_n310));
  OAI221_X1 g0110(.A(new_n308), .B1(new_n309), .B2(new_n263), .C1(new_n267), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n271), .ZN(new_n312));
  INV_X1    g0112(.A(new_n261), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n313), .A2(G244), .B1(new_n258), .B2(new_n255), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G200), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n312), .A2(G190), .A3(new_n314), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n289), .A2(G77), .A3(new_n290), .ZN(new_n318));
  INV_X1    g0118(.A(new_n277), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n319), .A2(new_n274), .B1(G20), .B2(G77), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT15), .B(G87), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n276), .B2(new_n321), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n322), .A2(new_n280), .B1(new_n266), .B2(new_n282), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n316), .A2(new_n317), .A3(new_n318), .A4(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G169), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n315), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n323), .A2(new_n318), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n326), .B(new_n327), .C1(G179), .C2(new_n315), .ZN(new_n328));
  AND4_X1   g0128(.A1(new_n302), .A2(new_n307), .A3(new_n324), .A4(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n263), .A2(G226), .A3(new_n264), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT69), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT69), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n263), .A2(new_n332), .A3(G226), .A4(new_n264), .ZN(new_n333));
  NAND2_X1  g0133(.A1(G33), .A2(G97), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n263), .A2(G232), .A3(G1698), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n331), .A2(new_n333), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n271), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n259), .B1(new_n310), .B2(new_n261), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT13), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT13), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n337), .A2(new_n342), .A3(new_n339), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(G190), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n342), .B1(new_n337), .B2(new_n339), .ZN(new_n345));
  AOI211_X1 g0145(.A(KEYINPUT13), .B(new_n338), .C1(new_n336), .C2(new_n271), .ZN(new_n346));
  OAI21_X1  g0146(.A(G200), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G68), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n274), .A2(G50), .B1(G20), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n266), .B2(new_n276), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n280), .ZN(new_n351));
  XOR2_X1   g0151(.A(new_n351), .B(KEYINPUT11), .Z(new_n352));
  NAND2_X1  g0152(.A1(new_n282), .A2(new_n348), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT70), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n354), .A2(KEYINPUT12), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(KEYINPUT12), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n353), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n357), .B(KEYINPUT71), .C1(KEYINPUT12), .C2(new_n353), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n289), .A2(G68), .A3(new_n290), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n358), .B(new_n359), .C1(KEYINPUT71), .C2(new_n357), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n352), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n344), .A2(new_n347), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n345), .A2(new_n346), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT14), .B1(new_n364), .B2(new_n325), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n341), .A2(G179), .A3(new_n343), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT14), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n367), .B(G169), .C1(new_n345), .C2(new_n346), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n365), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n361), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n363), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n277), .B1(new_n256), .B2(G20), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n372), .A2(new_n289), .B1(new_n282), .B2(new_n277), .ZN(new_n373));
  AND2_X1   g0173(.A1(G58), .A2(G68), .ZN(new_n374));
  OAI21_X1  g0174(.A(G20), .B1(new_n374), .B2(new_n201), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT72), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g0177(.A(G58), .B(G68), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n378), .A2(KEYINPUT72), .A3(G20), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n274), .A2(G159), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n377), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  AND2_X1   g0181(.A1(KEYINPUT3), .A2(G33), .ZN(new_n382));
  NOR2_X1   g0182(.A1(KEYINPUT3), .A2(G33), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT7), .B1(new_n384), .B2(new_n223), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  NOR4_X1   g0186(.A1(new_n382), .A2(new_n383), .A3(new_n386), .A4(G20), .ZN(new_n387));
  OAI21_X1  g0187(.A(G68), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n381), .B1(new_n388), .B2(KEYINPUT73), .ZN(new_n389));
  OR2_X1    g0189(.A1(KEYINPUT3), .A2(G33), .ZN(new_n390));
  NAND2_X1  g0190(.A1(KEYINPUT3), .A2(G33), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n223), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n386), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n390), .A2(KEYINPUT7), .A3(new_n223), .A4(new_n391), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n348), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT73), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT16), .B1(new_n389), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n380), .B1(new_n375), .B2(new_n376), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT72), .B1(new_n378), .B2(G20), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n401), .A2(new_n388), .A3(KEYINPUT16), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n280), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n373), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n259), .B1(new_n214), .B2(new_n261), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G87), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n268), .A2(new_n264), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n208), .A2(G1698), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n407), .B(new_n408), .C1(new_n382), .C2(new_n383), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n270), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(G179), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n405), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n313), .A2(G232), .B1(new_n258), .B2(new_n255), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n409), .A2(new_n406), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n271), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n412), .B1(new_n416), .B2(G169), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n404), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT18), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT16), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n401), .B1(new_n395), .B2(new_n396), .ZN(new_n422));
  AOI211_X1 g0222(.A(KEYINPUT73), .B(new_n348), .C1(new_n393), .C2(new_n394), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n395), .A2(new_n381), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n425), .A2(KEYINPUT16), .B1(new_n222), .B2(new_n279), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n417), .B1(new_n427), .B2(new_n373), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT18), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n420), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n413), .A2(new_n415), .A3(G190), .ZN(new_n432));
  OAI21_X1  g0232(.A(G200), .B1(new_n405), .B2(new_n410), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n373), .B(new_n435), .C1(new_n398), .C2(new_n403), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT17), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n436), .B(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n431), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n329), .A2(new_n371), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT74), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n329), .A2(new_n439), .A3(new_n371), .A4(KEYINPUT74), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g0244(.A(G244), .B(new_n264), .C1(new_n382), .C2(new_n383), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT4), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n263), .A2(KEYINPUT4), .A3(G244), .A4(new_n264), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G283), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n263), .A2(G250), .A3(G1698), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n447), .A2(new_n448), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n271), .ZN(new_n452));
  INV_X1    g0252(.A(G45), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(G1), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT5), .B(G41), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n255), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AND2_X1   g0256(.A1(KEYINPUT5), .A2(G41), .ZN(new_n457));
  NOR2_X1   g0257(.A1(KEYINPUT5), .A2(G41), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n454), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n260), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(new_n216), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n452), .A2(new_n456), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n325), .ZN(new_n464));
  INV_X1    g0264(.A(G33), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(G1), .ZN(new_n466));
  OAI21_X1  g0266(.A(G97), .B1(new_n288), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n281), .A2(new_n215), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT76), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT76), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n467), .A2(new_n471), .A3(new_n468), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n274), .A2(G77), .ZN(new_n474));
  AND2_X1   g0274(.A1(G97), .A2(G107), .ZN(new_n475));
  NOR2_X1   g0275(.A1(G97), .A2(G107), .ZN(new_n476));
  OAI22_X1  g0276(.A1(new_n475), .A2(new_n476), .B1(KEYINPUT75), .B2(KEYINPUT6), .ZN(new_n477));
  OR2_X1    g0277(.A1(new_n475), .A2(new_n476), .ZN(new_n478));
  NOR2_X1   g0278(.A1(KEYINPUT75), .A2(KEYINPUT6), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(KEYINPUT6), .B2(new_n215), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n477), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n474), .B1(new_n481), .B2(new_n223), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n309), .B1(new_n393), .B2(new_n394), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n280), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n473), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n461), .B1(new_n451), .B2(new_n271), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(new_n411), .A3(new_n456), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n464), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n485), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT77), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n463), .A2(G200), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n452), .A2(G190), .A3(new_n456), .A4(new_n462), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n489), .A2(new_n490), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n492), .A2(new_n484), .A3(new_n473), .ZN(new_n494));
  INV_X1    g0294(.A(G200), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n495), .B1(new_n486), .B2(new_n456), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT77), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n488), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT21), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n288), .A2(new_n466), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G116), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n282), .A2(new_n209), .ZN(new_n502));
  AOI21_X1  g0302(.A(G20), .B1(G33), .B2(G283), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n465), .A2(G97), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n503), .A2(new_n504), .B1(G20), .B2(new_n209), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n280), .A2(KEYINPUT20), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT20), .B1(new_n280), .B2(new_n505), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n501), .B(new_n502), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G169), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n456), .B1(new_n460), .B2(new_n210), .ZN(new_n510));
  OAI211_X1 g0310(.A(G264), .B(G1698), .C1(new_n382), .C2(new_n383), .ZN(new_n511));
  OAI211_X1 g0311(.A(G257), .B(new_n264), .C1(new_n382), .C2(new_n383), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n390), .A2(G303), .A3(new_n391), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT80), .B1(new_n514), .B2(new_n271), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(KEYINPUT80), .A3(new_n271), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n510), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n499), .B1(new_n509), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n510), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n514), .A2(KEYINPUT80), .A3(new_n271), .ZN(new_n521));
  OAI211_X1 g0321(.A(G190), .B(new_n520), .C1(new_n521), .C2(new_n515), .ZN(new_n522));
  INV_X1    g0322(.A(new_n508), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n522), .B(new_n523), .C1(new_n518), .C2(new_n495), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n518), .A2(G179), .A3(new_n508), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n520), .B1(new_n521), .B2(new_n515), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n526), .A2(new_n508), .A3(KEYINPUT21), .A4(G169), .ZN(new_n527));
  AND4_X1   g0327(.A1(new_n519), .A2(new_n524), .A3(new_n525), .A4(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n263), .A2(G238), .A3(new_n264), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G116), .ZN(new_n530));
  OAI211_X1 g0330(.A(G244), .B(G1698), .C1(new_n382), .C2(new_n383), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n271), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n255), .A2(new_n454), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n256), .A2(G45), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n260), .A2(G250), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n533), .A2(G190), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT79), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(KEYINPUT78), .A2(KEYINPUT19), .ZN(new_n542));
  NOR2_X1   g0342(.A1(KEYINPUT78), .A2(KEYINPUT19), .ZN(new_n543));
  OAI211_X1 g0343(.A(G33), .B(G97), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(G87), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n544), .A2(new_n223), .B1(new_n545), .B2(new_n476), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n223), .B(G68), .C1(new_n382), .C2(new_n383), .ZN(new_n547));
  OR2_X1    g0347(.A1(new_n542), .A2(new_n543), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n276), .A2(new_n215), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n280), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n321), .A2(new_n282), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n500), .A2(G87), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n533), .A2(new_n538), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G200), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n537), .B1(new_n532), .B2(new_n271), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n557), .A2(KEYINPUT79), .A3(G190), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n541), .A2(new_n554), .A3(new_n556), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n411), .ZN(new_n560));
  INV_X1    g0360(.A(new_n321), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n500), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n551), .A2(new_n552), .A3(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n560), .B(new_n563), .C1(G169), .C2(new_n557), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n263), .A2(G257), .A3(G1698), .ZN(new_n566));
  NAND2_X1  g0366(.A1(G33), .A2(G294), .ZN(new_n567));
  OAI211_X1 g0367(.A(G250), .B(new_n264), .C1(new_n382), .C2(new_n383), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n271), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n459), .A2(G264), .A3(new_n260), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n571), .A2(new_n456), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n325), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT83), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n571), .A2(new_n456), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n271), .B2(new_n569), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n573), .A2(new_n574), .B1(new_n576), .B2(G179), .ZN(new_n577));
  OAI21_X1  g0377(.A(KEYINPUT83), .B1(new_n576), .B2(new_n325), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n223), .B(G87), .C1(new_n382), .C2(new_n383), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT22), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT22), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n263), .A2(new_n581), .A3(new_n223), .A4(G87), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT23), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(G20), .B2(new_n309), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n223), .A2(KEYINPUT23), .A3(G107), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n530), .A2(G20), .ZN(new_n587));
  AND2_X1   g0387(.A1(KEYINPUT81), .A2(KEYINPUT24), .ZN(new_n588));
  NOR4_X1   g0388(.A1(new_n585), .A2(new_n586), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  OR2_X1    g0389(.A1(KEYINPUT81), .A2(KEYINPUT24), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n583), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n591), .B1(new_n583), .B2(new_n589), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n280), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT25), .ZN(new_n595));
  AOI211_X1 g0395(.A(G107), .B(new_n281), .C1(KEYINPUT82), .C2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n595), .A2(KEYINPUT82), .ZN(new_n597));
  OR2_X1    g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n598), .A2(new_n599), .B1(new_n500), .B2(G107), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n577), .A2(new_n578), .B1(new_n594), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(G190), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n570), .A2(new_n572), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n576), .B2(G200), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n604), .A2(new_n594), .A3(new_n600), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n565), .A2(new_n601), .A3(new_n606), .ZN(new_n607));
  AND4_X1   g0407(.A1(new_n444), .A2(new_n498), .A3(new_n528), .A4(new_n607), .ZN(G372));
  NAND3_X1  g0408(.A1(new_n464), .A2(new_n485), .A3(new_n487), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT26), .B1(new_n565), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT26), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n554), .A2(new_n556), .A3(new_n539), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n488), .A2(new_n611), .A3(new_n564), .A4(new_n612), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n610), .A2(new_n613), .A3(new_n564), .ZN(new_n614));
  INV_X1    g0414(.A(new_n601), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n525), .A2(new_n527), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n616), .A3(new_n519), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n612), .A2(new_n564), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n606), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(new_n498), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n614), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n444), .A2(new_n621), .ZN(new_n622));
  AOI211_X1 g0422(.A(KEYINPUT18), .B(new_n417), .C1(new_n427), .C2(new_n373), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n429), .B1(new_n404), .B2(new_n418), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n328), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n626), .B1(new_n369), .B2(new_n370), .ZN(new_n627));
  XNOR2_X1  g0427(.A(new_n436), .B(KEYINPUT17), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n362), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n625), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n302), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n631), .A2(new_n307), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n622), .A2(new_n632), .ZN(G369));
  NAND2_X1  g0433(.A1(new_n616), .A2(new_n519), .ZN(new_n634));
  INV_X1    g0434(.A(G13), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n635), .A2(G1), .A3(G20), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT84), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n637), .A2(new_n638), .A3(KEYINPUT27), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n638), .B1(new_n637), .B2(KEYINPUT27), .ZN(new_n640));
  OAI221_X1 g0440(.A(G213), .B1(KEYINPUT27), .B2(new_n637), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(G343), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n634), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n615), .A2(new_n605), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n615), .B2(new_n643), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n648), .B(KEYINPUT85), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n643), .A2(new_n508), .ZN(new_n650));
  MUX2_X1   g0450(.A(new_n634), .B(new_n528), .S(new_n650), .Z(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G330), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n644), .B1(new_n594), .B2(new_n600), .ZN(new_n654));
  OAI22_X1  g0454(.A1(new_n646), .A2(new_n654), .B1(new_n615), .B2(new_n644), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n649), .A2(new_n657), .ZN(G399));
  INV_X1    g0458(.A(new_n228), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(G41), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n476), .A2(new_n545), .A3(new_n209), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n661), .A2(G1), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n225), .B2(new_n661), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT28), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n643), .B1(new_n614), .B2(new_n620), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT87), .ZN(new_n668));
  OR3_X1    g0468(.A1(new_n667), .A2(new_n668), .A3(KEYINPUT29), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT88), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n617), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n615), .A2(new_n616), .A3(KEYINPUT88), .A4(new_n519), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n671), .A2(new_n498), .A3(new_n619), .A4(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n488), .A2(new_n611), .A3(new_n564), .A4(new_n559), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT26), .B1(new_n618), .B2(new_n609), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n674), .A2(new_n564), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n643), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT29), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n668), .B1(new_n667), .B2(KEYINPUT29), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n669), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT30), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n486), .A2(new_n576), .A3(new_n557), .ZN(new_n682));
  OAI211_X1 g0482(.A(G179), .B(new_n520), .C1(new_n521), .C2(new_n515), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(G179), .B1(new_n570), .B2(new_n572), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n463), .A2(new_n526), .A3(new_n685), .A4(new_n555), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n682), .A2(new_n683), .A3(new_n681), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n643), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT31), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT86), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n607), .A2(new_n498), .A3(new_n528), .A4(new_n644), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI211_X1 g0495(.A(KEYINPUT31), .B(new_n643), .C1(new_n687), .C2(new_n688), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n692), .B1(new_n691), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(G330), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n680), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n666), .B1(new_n702), .B2(G1), .ZN(G364));
  NAND2_X1  g0503(.A1(new_n223), .A2(G13), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT89), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n453), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n706), .A2(new_n256), .A3(new_n660), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(KEYINPUT90), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(KEYINPUT90), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n653), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(G330), .B2(new_n651), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n222), .B1(G20), .B2(new_n325), .ZN(new_n714));
  NOR2_X1   g0514(.A1(G13), .A2(G33), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G20), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n263), .A2(new_n228), .ZN(new_n720));
  INV_X1    g0520(.A(G355), .ZN(new_n721));
  OAI22_X1  g0521(.A1(new_n720), .A2(new_n721), .B1(G116), .B2(new_n228), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n250), .A2(G45), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n659), .A2(new_n263), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n453), .B2(new_n226), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n722), .B1(new_n723), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n711), .B1(new_n719), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n223), .A2(G179), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(new_n602), .A3(G200), .ZN(new_n730));
  INV_X1    g0530(.A(G283), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n223), .A2(new_n411), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G190), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n729), .A2(new_n734), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI22_X1  g0538(.A1(G311), .A2(new_n736), .B1(new_n738), .B2(G329), .ZN(new_n739));
  INV_X1    g0539(.A(G322), .ZN(new_n740));
  INV_X1    g0540(.A(new_n733), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n495), .A2(G190), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n739), .B(new_n384), .C1(new_n740), .C2(new_n744), .ZN(new_n745));
  OR3_X1    g0545(.A1(new_n741), .A2(KEYINPUT91), .A3(new_n495), .ZN(new_n746));
  OAI21_X1  g0546(.A(KEYINPUT91), .B1(new_n741), .B2(new_n495), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n746), .A2(G190), .A3(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI211_X1 g0549(.A(new_n732), .B(new_n745), .C1(G326), .C2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n746), .A2(new_n602), .A3(new_n747), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  XNOR2_X1  g0552(.A(KEYINPUT33), .B(G317), .ZN(new_n753));
  OAI21_X1  g0553(.A(G20), .B1(new_n742), .B2(G179), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT93), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n752), .A2(new_n753), .B1(new_n759), .B2(G294), .ZN(new_n760));
  INV_X1    g0560(.A(G303), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n729), .A2(G190), .A3(G200), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n762), .A2(KEYINPUT92), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(KEYINPUT92), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT94), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n750), .B(new_n760), .C1(new_n761), .C2(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G50), .A2(new_n749), .B1(new_n752), .B2(G68), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n263), .B1(new_n266), .B2(new_n735), .C1(new_n744), .C2(new_n213), .ZN(new_n770));
  INV_X1    g0570(.A(G159), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n737), .A2(KEYINPUT32), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(KEYINPUT32), .B1(new_n737), .B2(new_n771), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(new_n309), .B2(new_n730), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n770), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n765), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G87), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n759), .A2(G97), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n769), .A2(new_n775), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n768), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n728), .B1(new_n780), .B2(new_n714), .ZN(new_n781));
  INV_X1    g0581(.A(new_n717), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n781), .B1(new_n651), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n713), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(G396));
  NAND2_X1  g0585(.A1(new_n766), .A2(G107), .ZN(new_n786));
  INV_X1    g0586(.A(G294), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n744), .A2(new_n787), .B1(new_n735), .B2(new_n209), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n730), .A2(new_n545), .ZN(new_n789));
  INV_X1    g0589(.A(G311), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n384), .B1(new_n737), .B2(new_n790), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G283), .A2(new_n752), .B1(new_n749), .B2(G303), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n786), .A2(new_n792), .A3(new_n778), .A4(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G143), .A2(new_n743), .B1(new_n736), .B2(G159), .ZN(new_n795));
  INV_X1    g0595(.A(G137), .ZN(new_n796));
  INV_X1    g0596(.A(G150), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n795), .B1(new_n748), .B2(new_n796), .C1(new_n797), .C2(new_n751), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT34), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G132), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n263), .B1(new_n737), .B2(new_n801), .C1(new_n730), .C2(new_n348), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(new_n759), .B2(G58), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n800), .B(new_n803), .C1(new_n202), .C2(new_n767), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n798), .A2(new_n799), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n794), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT96), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n806), .A2(new_n807), .ZN(new_n810));
  INV_X1    g0610(.A(new_n714), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n714), .A2(new_n715), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n710), .B1(new_n266), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT95), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n327), .A2(new_n643), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n324), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n328), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n626), .A2(new_n644), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n815), .B1(new_n821), .B2(new_n716), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n812), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n667), .B(new_n821), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n701), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n711), .B1(new_n701), .B2(new_n824), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G384));
  INV_X1    g0628(.A(KEYINPUT102), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n341), .A2(new_n343), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n367), .B1(new_n830), .B2(G169), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n368), .A2(new_n366), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n370), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n370), .A2(new_n643), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n833), .A2(new_n362), .A3(new_n834), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n370), .B(new_n643), .C1(new_n369), .C2(new_n363), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n820), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n691), .A2(new_n696), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n694), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n837), .A2(new_n839), .A3(KEYINPUT101), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(KEYINPUT101), .B1(new_n837), .B2(new_n839), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n421), .B1(new_n395), .B2(new_n381), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n426), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n641), .B1(new_n844), .B2(new_n373), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n431), .B2(new_n438), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n417), .B1(new_n844), .B2(new_n373), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT37), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n847), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n641), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n404), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n419), .A2(new_n851), .A3(new_n436), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n849), .A2(new_n436), .B1(new_n852), .B2(new_n848), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n846), .A2(new_n853), .A3(KEYINPUT38), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT38), .B1(new_n846), .B2(new_n853), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g0656(.A1(new_n841), .A2(new_n842), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n829), .B1(new_n857), .B2(KEYINPUT40), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n837), .A2(new_n839), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT101), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n855), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n846), .A2(new_n853), .A3(KEYINPUT38), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n861), .A2(new_n864), .A3(new_n840), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT40), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n865), .A2(KEYINPUT102), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n858), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n641), .B1(new_n427), .B2(new_n373), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT99), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT37), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n373), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n872), .B(new_n434), .C1(new_n424), .C2(new_n426), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n428), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n871), .A2(new_n874), .A3(new_n851), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n848), .B1(new_n851), .B2(KEYINPUT99), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n852), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT100), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT100), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n875), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n851), .B1(new_n625), .B2(new_n628), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n879), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  XOR2_X1   g0684(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n885));
  AOI21_X1  g0685(.A(new_n854), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OR3_X1    g0686(.A1(new_n886), .A2(new_n866), .A3(new_n859), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n868), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n444), .A2(new_n839), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(G330), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n889), .B2(new_n888), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n819), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n667), .B2(new_n821), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n835), .A2(new_n836), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NOR3_X1   g0697(.A1(new_n856), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n431), .B2(new_n641), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT39), .ZN(new_n900));
  INV_X1    g0700(.A(new_n885), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n882), .B1(new_n878), .B2(KEYINPUT100), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n901), .B1(new_n902), .B2(new_n881), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n900), .B1(new_n903), .B2(new_n854), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n369), .A2(new_n370), .A3(new_n644), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n856), .A2(KEYINPUT39), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n904), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n899), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n444), .A2(new_n669), .A3(new_n679), .A4(new_n678), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n910), .A2(new_n632), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n909), .B(new_n911), .Z(new_n912));
  AOI22_X1  g0712(.A1(new_n893), .A2(new_n912), .B1(G1), .B2(new_n705), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n912), .B2(new_n893), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT35), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n481), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n916), .A2(G116), .A3(new_n224), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n915), .B2(new_n481), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n918), .A2(KEYINPUT36), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(KEYINPUT36), .ZN(new_n920));
  OAI21_X1  g0720(.A(G77), .B1(new_n213), .B2(new_n348), .ZN(new_n921));
  OAI22_X1  g0721(.A1(new_n921), .A2(new_n225), .B1(G50), .B2(new_n348), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(G1), .A3(new_n635), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT97), .Z(new_n924));
  NAND4_X1  g0724(.A1(new_n914), .A2(new_n919), .A3(new_n920), .A4(new_n924), .ZN(G367));
  OAI21_X1  g0725(.A(new_n498), .B1(new_n489), .B2(new_n644), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n609), .B2(new_n644), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n928), .A2(new_n647), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n930), .A2(KEYINPUT42), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n493), .A2(new_n497), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n601), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n643), .B1(new_n933), .B2(new_n609), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(new_n930), .B2(KEYINPUT42), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n644), .A2(new_n554), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n618), .A2(new_n936), .ZN(new_n937));
  OR3_X1    g0737(.A1(new_n564), .A2(new_n644), .A3(new_n554), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n931), .A2(new_n935), .B1(KEYINPUT43), .B2(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n656), .A2(new_n928), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n944), .B(new_n945), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n660), .B(KEYINPUT41), .Z(new_n947));
  NAND2_X1  g0747(.A1(new_n649), .A2(new_n928), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT44), .Z(new_n949));
  NOR2_X1   g0749(.A1(new_n649), .A2(new_n928), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT45), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n657), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n645), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n647), .B1(new_n655), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n653), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n702), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n952), .A2(new_n657), .ZN(new_n959));
  OR3_X1    g0759(.A1(new_n954), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n947), .B1(new_n960), .B2(new_n702), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n706), .A2(new_n256), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n946), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n718), .B1(new_n228), .B2(new_n321), .C1(new_n237), .C2(new_n725), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n965), .A2(KEYINPUT103), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(KEYINPUT103), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n966), .A2(new_n967), .A3(new_n710), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n730), .A2(new_n215), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n263), .B1(new_n738), .B2(G317), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n970), .B1(new_n731), .B2(new_n735), .C1(new_n744), .C2(new_n761), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n969), .B(new_n971), .C1(G311), .C2(new_n749), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n766), .A2(KEYINPUT46), .A3(G116), .ZN(new_n973));
  XOR2_X1   g0773(.A(KEYINPUT104), .B(KEYINPUT46), .Z(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n765), .B2(new_n209), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n752), .A2(G294), .B1(new_n759), .B2(G107), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n972), .A2(new_n973), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  AOI22_X1  g0777(.A1(G143), .A2(new_n749), .B1(new_n752), .B2(G159), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n759), .A2(G68), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n743), .A2(G150), .B1(new_n738), .B2(G137), .ZN(new_n980));
  INV_X1    g0780(.A(new_n730), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(G77), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n384), .B1(new_n736), .B2(G50), .ZN(new_n983));
  AND3_X1   g0783(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n776), .A2(G58), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n978), .A2(new_n979), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n977), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT47), .Z(new_n988));
  OAI221_X1 g0788(.A(new_n968), .B1(new_n782), .B2(new_n939), .C1(new_n988), .C2(new_n811), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n964), .A2(new_n989), .ZN(G387));
  OAI22_X1  g0790(.A1(new_n720), .A2(new_n663), .B1(G107), .B2(new_n228), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n241), .A2(new_n453), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n277), .A2(G50), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT50), .ZN(new_n994));
  AOI211_X1 g0794(.A(G45), .B(new_n662), .C1(G68), .C2(G77), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n725), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n991), .B1(new_n992), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n711), .B1(new_n997), .B2(new_n719), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n752), .A2(new_n319), .B1(new_n776), .B2(G77), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n749), .A2(G159), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n263), .B1(new_n744), .B2(new_n202), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n735), .A2(new_n348), .B1(new_n737), .B2(new_n797), .ZN(new_n1002));
  NOR3_X1   g0802(.A1(new_n1001), .A2(new_n969), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n759), .A2(new_n561), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n999), .A2(new_n1000), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n263), .B1(new_n738), .B2(G326), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n731), .A2(new_n758), .B1(new_n765), .B2(new_n787), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G317), .A2(new_n743), .B1(new_n736), .B2(G303), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n748), .B2(new_n740), .C1(new_n790), .C2(new_n751), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT48), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1007), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n1010), .B2(new_n1009), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT49), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1006), .B1(new_n209), .B2(new_n730), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1005), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n998), .B1(new_n1016), .B2(new_n714), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n655), .B2(new_n782), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT105), .Z(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n957), .B2(new_n963), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n958), .A2(new_n660), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n702), .A2(new_n957), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(G393));
  OAI21_X1  g0823(.A(new_n958), .B1(new_n954), .B2(new_n959), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n960), .A2(new_n660), .A3(new_n1024), .ZN(new_n1025));
  NOR3_X1   g0825(.A1(new_n954), .A2(new_n962), .A3(new_n959), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n928), .A2(new_n717), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n245), .A2(new_n725), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n719), .B(new_n1028), .C1(G97), .C2(new_n659), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n748), .A2(new_n797), .B1(new_n771), .B2(new_n744), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT51), .ZN(new_n1031));
  INV_X1    g0831(.A(G143), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n263), .B1(new_n737), .B2(new_n1032), .C1(new_n735), .C2(new_n277), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n789), .B(new_n1033), .C1(new_n752), .C2(G50), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G77), .A2(new_n759), .B1(new_n776), .B2(G68), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1031), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n749), .A2(G317), .B1(G311), .B2(new_n743), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT52), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n263), .B1(new_n738), .B2(G322), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n309), .B2(new_n730), .C1(new_n765), .C2(new_n731), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1040), .A2(KEYINPUT106), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(KEYINPUT106), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n751), .A2(new_n761), .B1(new_n787), .B2(new_n735), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G116), .B2(new_n759), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1036), .B1(new_n1038), .B2(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT107), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n710), .B(new_n1029), .C1(new_n1047), .C2(new_n714), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1026), .B1(new_n1027), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1025), .A2(new_n1049), .ZN(G390));
  AOI21_X1  g0850(.A(new_n699), .B1(new_n838), .B2(new_n694), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n444), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n910), .A2(new_n632), .A3(new_n1052), .ZN(new_n1053));
  OAI211_X1 g0853(.A(G330), .B(new_n821), .C1(new_n695), .C2(new_n697), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n897), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1051), .A2(new_n837), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n621), .A2(new_n644), .A3(new_n821), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n819), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1057), .A2(KEYINPUT109), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT109), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1054), .A2(new_n897), .B1(new_n837), .B2(new_n1051), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1061), .B1(new_n1062), .B2(new_n895), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1054), .A2(new_n897), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n677), .A2(new_n818), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1051), .A2(new_n821), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n897), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1066), .A2(new_n819), .A3(new_n1067), .A4(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1053), .B1(new_n1064), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n906), .B1(new_n1059), .B2(new_n896), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n904), .B2(new_n907), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n905), .B1(new_n903), .B2(new_n854), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n897), .B1(new_n1067), .B2(new_n819), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n837), .B(new_n1051), .C1(new_n1073), .C2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1066), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1078), .A2(new_n1073), .A3(KEYINPUT108), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT108), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n907), .B1(new_n886), .B2(KEYINPUT39), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1072), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n884), .A2(new_n885), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n906), .B1(new_n1084), .B2(new_n863), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n818), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n643), .B(new_n1086), .C1(new_n673), .C2(new_n676), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n896), .B1(new_n1087), .B2(new_n894), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1065), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1080), .B1(new_n1083), .B2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1071), .B(new_n1077), .C1(new_n1079), .C2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(KEYINPUT110), .ZN(new_n1092));
  OAI21_X1  g0892(.A(KEYINPUT108), .B1(new_n1078), .B2(new_n1073), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1083), .A2(new_n1089), .A3(new_n1080), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT110), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1095), .A2(new_n1096), .A3(new_n1077), .A4(new_n1071), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1092), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1095), .A2(new_n1077), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1071), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n661), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1099), .A2(new_n962), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n813), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n765), .A2(new_n797), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT53), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n749), .A2(G128), .ZN(new_n1107));
  INV_X1    g0907(.A(G125), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n263), .B1(new_n737), .B2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(KEYINPUT54), .B(G143), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n744), .A2(new_n801), .B1(new_n735), .B2(new_n1110), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1109), .B(new_n1111), .C1(G50), .C2(new_n981), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n752), .A2(G137), .B1(new_n759), .B2(G159), .ZN(new_n1113));
  AND4_X1   g0913(.A1(new_n1106), .A2(new_n1107), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n263), .B1(new_n766), .B2(G87), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT111), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(G116), .A2(new_n743), .B1(new_n736), .B2(G97), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n1117), .B1(new_n348), .B2(new_n730), .C1(new_n787), .C2(new_n737), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n309), .A2(new_n751), .B1(new_n748), .B2(new_n731), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1118), .B(new_n1119), .C1(G77), .C2(new_n759), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1114), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n711), .B1(new_n319), .B2(new_n1104), .C1(new_n1121), .C2(new_n811), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n1081), .B2(new_n715), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1103), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1102), .A2(new_n1124), .ZN(G378));
  AND3_X1   g0925(.A1(new_n865), .A2(KEYINPUT102), .A3(new_n866), .ZN(new_n1126));
  AOI21_X1  g0926(.A(KEYINPUT102), .B1(new_n865), .B2(new_n866), .ZN(new_n1127));
  OAI211_X1 g0927(.A(G330), .B(new_n887), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n302), .A2(new_n307), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n850), .A2(new_n292), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1129), .B(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1131), .B(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1128), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n868), .A2(G330), .A3(new_n887), .A4(new_n1133), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT116), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n909), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n909), .ZN(new_n1140));
  AOI211_X1 g0940(.A(KEYINPUT116), .B(new_n1140), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n963), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1134), .A2(new_n715), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n711), .B1(G50), .B2(new_n1104), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1145));
  INV_X1    g0945(.A(G41), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1145), .B1(new_n384), .B2(new_n1146), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n751), .A2(new_n215), .B1(new_n765), .B2(new_n266), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n730), .A2(new_n213), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  AOI211_X1 g0950(.A(G41), .B(new_n263), .C1(new_n736), .C2(new_n561), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n743), .A2(G107), .B1(new_n738), .B2(G283), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n979), .A2(new_n1150), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1148), .B(new_n1153), .C1(G116), .C2(new_n749), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT112), .Z(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT113), .B(KEYINPUT58), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1147), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n751), .A2(new_n801), .B1(new_n796), .B2(new_n735), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT114), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1110), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n776), .A2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT115), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n749), .A2(G125), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n759), .A2(G150), .B1(G128), .B2(new_n743), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1159), .A2(new_n1162), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1165), .A2(KEYINPUT59), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(KEYINPUT59), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n981), .A2(G159), .ZN(new_n1168));
  AOI211_X1 g0968(.A(G33), .B(G41), .C1(new_n738), .C2(G124), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1157), .B1(new_n1166), .B2(new_n1170), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1144), .B1(new_n1171), .B2(new_n714), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1143), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1142), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT57), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1053), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1175), .B1(new_n1098), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1137), .A2(new_n909), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1135), .A2(new_n1136), .A3(new_n1140), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n661), .B1(new_n1177), .B2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1053), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1175), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1174), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(G375));
  NAND2_X1  g0986(.A1(new_n1064), .A2(new_n1070), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n1053), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n947), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(new_n1190), .A3(new_n1100), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT117), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n897), .A2(new_n715), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1004), .B1(new_n731), .B2(new_n744), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT118), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n263), .B1(new_n738), .B2(G303), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1196), .B(new_n982), .C1(new_n309), .C2(new_n735), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n751), .A2(new_n209), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(G294), .C2(new_n749), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1195), .B(new_n1199), .C1(new_n215), .C2(new_n767), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(G150), .A2(new_n736), .B1(new_n738), .B2(G128), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1201), .B(new_n263), .C1(new_n796), .C2(new_n744), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1149), .B(new_n1202), .C1(new_n752), .C2(new_n1160), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n749), .A2(G132), .B1(new_n759), .B2(G50), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(new_n771), .C2(new_n767), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n811), .B1(new_n1200), .B2(new_n1205), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n710), .B(new_n1206), .C1(new_n348), .C2(new_n813), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT119), .Z(new_n1208));
  AOI22_X1  g1008(.A1(new_n1187), .A2(new_n963), .B1(new_n1193), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1192), .A2(new_n1209), .ZN(G381));
  INV_X1    g1010(.A(G390), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n827), .ZN(new_n1212));
  NOR4_X1   g1012(.A1(new_n1212), .A2(G387), .A3(G396), .A4(G393), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT120), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1102), .A2(new_n1214), .A3(new_n1124), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1214), .B1(new_n1102), .B2(new_n1124), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(G375), .A2(new_n1218), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1213), .A2(new_n1219), .A3(new_n1209), .A4(new_n1192), .ZN(G407));
  INV_X1    g1020(.A(G213), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1221), .A2(G343), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1219), .A2(new_n1222), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT121), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1224), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1025(.A(KEYINPUT126), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1222), .A2(G2897), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1100), .A2(KEYINPUT60), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1228), .A2(new_n1189), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n660), .B1(new_n1228), .B2(new_n1189), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1209), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n827), .ZN(new_n1232));
  OAI211_X1 g1032(.A(G384), .B(new_n1209), .C1(new_n1229), .C2(new_n1230), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1234), .A2(KEYINPUT123), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT123), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1227), .B1(new_n1235), .B2(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1237), .A2(new_n1227), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT116), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(new_n909), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1098), .A2(new_n1176), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1242), .A2(new_n1190), .A3(new_n1243), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1180), .A2(new_n963), .B1(new_n1143), .B2(new_n1172), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1185), .A2(G378), .B1(new_n1217), .B2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(KEYINPUT125), .B1(new_n1247), .B2(new_n1222), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1174), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1243), .A2(KEYINPUT57), .A3(new_n1180), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n660), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT57), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1249), .B(G378), .C1(new_n1251), .C2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G378), .A2(KEYINPUT120), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1102), .A2(new_n1214), .A3(new_n1124), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1182), .A2(new_n947), .A3(new_n1183), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1245), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1254), .B(new_n1255), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1253), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT125), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1222), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1240), .B1(new_n1248), .B2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1226), .B1(new_n1263), .B2(KEYINPUT61), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1240), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1260), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1266));
  AOI211_X1 g1066(.A(KEYINPUT125), .B(new_n1222), .C1(new_n1253), .C2(new_n1258), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1265), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT61), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(KEYINPUT126), .A3(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT62), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1271), .B1(new_n1272), .B2(new_n1234), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1234), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1248), .A2(new_n1274), .A3(new_n1262), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1273), .B1(new_n1275), .B2(new_n1271), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1264), .A2(new_n1270), .A3(new_n1276), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(G393), .B(new_n784), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G390), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(G390), .A2(new_n1278), .ZN(new_n1281));
  OAI21_X1  g1081(.A(G387), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  OR2_X1    g1082(.A1(G390), .A2(new_n1278), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1283), .A2(new_n964), .A3(new_n989), .A4(new_n1279), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(KEYINPUT127), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1277), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1282), .A2(new_n1284), .A3(new_n1269), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT124), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1282), .A2(new_n1284), .A3(KEYINPUT124), .A4(new_n1269), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(new_n1290), .A2(new_n1291), .B1(new_n1265), .B2(new_n1272), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1248), .A2(KEYINPUT63), .A3(new_n1262), .A4(new_n1274), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1272), .A2(new_n1234), .ZN(new_n1294));
  XOR2_X1   g1094(.A(KEYINPUT122), .B(KEYINPUT63), .Z(new_n1295));
  OAI211_X1 g1095(.A(new_n1292), .B(new_n1293), .C1(new_n1294), .C2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1287), .A2(new_n1296), .ZN(G405));
  OAI21_X1  g1097(.A(new_n1253), .B1(new_n1218), .B2(new_n1185), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1298), .B(new_n1234), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1299), .B(new_n1285), .ZN(G402));
endmodule


