//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(KEYINPUT64), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n223), .A2(KEYINPUT64), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n212), .B(new_n217), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT65), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G68), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NOR2_X1   g0048(.A1(G20), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G150), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT8), .B(G58), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n207), .A2(G33), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G50), .A2(G58), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n207), .B1(new_n254), .B2(new_n219), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n215), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(new_n258), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n206), .A2(G20), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G50), .A3(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(G50), .B2(new_n261), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  OR2_X1    g0067(.A1(new_n267), .A2(KEYINPUT9), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  INV_X1    g0069(.A(G45), .ZN(new_n270));
  AOI21_X1  g0070(.A(G1), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(G1), .A3(G13), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(new_n273), .A3(G274), .ZN(new_n274));
  INV_X1    g0074(.A(G226), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n274), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  OR2_X1    g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  AOI21_X1  g0080(.A(G1698), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NOR2_X1   g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n281), .A2(G222), .B1(new_n284), .B2(G77), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n286), .B1(new_n279), .B2(new_n280), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  XOR2_X1   g0088(.A(KEYINPUT66), .B(G223), .Z(new_n289));
  OAI21_X1  g0089(.A(new_n285), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n278), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G200), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(G190), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n267), .A2(KEYINPUT9), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n268), .A2(new_n294), .A3(new_n295), .A4(new_n296), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT10), .ZN(new_n298));
  INV_X1    g0098(.A(G179), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n292), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  OAI22_X1  g0101(.A1(new_n292), .A2(G169), .B1(new_n260), .B2(new_n266), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n251), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n305), .A2(new_n249), .B1(G20), .B2(G77), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT15), .B(G87), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n306), .B1(new_n252), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n258), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n264), .A2(G77), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n263), .A2(new_n311), .B1(new_n221), .B2(new_n262), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n287), .A2(G238), .B1(new_n284), .B2(G107), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n281), .A2(G232), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n273), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n274), .B1(new_n222), .B2(new_n277), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n313), .B1(new_n318), .B2(G169), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n316), .A2(G179), .A3(new_n317), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n313), .B1(new_n318), .B2(G190), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n293), .B2(new_n318), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n304), .A2(new_n325), .ZN(new_n326));
  OAI211_X1 g0126(.A(G232), .B(G1698), .C1(new_n282), .C2(new_n283), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT67), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT3), .B(G33), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT67), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n329), .A2(new_n330), .A3(G232), .A4(G1698), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g0132(.A(G226), .B(new_n286), .C1(new_n282), .C2(new_n283), .ZN(new_n333));
  NAND2_X1  g0133(.A1(G33), .A2(G97), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n273), .B1(new_n332), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n274), .B1(new_n220), .B2(new_n277), .ZN(new_n338));
  OAI21_X1  g0138(.A(KEYINPUT13), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n338), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT13), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n335), .B1(new_n331), .B2(new_n328), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n340), .B(new_n341), .C1(new_n342), .C2(new_n273), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT14), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(new_n345), .A3(G169), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT70), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n344), .A2(G169), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT14), .ZN(new_n349));
  INV_X1    g0149(.A(G169), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n350), .B1(new_n339), .B2(new_n343), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT70), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(new_n352), .A3(new_n345), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n339), .A2(new_n343), .A3(G179), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n347), .A2(new_n349), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT69), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n249), .A2(G50), .B1(G20), .B2(new_n219), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n221), .B2(new_n252), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(KEYINPUT11), .A3(new_n258), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n206), .A2(new_n219), .A3(G13), .A4(G20), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT12), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n263), .A2(G68), .A3(new_n264), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n359), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT11), .B1(new_n358), .B2(new_n258), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n356), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n362), .A2(new_n361), .ZN(new_n366));
  INV_X1    g0166(.A(new_n364), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT69), .A4(new_n359), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n355), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n339), .A2(new_n343), .A3(G190), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT68), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT68), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n339), .A2(new_n343), .A3(new_n374), .A4(G190), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n293), .B1(new_n339), .B2(new_n343), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n370), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n251), .B1(new_n206), .B2(G20), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n380), .A2(new_n263), .B1(new_n262), .B2(new_n251), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n249), .A2(G159), .ZN(new_n383));
  AND2_X1   g0183(.A1(G58), .A2(G68), .ZN(new_n384));
  NOR2_X1   g0184(.A1(G58), .A2(G68), .ZN(new_n385));
  OAI21_X1  g0185(.A(G20), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n383), .B1(new_n386), .B2(KEYINPUT72), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT72), .ZN(new_n388));
  XNOR2_X1  g0188(.A(G58), .B(G68), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n388), .B1(new_n389), .B2(G20), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT7), .B1(new_n329), .B2(G20), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n284), .A2(new_n393), .A3(new_n207), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n392), .A2(new_n394), .A3(G68), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT16), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n259), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT71), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(new_n392), .B2(new_n394), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n329), .A2(G20), .ZN(new_n401));
  NOR2_X1   g0201(.A1(KEYINPUT71), .A2(KEYINPUT7), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(G68), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n391), .B(KEYINPUT16), .C1(new_n400), .C2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n382), .B1(new_n398), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n275), .A2(G1698), .ZN(new_n407));
  OAI221_X1 g0207(.A(new_n407), .B1(G223), .B2(G1698), .C1(new_n282), .C2(new_n283), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G87), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n273), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n274), .B1(new_n233), .B2(new_n277), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(new_n350), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n410), .A2(new_n411), .A3(new_n299), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT18), .B1(new_n406), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n393), .B1(new_n284), .B2(new_n207), .ZN(new_n417));
  NOR4_X1   g0217(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT7), .A4(G20), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n417), .A2(new_n418), .A3(new_n219), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n386), .A2(KEYINPUT72), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n389), .A2(new_n388), .A3(G20), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(new_n421), .A3(new_n383), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n397), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n423), .A2(new_n405), .A3(new_n258), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n381), .ZN(new_n425));
  INV_X1    g0225(.A(new_n415), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT18), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n416), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT73), .ZN(new_n430));
  INV_X1    g0230(.A(G190), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n412), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n293), .B1(new_n410), .B2(new_n411), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT17), .B1(new_n406), .B2(new_n434), .ZN(new_n435));
  AND4_X1   g0235(.A1(KEYINPUT17), .A2(new_n424), .A3(new_n381), .A4(new_n434), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n430), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n424), .A2(new_n381), .A3(new_n434), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n406), .A2(KEYINPUT17), .A3(new_n434), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT73), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n429), .B1(new_n437), .B2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n326), .A2(new_n371), .A3(new_n379), .A4(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT77), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n269), .A2(KEYINPUT5), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n206), .A2(G45), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT5), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G41), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n450), .A2(KEYINPUT77), .A3(new_n206), .A4(G45), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n269), .A2(KEYINPUT5), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n448), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n453), .A2(KEYINPUT80), .A3(G270), .A4(new_n273), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n206), .B(G45), .C1(new_n269), .C2(KEYINPUT5), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n455), .A2(new_n445), .B1(KEYINPUT5), .B2(new_n269), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n456), .A2(G274), .A3(new_n273), .A4(new_n451), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n291), .B1(new_n456), .B2(new_n451), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT80), .B1(new_n459), .B2(G270), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n462), .B(new_n207), .C1(G33), .C2(new_n202), .ZN(new_n463));
  INV_X1    g0263(.A(G116), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G20), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n463), .A2(new_n258), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT20), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n466), .B(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n261), .A2(G116), .ZN(new_n469));
  INV_X1    g0269(.A(G33), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(G1), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n262), .A2(new_n258), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n469), .B1(new_n472), .B2(G116), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(G264), .B(G1698), .C1(new_n282), .C2(new_n283), .ZN(new_n475));
  OAI211_X1 g0275(.A(G257), .B(new_n286), .C1(new_n282), .C2(new_n283), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n279), .A2(G303), .A3(new_n280), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n299), .B1(new_n478), .B2(new_n291), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n461), .A2(new_n474), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n453), .A2(G270), .A3(new_n273), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT80), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n478), .A2(new_n291), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n483), .A2(new_n484), .A3(new_n457), .A4(new_n454), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT21), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n350), .B1(new_n468), .B2(new_n473), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n486), .B1(new_n485), .B2(new_n487), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n480), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n485), .A2(G200), .ZN(new_n491));
  INV_X1    g0291(.A(new_n458), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n492), .A2(G190), .A3(new_n484), .A4(new_n483), .ZN(new_n493));
  INV_X1    g0293(.A(new_n474), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n490), .A2(new_n495), .A3(KEYINPUT81), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT81), .ZN(new_n497));
  AND4_X1   g0297(.A1(new_n483), .A2(new_n492), .A3(new_n474), .A4(new_n479), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n485), .A2(new_n487), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT21), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n497), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n329), .A2(new_n207), .A3(G87), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT22), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT22), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n329), .A2(new_n508), .A3(new_n207), .A4(G87), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g0310(.A(KEYINPUT82), .B(KEYINPUT24), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT23), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(new_n203), .A3(G20), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT83), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n512), .B2(new_n203), .ZN(new_n516));
  AOI21_X1  g0316(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n517));
  OAI22_X1  g0317(.A1(new_n513), .A2(new_n514), .B1(new_n517), .B2(G20), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n510), .A2(new_n511), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n511), .B1(new_n510), .B2(new_n519), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n258), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(G257), .B(G1698), .C1(new_n282), .C2(new_n283), .ZN(new_n523));
  OAI211_X1 g0323(.A(G250), .B(new_n286), .C1(new_n282), .C2(new_n283), .ZN(new_n524));
  INV_X1    g0324(.A(G294), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n523), .B(new_n524), .C1(new_n470), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n291), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n453), .A2(G264), .A3(new_n273), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(new_n528), .A3(new_n457), .ZN(new_n529));
  OR2_X1    g0329(.A1(new_n529), .A2(new_n431), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n262), .A2(new_n203), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(KEYINPUT84), .A3(KEYINPUT25), .ZN(new_n532));
  XNOR2_X1  g0332(.A(KEYINPUT84), .B(KEYINPUT25), .ZN(new_n533));
  INV_X1    g0333(.A(new_n472), .ZN(new_n534));
  OAI221_X1 g0334(.A(new_n532), .B1(new_n531), .B2(new_n533), .C1(new_n534), .C2(new_n203), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n529), .A2(G200), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n522), .A2(new_n530), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n510), .A2(new_n519), .ZN(new_n539));
  INV_X1    g0339(.A(new_n511), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n510), .A2(new_n511), .A3(new_n519), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n535), .B1(new_n543), .B2(new_n258), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n529), .A2(new_n350), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(G179), .B2(new_n529), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n538), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n261), .A2(G97), .ZN(new_n548));
  XNOR2_X1  g0348(.A(new_n548), .B(KEYINPUT75), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n472), .A2(G97), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n392), .A2(new_n394), .A3(G107), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n249), .A2(G77), .ZN(new_n553));
  XNOR2_X1  g0353(.A(new_n553), .B(KEYINPUT74), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G97), .A2(G107), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT6), .B1(new_n204), .B2(new_n555), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n203), .A2(KEYINPUT6), .A3(G97), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n552), .B(new_n554), .C1(new_n207), .C2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n551), .B1(new_n559), .B2(new_n258), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n453), .A2(G257), .A3(new_n273), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n457), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(G250), .B(G1698), .C1(new_n282), .C2(new_n283), .ZN(new_n565));
  XNOR2_X1  g0365(.A(new_n565), .B(KEYINPUT76), .ZN(new_n566));
  OAI211_X1 g0366(.A(G244), .B(new_n286), .C1(new_n282), .C2(new_n283), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT4), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n329), .A2(KEYINPUT4), .A3(G244), .A4(new_n286), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(new_n462), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n291), .B1(new_n566), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n564), .A2(new_n572), .A3(new_n299), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n569), .A2(new_n570), .A3(new_n462), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT76), .ZN(new_n575));
  XNOR2_X1  g0375(.A(new_n565), .B(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n273), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n350), .B1(new_n577), .B2(new_n563), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n561), .A2(new_n573), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n564), .A2(new_n572), .A3(G190), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n567), .A2(new_n568), .B1(G33), .B2(G283), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT76), .B1(new_n287), .B2(G250), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n565), .A2(new_n575), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n581), .B(new_n570), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n563), .B1(new_n291), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n580), .B(new_n560), .C1(new_n585), .C2(new_n293), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n287), .A2(G244), .B1(G33), .B2(G116), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n281), .A2(G238), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n291), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT79), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n273), .A2(G250), .A3(new_n447), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT78), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n593), .A2(new_n594), .A3(new_n273), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n594), .B1(new_n593), .B2(new_n273), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n591), .B(new_n592), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n599));
  OAI21_X1  g0399(.A(KEYINPUT78), .B1(new_n291), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n593), .A2(new_n273), .A3(new_n594), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n591), .B1(new_n602), .B2(new_n592), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n299), .B(new_n590), .C1(new_n598), .C2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n329), .A2(new_n207), .A3(G68), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT19), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n207), .B1(new_n334), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(G87), .B2(new_n204), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n606), .B1(new_n252), .B2(new_n202), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n605), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n610), .A2(new_n258), .B1(new_n262), .B2(new_n307), .ZN(new_n611));
  OR2_X1    g0411(.A1(new_n534), .A2(new_n307), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n273), .B1(new_n587), .B2(new_n588), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT79), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n614), .B1(new_n616), .B2(new_n597), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n604), .B(new_n613), .C1(G169), .C2(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(G190), .B(new_n590), .C1(new_n598), .C2(new_n603), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n472), .A2(G87), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n611), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n619), .B(new_n622), .C1(new_n293), .C2(new_n617), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n579), .A2(new_n586), .A3(new_n618), .A4(new_n623), .ZN(new_n624));
  NOR4_X1   g0424(.A1(new_n444), .A2(new_n505), .A3(new_n547), .A4(new_n624), .ZN(G372));
  INV_X1    g0425(.A(new_n303), .ZN(new_n626));
  INV_X1    g0426(.A(new_n429), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n379), .A2(new_n321), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n371), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT73), .B1(new_n440), .B2(new_n441), .ZN(new_n630));
  INV_X1    g0430(.A(new_n442), .ZN(new_n631));
  OAI22_X1  g0431(.A1(new_n629), .A2(KEYINPUT87), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n355), .A2(new_n370), .B1(new_n379), .B2(new_n321), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT87), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n627), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n626), .B1(new_n636), .B2(new_n298), .ZN(new_n637));
  INV_X1    g0437(.A(new_n618), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n590), .B1(new_n598), .B2(new_n603), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n639), .A2(new_n350), .B1(new_n611), .B2(new_n612), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n621), .B1(new_n617), .B2(G190), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n639), .A2(G200), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n640), .A2(new_n604), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n561), .A2(new_n573), .A3(new_n578), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n638), .B1(new_n645), .B2(KEYINPUT26), .ZN(new_n646));
  XOR2_X1   g0446(.A(KEYINPUT86), .B(KEYINPUT26), .Z(new_n647));
  NAND3_X1  g0447(.A1(new_n643), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n544), .A2(new_n546), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT85), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n490), .A2(new_n650), .ZN(new_n651));
  OAI211_X1 g0451(.A(KEYINPUT85), .B(new_n480), .C1(new_n488), .C2(new_n489), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n643), .A2(new_n538), .A3(new_n579), .A4(new_n586), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n646), .B(new_n648), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n637), .B1(new_n444), .B2(new_n656), .ZN(G369));
  AND2_X1   g0457(.A1(new_n651), .A2(new_n652), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G213), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G343), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n494), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n658), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n505), .B2(new_n666), .ZN(new_n668));
  XOR2_X1   g0468(.A(KEYINPUT88), .B(G330), .Z(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n544), .A2(new_n665), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT89), .B1(new_n547), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n522), .A2(new_n536), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n673), .B(new_n545), .C1(G179), .C2(new_n529), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT89), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n664), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n674), .A2(new_n675), .A3(new_n538), .A4(new_n676), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n672), .B(new_n677), .C1(new_n674), .C2(new_n665), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n668), .A2(new_n670), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n490), .A2(new_n665), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(new_n672), .B2(new_n677), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n674), .A2(new_n664), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n679), .A2(new_n683), .ZN(G399));
  INV_X1    g0484(.A(new_n210), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G41), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n204), .A2(G87), .A3(G116), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G1), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n213), .B2(new_n687), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT28), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n651), .A2(new_n652), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n654), .B1(new_n692), .B2(new_n674), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n618), .A2(new_n623), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT26), .B1(new_n694), .B2(new_n579), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n695), .A2(new_n648), .A3(new_n618), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n665), .B1(new_n693), .B2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT29), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT91), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT91), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n697), .A2(new_n701), .A3(new_n698), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT26), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n644), .A2(new_n704), .A3(new_n618), .A4(new_n623), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n618), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n647), .B1(new_n643), .B2(new_n644), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT92), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n647), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n694), .B2(new_n579), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT92), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n710), .A2(new_n711), .A3(new_n618), .A4(new_n705), .ZN(new_n712));
  INV_X1    g0512(.A(new_n538), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n624), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n674), .A2(new_n502), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n708), .A2(new_n712), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(KEYINPUT29), .A3(new_n665), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n703), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT93), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n624), .A2(new_n547), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n721), .B(new_n665), .C1(new_n496), .C2(new_n504), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n529), .A2(new_n299), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n585), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT90), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n639), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n617), .A2(KEYINPUT90), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n724), .A2(new_n485), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n479), .A2(new_n527), .A3(new_n528), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n639), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n730), .A2(KEYINPUT30), .A3(new_n461), .A4(new_n585), .ZN(new_n731));
  INV_X1    g0531(.A(new_n729), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n585), .A2(new_n461), .A3(new_n617), .A4(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT30), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n728), .A2(new_n731), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT31), .B1(new_n736), .B2(new_n664), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n664), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n722), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n670), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OR3_X1    g0542(.A1(new_n719), .A2(new_n720), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n720), .B1(new_n719), .B2(new_n742), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n691), .B1(new_n745), .B2(G1), .ZN(G364));
  AND2_X1   g0546(.A1(new_n207), .A2(G13), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n206), .B1(new_n747), .B2(G45), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n686), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n750), .B1(new_n668), .B2(new_n670), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(new_n670), .B2(new_n668), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G13), .A2(G33), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n215), .B1(G20), .B2(new_n350), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n685), .A2(new_n284), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n758), .A2(G355), .B1(new_n464), .B2(new_n685), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n244), .A2(new_n270), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n685), .A2(new_n329), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(G45), .B2(new_n213), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n759), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT94), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n757), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(new_n764), .B2(new_n763), .ZN(new_n766));
  INV_X1    g0566(.A(new_n756), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n207), .A2(new_n299), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n769), .A2(new_n293), .A3(G190), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n769), .A2(G190), .A3(G200), .ZN(new_n771));
  AOI22_X1  g0571(.A1(G68), .A2(new_n770), .B1(new_n771), .B2(G77), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n207), .A2(G179), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(new_n431), .A3(G200), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n772), .B1(new_n203), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G87), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n773), .A2(G190), .A3(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n768), .A2(G190), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n293), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G50), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n329), .B1(new_n776), .B2(new_n777), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n778), .A2(G200), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G58), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G179), .A2(G200), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n207), .B1(new_n787), .B2(G190), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n202), .ZN(new_n789));
  NOR4_X1   g0589(.A1(new_n775), .A2(new_n782), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n787), .A2(G20), .A3(new_n431), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n791), .A2(KEYINPUT95), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(KEYINPUT95), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G159), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT32), .ZN(new_n797));
  AOI21_X1  g0597(.A(KEYINPUT96), .B1(new_n790), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n774), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n771), .A2(G311), .B1(G283), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G303), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n801), .B2(new_n777), .ZN(new_n802));
  XNOR2_X1  g0602(.A(KEYINPUT33), .B(G317), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n329), .B1(new_n770), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n788), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n783), .A2(G322), .B1(G294), .B2(new_n805), .ZN(new_n806));
  XOR2_X1   g0606(.A(KEYINPUT97), .B(G326), .Z(new_n807));
  OAI211_X1 g0607(.A(new_n804), .B(new_n806), .C1(new_n780), .C2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n794), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n802), .B(new_n808), .C1(G329), .C2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n798), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n790), .A2(KEYINPUT96), .A3(new_n797), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n767), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n750), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n766), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n755), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n668), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n752), .A2(new_n817), .ZN(G396));
  NOR2_X1   g0618(.A1(new_n322), .A2(new_n664), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n313), .A2(new_n664), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n324), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n322), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n697), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n325), .A2(new_n664), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n825), .B1(new_n656), .B2(new_n827), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n828), .A2(new_n741), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n750), .B1(new_n828), .B2(new_n741), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n756), .A2(new_n753), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n750), .B1(G77), .B2(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G150), .A2(new_n770), .B1(new_n771), .B2(G159), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n783), .A2(G143), .ZN(new_n836));
  INV_X1    g0636(.A(G137), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n835), .B(new_n836), .C1(new_n837), .C2(new_n780), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT34), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n774), .A2(new_n219), .B1(new_n777), .B2(new_n781), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(G58), .B2(new_n805), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(G132), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n329), .B1(new_n794), .B2(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT98), .ZN(new_n847));
  INV_X1    g0647(.A(new_n777), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n329), .B(new_n789), .C1(G107), .C2(new_n848), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n849), .B1(new_n525), .B2(new_n784), .C1(new_n801), .C2(new_n780), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n771), .A2(G116), .B1(G87), .B2(new_n799), .ZN(new_n851));
  INV_X1    g0651(.A(G283), .ZN(new_n852));
  INV_X1    g0652(.A(new_n770), .ZN(new_n853));
  INV_X1    g0653(.A(G311), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n851), .B1(new_n852), .B2(new_n853), .C1(new_n854), .C2(new_n794), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n844), .A2(new_n847), .B1(new_n850), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n834), .B1(new_n856), .B2(new_n756), .ZN(new_n857));
  INV_X1    g0657(.A(new_n824), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n857), .B1(new_n858), .B2(new_n754), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT99), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n831), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(G384));
  INV_X1    g0662(.A(new_n558), .ZN(new_n863));
  OR2_X1    g0663(.A1(new_n863), .A2(KEYINPUT35), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(KEYINPUT35), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n864), .A2(G116), .A3(new_n216), .A4(new_n865), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n866), .B(KEYINPUT36), .Z(new_n867));
  OAI211_X1 g0667(.A(new_n214), .B(G77), .C1(new_n785), .C2(new_n219), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n781), .A2(G68), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n206), .B(G13), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n819), .B1(new_n655), .B2(new_n826), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n370), .A2(new_n664), .ZN(new_n874));
  INV_X1    g0674(.A(new_n353), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n354), .B1(new_n351), .B2(new_n345), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n352), .B1(new_n351), .B2(new_n345), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n379), .B(new_n874), .C1(new_n878), .C2(new_n369), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n377), .B(new_n370), .C1(new_n373), .C2(new_n375), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n370), .B(new_n664), .C1(new_n355), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT71), .B1(new_n417), .B2(new_n418), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n284), .A2(new_n207), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n219), .B1(new_n884), .B2(new_n402), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n422), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n259), .B1(new_n886), .B2(KEYINPUT16), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n391), .B1(new_n400), .B2(new_n404), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n397), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n382), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n438), .B1(new_n890), .B2(new_n662), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n415), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT37), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n425), .A2(new_n426), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n662), .B(KEYINPUT100), .Z(new_n895));
  NAND2_X1  g0695(.A1(new_n425), .A2(new_n895), .ZN(new_n896));
  XOR2_X1   g0696(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n897));
  NAND4_X1  g0697(.A1(new_n894), .A2(new_n896), .A3(new_n438), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n890), .A2(new_n662), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(KEYINPUT38), .B(new_n899), .C1(new_n443), .C2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n899), .B1(new_n443), .B2(new_n901), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n873), .B(new_n882), .C1(new_n903), .C2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT39), .ZN(new_n908));
  INV_X1    g0708(.A(new_n898), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n416), .A2(new_n428), .A3(new_n440), .A4(new_n441), .ZN(new_n910));
  INV_X1    g0710(.A(new_n896), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n909), .A2(KEYINPUT102), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n894), .A2(new_n896), .A3(new_n438), .ZN(new_n913));
  INV_X1    g0713(.A(new_n897), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT102), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(new_n916), .A3(new_n898), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT38), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n908), .B1(new_n903), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n355), .A2(new_n370), .A3(new_n665), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n904), .A2(new_n905), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(KEYINPUT39), .A3(new_n902), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n919), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n627), .A2(new_n895), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n907), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n633), .A2(new_n634), .B1(new_n437), .B2(new_n442), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n629), .A2(KEYINPUT87), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n429), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n298), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n303), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n710), .A2(new_n618), .A3(new_n705), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n932), .A2(KEYINPUT92), .B1(new_n714), .B2(new_n715), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n664), .B1(new_n933), .B2(new_n712), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n444), .B1(KEYINPUT29), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n931), .B1(new_n703), .B2(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n926), .B(new_n936), .Z(new_n937));
  AOI21_X1  g0737(.A(new_n824), .B1(new_n879), .B2(new_n881), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n740), .B(new_n938), .C1(new_n903), .C2(new_n918), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n938), .A2(new_n740), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT40), .B1(new_n922), .B2(new_n902), .ZN(new_n941));
  AOI22_X1  g0741(.A1(KEYINPUT40), .A2(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AND4_X1   g0742(.A1(new_n371), .A2(new_n326), .A3(new_n379), .A4(new_n443), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n740), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n942), .B(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n945), .A2(new_n669), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n937), .A2(new_n946), .B1(new_n206), .B2(new_n747), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n937), .A2(new_n946), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n871), .B1(new_n947), .B2(new_n948), .ZN(G367));
  INV_X1    g0749(.A(new_n771), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n284), .B1(new_n202), .B2(new_n774), .C1(new_n950), .C2(new_n852), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(G317), .B2(new_n809), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n848), .A2(KEYINPUT46), .A3(G116), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT46), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n777), .B2(new_n464), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n953), .B(new_n955), .C1(new_n853), .C2(new_n525), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT108), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n784), .A2(new_n801), .B1(new_n788), .B2(new_n203), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(G311), .B2(new_n779), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n952), .A2(new_n958), .A3(new_n959), .A4(new_n961), .ZN(new_n962));
  AOI22_X1  g0762(.A1(G50), .A2(new_n771), .B1(new_n770), .B2(G159), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT109), .Z(new_n964));
  OAI21_X1  g0764(.A(new_n329), .B1(new_n777), .B2(new_n785), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(G77), .B2(new_n799), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n964), .B(new_n966), .C1(new_n837), .C2(new_n794), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n788), .A2(new_n219), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(new_n779), .B2(G143), .ZN(new_n969));
  INV_X1    g0769(.A(G150), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n969), .B1(new_n970), .B2(new_n784), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n962), .B1(new_n967), .B2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT47), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n756), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n621), .A2(new_n664), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT103), .Z(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n694), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n638), .B2(new_n976), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n755), .ZN(new_n979));
  INV_X1    g0779(.A(new_n761), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n757), .B1(new_n210), .B2(new_n307), .C1(new_n980), .C2(new_n239), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n974), .A2(new_n750), .A3(new_n979), .A4(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT106), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n560), .A2(new_n665), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n579), .A2(new_n586), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n578), .A2(new_n573), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n986), .B(KEYINPUT104), .C1(new_n987), .C2(new_n985), .ZN(new_n988));
  OR3_X1    g0788(.A1(new_n985), .A2(new_n987), .A3(KEYINPUT104), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n983), .B1(new_n683), .B2(new_n991), .ZN(new_n992));
  NOR4_X1   g0792(.A1(new_n681), .A2(new_n990), .A3(KEYINPUT106), .A4(new_n682), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT45), .ZN(new_n994));
  OR3_X1    g0794(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n990), .B1(new_n681), .B2(new_n682), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT44), .Z(new_n997));
  OAI21_X1  g0797(.A(new_n994), .B1(new_n992), .B2(new_n993), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n995), .A2(new_n997), .A3(new_n679), .A4(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(KEYINPUT107), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n995), .A2(new_n998), .A3(new_n997), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n679), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1001), .A2(KEYINPUT107), .A3(new_n1002), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n668), .A2(new_n670), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n681), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n680), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1008), .B1(new_n678), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1007), .B(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n745), .B1(new_n1006), .B2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n686), .B(KEYINPUT41), .Z(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n749), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT43), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n978), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n991), .A2(new_n681), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1018), .A2(KEYINPUT42), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT105), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n579), .B1(new_n990), .B2(new_n674), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1018), .A2(KEYINPUT42), .B1(new_n1021), .B2(new_n665), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1017), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n978), .A2(new_n1016), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n679), .A2(new_n990), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1027), .B(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n982), .B1(new_n1015), .B2(new_n1030), .ZN(G387));
  AOI21_X1  g0831(.A(new_n1011), .B1(new_n743), .B2(new_n744), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1032), .A2(new_n687), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1011), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1033), .B1(new_n745), .B2(new_n1034), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n678), .A2(new_n816), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n688), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n758), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(G107), .B2(new_n210), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n236), .A2(new_n270), .ZN(new_n1040));
  AOI211_X1 g0840(.A(G45), .B(new_n1037), .C1(G68), .C2(G77), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n251), .A2(G50), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n980), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1039), .B1(new_n1040), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n757), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n750), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n777), .A2(new_n221), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n771), .B2(G68), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n794), .B2(new_n970), .C1(new_n251), .C2(new_n853), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n329), .B1(new_n202), .B2(new_n774), .C1(new_n784), .C2(new_n781), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n780), .A2(new_n795), .B1(new_n788), .B2(new_n307), .ZN(new_n1053));
  NOR3_X1   g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT111), .Z(new_n1055));
  AOI21_X1  g0855(.A(new_n329), .B1(new_n799), .B2(G116), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n777), .A2(new_n525), .B1(new_n788), .B2(new_n852), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G303), .A2(new_n771), .B1(new_n770), .B2(G311), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n783), .A2(G317), .ZN(new_n1059));
  INV_X1    g0859(.A(G322), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1058), .B(new_n1059), .C1(new_n1060), .C2(new_n780), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT48), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1057), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n1062), .B2(new_n1061), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT49), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1056), .B1(new_n794), .B2(new_n807), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1055), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1048), .B1(new_n1068), .B2(new_n756), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1034), .A2(new_n749), .B1(new_n1036), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1035), .A2(new_n1070), .ZN(G393));
  OAI221_X1 g0871(.A(new_n757), .B1(new_n202), .B2(new_n210), .C1(new_n980), .C2(new_n247), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n329), .B1(new_n799), .B2(G107), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n950), .B2(new_n525), .C1(new_n801), .C2(new_n853), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G311), .A2(new_n783), .B1(new_n779), .B2(G317), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT52), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1074), .B(new_n1076), .C1(G116), .C2(new_n805), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n794), .A2(new_n1060), .B1(new_n852), .B2(new_n777), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT113), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G150), .A2(new_n779), .B1(new_n783), .B2(G159), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT51), .Z(new_n1081));
  NAND2_X1  g0881(.A1(new_n805), .A2(G77), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1082), .B(new_n329), .C1(new_n776), .C2(new_n774), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n771), .A2(new_n305), .B1(G68), .B2(new_n848), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n781), .B2(new_n853), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1083), .B(new_n1085), .C1(G143), .C2(new_n809), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1077), .A2(new_n1079), .B1(new_n1081), .B2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n750), .B(new_n1072), .C1(new_n1087), .C2(new_n767), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n990), .B2(new_n755), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT112), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n999), .A2(new_n1090), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(new_n1003), .Z(new_n1092));
  AOI21_X1  g0892(.A(new_n1089), .B1(new_n1092), .B2(new_n749), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1032), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n686), .B1(new_n1094), .B2(new_n1006), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1092), .A2(new_n1032), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1093), .B1(new_n1095), .B2(new_n1096), .ZN(G390));
  INV_X1    g0897(.A(G330), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n664), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1099), .A2(new_n737), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1098), .B1(new_n1100), .B2(new_n722), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n938), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n714), .B1(new_n658), .B2(new_n649), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n696), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n827), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n882), .B1(new_n1106), .B2(new_n819), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1107), .A2(new_n920), .B1(new_n919), .B2(new_n923), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n920), .B1(new_n903), .B2(new_n918), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n717), .A2(new_n665), .A3(new_n823), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n820), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1109), .B1(new_n1111), .B2(new_n882), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1103), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1109), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n819), .B1(new_n934), .B2(new_n823), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n882), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n919), .A2(new_n923), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n920), .B1(new_n872), .B2(new_n1116), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n740), .A2(new_n670), .A3(new_n858), .A4(new_n882), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1117), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1113), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1123), .A2(new_n748), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1118), .A2(new_n753), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n750), .B1(new_n305), .B2(new_n833), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT54), .B(G143), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n853), .A2(new_n837), .B1(new_n950), .B2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n284), .B(new_n1128), .C1(G50), .C2(new_n799), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n784), .A2(new_n845), .B1(new_n788), .B2(new_n795), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(G128), .B2(new_n779), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n809), .A2(G125), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n777), .A2(new_n970), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1133), .B(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1129), .A2(new_n1131), .A3(new_n1132), .A4(new_n1135), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1082), .B1(new_n780), .B2(new_n852), .C1(new_n464), .C2(new_n784), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n950), .A2(new_n202), .B1(new_n219), .B2(new_n774), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G107), .B2(new_n770), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n284), .B1(new_n777), .B2(new_n776), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT117), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1139), .B(new_n1141), .C1(new_n525), .C2(new_n794), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1136), .B1(new_n1137), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1126), .B1(new_n1143), .B2(new_n756), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT118), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1124), .B1(new_n1125), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT114), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n740), .A2(new_n670), .A3(new_n858), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1148), .A2(new_n1116), .B1(new_n938), .B2(new_n1101), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1121), .A2(new_n820), .A3(new_n1110), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n882), .B1(new_n1101), .B2(new_n858), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n1149), .A2(new_n872), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n943), .A2(new_n1101), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1152), .A2(new_n936), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1147), .B1(new_n1123), .B2(new_n1154), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1121), .A2(new_n820), .A3(new_n1110), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1151), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n669), .B(new_n824), .C1(new_n1100), .C2(new_n722), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1102), .B1(new_n1158), .B2(new_n882), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1156), .A2(new_n1157), .B1(new_n1159), .B2(new_n873), .ZN(new_n1160));
  AOI211_X1 g0960(.A(KEYINPUT91), .B(KEYINPUT29), .C1(new_n655), .C2(new_n665), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n701), .B1(new_n697), .B2(new_n698), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n943), .A2(new_n718), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n637), .B(new_n1153), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1160), .A2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1166), .A2(KEYINPUT114), .A3(new_n1122), .A4(new_n1113), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1155), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n687), .B1(new_n1123), .B2(new_n1154), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1168), .A2(KEYINPUT115), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(KEYINPUT115), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1146), .B1(new_n1170), .B2(new_n1171), .ZN(G378));
  INV_X1    g0972(.A(new_n1165), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1168), .A2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n267), .A2(new_n662), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n304), .B(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1177), .B(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n942), .B2(new_n1098), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n940), .A2(new_n941), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT40), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n918), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n902), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1183), .B1(new_n940), .B2(new_n1185), .ZN(new_n1186));
  OAI211_X1 g0986(.A(G330), .B(new_n1179), .C1(new_n1182), .C2(new_n1186), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1181), .A2(new_n1187), .A3(new_n926), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n926), .B1(new_n1181), .B2(new_n1187), .ZN(new_n1189));
  OAI21_X1  g0989(.A(KEYINPUT57), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT121), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1174), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT57), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1165), .B1(new_n1155), .B2(new_n1167), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1194), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(KEYINPUT121), .B1(new_n1195), .B2(new_n1190), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1193), .A2(new_n1197), .A3(new_n1198), .A4(new_n686), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n814), .B1(new_n781), .B2(new_n832), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n783), .A2(G128), .B1(G150), .B2(new_n805), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n770), .A2(G132), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1203), .B1(new_n777), .B2(new_n1127), .C1(new_n950), .C2(new_n837), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1202), .B(new_n1204), .C1(G125), .C2(new_n779), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n809), .A2(G124), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n470), .A2(new_n269), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT119), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G159), .B2(new_n799), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .A4(new_n1212), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n950), .A2(new_n307), .B1(new_n785), .B2(new_n774), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G97), .B2(new_n770), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n852), .B2(new_n794), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n284), .A2(new_n269), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1049), .A2(new_n1217), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n784), .A2(new_n203), .B1(new_n780), .B2(new_n464), .ZN(new_n1219));
  NOR4_X1   g1019(.A1(new_n1216), .A2(new_n968), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1220), .A2(KEYINPUT58), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(KEYINPUT58), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1211), .A2(new_n781), .A3(new_n1217), .ZN(new_n1223));
  AND4_X1   g1023(.A1(new_n1213), .A2(new_n1221), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1200), .B1(new_n767), .B2(new_n1224), .C1(new_n1179), .C2(new_n754), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n1196), .B2(new_n748), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT120), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1226), .B(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1199), .A2(new_n1228), .ZN(G375));
  NAND2_X1  g1029(.A1(new_n1160), .A2(new_n1165), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1154), .A2(new_n1230), .A3(new_n1014), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1152), .A2(new_n749), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1116), .A2(new_n753), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT122), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n814), .B1(new_n219), .B2(new_n832), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G107), .A2(new_n771), .B1(new_n770), .B2(G116), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n525), .B2(new_n780), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT123), .Z(new_n1238));
  OAI221_X1 g1038(.A(new_n284), .B1(new_n777), .B2(new_n202), .C1(new_n221), .C2(new_n774), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n784), .A2(new_n852), .B1(new_n788), .B2(new_n307), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1239), .B(new_n1240), .C1(G303), .C2(new_n809), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n329), .B1(new_n774), .B2(new_n785), .ZN(new_n1242));
  XOR2_X1   g1042(.A(new_n1242), .B(KEYINPUT124), .Z(new_n1243));
  AOI22_X1  g1043(.A1(new_n783), .A2(G137), .B1(G50), .B2(new_n805), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n845), .B2(new_n780), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n771), .A2(G150), .B1(G159), .B2(new_n848), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n853), .B2(new_n1127), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1245), .B(new_n1247), .C1(G128), .C2(new_n809), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1238), .A2(new_n1241), .B1(new_n1243), .B2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1234), .B(new_n1235), .C1(new_n767), .C2(new_n1249), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1232), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1231), .A2(new_n1251), .ZN(G381));
  NOR2_X1   g1052(.A1(G393), .A2(G396), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1254), .A2(new_n1146), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1256));
  NOR4_X1   g1056(.A1(new_n1256), .A2(G384), .A3(G390), .A4(G381), .ZN(new_n1257));
  INV_X1    g1057(.A(G387), .ZN(new_n1258));
  INV_X1    g1058(.A(G375), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(G407));
  NAND2_X1  g1060(.A1(new_n1254), .A2(new_n1146), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n663), .A2(G213), .ZN(new_n1262));
  OR3_X1    g1062(.A1(G375), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(G407), .A2(G213), .A3(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT125), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(G407), .A2(new_n1263), .A3(KEYINPUT125), .A4(G213), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(G409));
  XNOR2_X1  g1068(.A(G387), .B(G390), .ZN(new_n1269));
  AND2_X1   g1069(.A1(G393), .A2(G396), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1270), .A2(new_n1253), .ZN(new_n1271));
  XOR2_X1   g1071(.A(new_n1269), .B(new_n1271), .Z(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT60), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1230), .B1(new_n1166), .B2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1160), .A2(new_n1165), .A3(KEYINPUT60), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1275), .A2(new_n686), .A3(new_n1276), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1277), .A2(G384), .A3(new_n1251), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G384), .B1(new_n1277), .B2(new_n1251), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1199), .A2(new_n1228), .A3(G378), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1196), .B1(new_n1168), .B2(new_n1173), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1226), .B1(new_n1282), .B2(new_n1014), .ZN(new_n1283));
  OAI21_X1  g1083(.A(KEYINPUT126), .B1(new_n1283), .B2(new_n1261), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT126), .ZN(new_n1285));
  NOR3_X1   g1085(.A1(new_n1195), .A2(new_n1013), .A3(new_n1196), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1255), .B(new_n1285), .C1(new_n1226), .C2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1284), .A2(new_n1287), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1262), .B(new_n1280), .C1(new_n1281), .C2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT127), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1199), .A2(new_n1228), .A3(G378), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(new_n1284), .A3(new_n1287), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1293), .A2(KEYINPUT127), .A3(new_n1262), .A4(new_n1280), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT62), .B1(new_n1291), .B2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1262), .B1(new_n1281), .B2(new_n1288), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n663), .A2(G213), .A3(G2897), .ZN(new_n1297));
  XOR2_X1   g1097(.A(new_n1280), .B(new_n1297), .Z(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT61), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1289), .A2(KEYINPUT62), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1273), .B1(new_n1295), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT63), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1291), .A2(new_n1303), .A3(new_n1294), .ZN(new_n1304));
  OR2_X1    g1104(.A1(new_n1289), .A2(new_n1303), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1304), .A2(new_n1272), .A3(new_n1299), .A4(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1302), .A2(new_n1306), .ZN(G405));
  NOR2_X1   g1107(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1308));
  OR3_X1    g1108(.A1(new_n1308), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1280), .B1(new_n1308), .B2(new_n1281), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1273), .A2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1272), .A2(new_n1310), .A3(new_n1309), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(G402));
endmodule


