

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U552 ( .A1(n700), .A2(n699), .ZN(n702) );
  XNOR2_X1 U553 ( .A(n724), .B(n723), .ZN(n728) );
  AND2_X1 U554 ( .A1(n750), .A2(n741), .ZN(n743) );
  AND2_X1 U555 ( .A1(n765), .A2(n763), .ZN(n764) );
  INV_X1 U556 ( .A(KEYINPUT33), .ZN(n763) );
  INV_X1 U557 ( .A(n995), .ZN(n771) );
  INV_X1 U558 ( .A(n553), .ZN(n894) );
  AND2_X1 U559 ( .A1(n523), .A2(n827), .ZN(n520) );
  AND2_X1 U560 ( .A1(n729), .A2(G1341), .ZN(n521) );
  XOR2_X1 U561 ( .A(G2104), .B(KEYINPUT66), .Z(n522) );
  AND2_X1 U562 ( .A1(n808), .A2(n822), .ZN(n523) );
  AND2_X1 U563 ( .A1(n784), .A2(n783), .ZN(n524) );
  AND2_X1 U564 ( .A1(n762), .A2(n986), .ZN(n525) );
  INV_X1 U565 ( .A(KEYINPUT64), .ZN(n701) );
  BUF_X1 U566 ( .A(n703), .Z(n714) );
  NOR2_X1 U567 ( .A1(n708), .A2(n707), .ZN(n709) );
  INV_X1 U568 ( .A(KEYINPUT29), .ZN(n723) );
  OR2_X1 U569 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U570 ( .A(n737), .B(KEYINPUT31), .ZN(n738) );
  INV_X1 U571 ( .A(KEYINPUT101), .ZN(n742) );
  INV_X1 U572 ( .A(n984), .ZN(n760) );
  AND2_X1 U573 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U574 ( .A1(n691), .A2(n690), .ZN(n695) );
  NOR2_X1 U575 ( .A1(n695), .A2(n786), .ZN(n703) );
  INV_X1 U576 ( .A(n703), .ZN(n729) );
  NAND2_X1 U577 ( .A1(n729), .A2(G8), .ZN(n781) );
  INV_X1 U578 ( .A(KEYINPUT105), .ZN(n769) );
  AND2_X1 U579 ( .A1(G40), .A2(n692), .ZN(n694) );
  AND2_X1 U580 ( .A1(G2105), .A2(n522), .ZN(n552) );
  XOR2_X1 U581 ( .A(KEYINPUT65), .B(n526), .Z(n641) );
  NOR2_X1 U582 ( .A1(n522), .A2(G2105), .ZN(n612) );
  XOR2_X1 U583 ( .A(KEYINPUT1), .B(n533), .Z(n653) );
  NOR2_X1 U584 ( .A1(n577), .A2(n576), .ZN(n579) );
  BUF_X1 U585 ( .A(n612), .Z(n889) );
  NOR2_X1 U586 ( .A1(G651), .A2(n655), .ZN(n649) );
  NAND2_X1 U587 ( .A1(n579), .A2(n578), .ZN(n688) );
  AND2_X1 U588 ( .A1(n555), .A2(n554), .ZN(n692) );
  NOR2_X1 U589 ( .A1(G651), .A2(G543), .ZN(n526) );
  NAND2_X1 U590 ( .A1(n641), .A2(G89), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n527), .B(KEYINPUT4), .ZN(n530) );
  XNOR2_X1 U592 ( .A(G543), .B(KEYINPUT0), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n528), .B(KEYINPUT67), .ZN(n655) );
  INV_X1 U594 ( .A(G651), .ZN(n532) );
  NOR2_X1 U595 ( .A1(n655), .A2(n532), .ZN(n642) );
  NAND2_X1 U596 ( .A1(G76), .A2(n642), .ZN(n529) );
  NAND2_X1 U597 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n531), .B(KEYINPUT5), .ZN(n538) );
  NOR2_X1 U599 ( .A1(G543), .A2(n532), .ZN(n533) );
  NAND2_X1 U600 ( .A1(G63), .A2(n653), .ZN(n535) );
  NAND2_X1 U601 ( .A1(G51), .A2(n649), .ZN(n534) );
  NAND2_X1 U602 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U603 ( .A(KEYINPUT6), .B(n536), .Z(n537) );
  NAND2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n539), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U606 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U607 ( .A1(G102), .A2(n612), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n540), .B(KEYINPUT88), .ZN(n547) );
  NAND2_X1 U609 ( .A1(n552), .A2(G126), .ZN(n542) );
  AND2_X1 U610 ( .A1(G2105), .A2(G2104), .ZN(n893) );
  NAND2_X1 U611 ( .A1(G114), .A2(n893), .ZN(n541) );
  AND2_X1 U612 ( .A1(n542), .A2(n541), .ZN(n545) );
  NOR2_X1 U613 ( .A1(G2105), .A2(G2104), .ZN(n543) );
  XOR2_X1 U614 ( .A(KEYINPUT17), .B(n543), .Z(n606) );
  NAND2_X1 U615 ( .A1(n606), .A2(G138), .ZN(n544) );
  AND2_X1 U616 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U617 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U618 ( .A(n548), .B(KEYINPUT89), .ZN(n689) );
  BUF_X1 U619 ( .A(n689), .Z(G164) );
  NAND2_X1 U620 ( .A1(n893), .A2(G113), .ZN(n551) );
  NAND2_X1 U621 ( .A1(G101), .A2(n612), .ZN(n549) );
  XOR2_X1 U622 ( .A(KEYINPUT23), .B(n549), .Z(n550) );
  AND2_X1 U623 ( .A1(n551), .A2(n550), .ZN(n693) );
  NAND2_X1 U624 ( .A1(G137), .A2(n606), .ZN(n555) );
  INV_X1 U625 ( .A(n552), .ZN(n553) );
  NAND2_X1 U626 ( .A1(G125), .A2(n894), .ZN(n554) );
  AND2_X1 U627 ( .A1(n693), .A2(n692), .ZN(G160) );
  XNOR2_X1 U628 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n560) );
  NAND2_X1 U629 ( .A1(G90), .A2(n641), .ZN(n557) );
  NAND2_X1 U630 ( .A1(G77), .A2(n642), .ZN(n556) );
  NAND2_X1 U631 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U632 ( .A(n558), .B(KEYINPUT9), .ZN(n559) );
  XNOR2_X1 U633 ( .A(n560), .B(n559), .ZN(n566) );
  NAND2_X1 U634 ( .A1(n653), .A2(G64), .ZN(n561) );
  XNOR2_X1 U635 ( .A(n561), .B(KEYINPUT68), .ZN(n563) );
  NAND2_X1 U636 ( .A1(G52), .A2(n649), .ZN(n562) );
  NAND2_X1 U637 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U638 ( .A(KEYINPUT69), .B(n564), .Z(n565) );
  NOR2_X1 U639 ( .A1(n566), .A2(n565), .ZN(G171) );
  INV_X1 U640 ( .A(G132), .ZN(G219) );
  INV_X1 U641 ( .A(G82), .ZN(G220) );
  INV_X1 U642 ( .A(G120), .ZN(G236) );
  INV_X1 U643 ( .A(G69), .ZN(G235) );
  INV_X1 U644 ( .A(G108), .ZN(G238) );
  NAND2_X1 U645 ( .A1(G94), .A2(G452), .ZN(n567) );
  XOR2_X1 U646 ( .A(KEYINPUT72), .B(n567), .Z(G173) );
  NAND2_X1 U647 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U648 ( .A(n568), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U649 ( .A(G223), .ZN(n844) );
  NAND2_X1 U650 ( .A1(n844), .A2(G567), .ZN(n569) );
  XOR2_X1 U651 ( .A(KEYINPUT11), .B(n569), .Z(G234) );
  XNOR2_X1 U652 ( .A(KEYINPUT73), .B(KEYINPUT13), .ZN(n574) );
  NAND2_X1 U653 ( .A1(n641), .A2(G81), .ZN(n570) );
  XNOR2_X1 U654 ( .A(n570), .B(KEYINPUT12), .ZN(n572) );
  NAND2_X1 U655 ( .A1(G68), .A2(n642), .ZN(n571) );
  NAND2_X1 U656 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U657 ( .A(n574), .B(n573), .ZN(n577) );
  NAND2_X1 U658 ( .A1(n653), .A2(G56), .ZN(n575) );
  XOR2_X1 U659 ( .A(KEYINPUT14), .B(n575), .Z(n576) );
  NAND2_X1 U660 ( .A1(n649), .A2(G43), .ZN(n578) );
  INV_X1 U661 ( .A(G860), .ZN(n599) );
  OR2_X1 U662 ( .A1(n688), .A2(n599), .ZN(G153) );
  INV_X1 U663 ( .A(G171), .ZN(G301) );
  NAND2_X1 U664 ( .A1(G66), .A2(n653), .ZN(n581) );
  NAND2_X1 U665 ( .A1(G54), .A2(n649), .ZN(n580) );
  NAND2_X1 U666 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U667 ( .A1(G92), .A2(n641), .ZN(n583) );
  NAND2_X1 U668 ( .A1(G79), .A2(n642), .ZN(n582) );
  NAND2_X1 U669 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U670 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U671 ( .A(n586), .B(KEYINPUT15), .ZN(n988) );
  INV_X1 U672 ( .A(G868), .ZN(n670) );
  NAND2_X1 U673 ( .A1(n988), .A2(n670), .ZN(n587) );
  XNOR2_X1 U674 ( .A(n587), .B(KEYINPUT74), .ZN(n589) );
  NAND2_X1 U675 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U676 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U677 ( .A1(G65), .A2(n653), .ZN(n591) );
  NAND2_X1 U678 ( .A1(G53), .A2(n649), .ZN(n590) );
  NAND2_X1 U679 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U680 ( .A1(G91), .A2(n641), .ZN(n593) );
  NAND2_X1 U681 ( .A1(G78), .A2(n642), .ZN(n592) );
  NAND2_X1 U682 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U683 ( .A1(n595), .A2(n594), .ZN(n976) );
  INV_X1 U684 ( .A(n976), .ZN(G299) );
  XNOR2_X1 U685 ( .A(KEYINPUT75), .B(G868), .ZN(n596) );
  NOR2_X1 U686 ( .A1(G286), .A2(n596), .ZN(n598) );
  NOR2_X1 U687 ( .A1(G868), .A2(G299), .ZN(n597) );
  NOR2_X1 U688 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U689 ( .A1(n599), .A2(G559), .ZN(n600) );
  INV_X1 U690 ( .A(n988), .ZN(n913) );
  NAND2_X1 U691 ( .A1(n600), .A2(n913), .ZN(n601) );
  XNOR2_X1 U692 ( .A(n601), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U693 ( .A1(n988), .A2(n670), .ZN(n602) );
  XOR2_X1 U694 ( .A(KEYINPUT76), .B(n602), .Z(n603) );
  NOR2_X1 U695 ( .A1(G559), .A2(n603), .ZN(n605) );
  NOR2_X1 U696 ( .A1(G868), .A2(n688), .ZN(n604) );
  NOR2_X1 U697 ( .A1(n605), .A2(n604), .ZN(G282) );
  NAND2_X1 U698 ( .A1(G111), .A2(n893), .ZN(n608) );
  BUF_X1 U699 ( .A(n606), .Z(n890) );
  NAND2_X1 U700 ( .A1(G135), .A2(n890), .ZN(n607) );
  NAND2_X1 U701 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U702 ( .A1(n894), .A2(G123), .ZN(n609) );
  XOR2_X1 U703 ( .A(KEYINPUT18), .B(n609), .Z(n610) );
  NOR2_X1 U704 ( .A1(n611), .A2(n610), .ZN(n614) );
  NAND2_X1 U705 ( .A1(n889), .A2(G99), .ZN(n613) );
  NAND2_X1 U706 ( .A1(n614), .A2(n613), .ZN(n925) );
  XOR2_X1 U707 ( .A(n925), .B(G2096), .Z(n616) );
  XNOR2_X1 U708 ( .A(G2100), .B(KEYINPUT77), .ZN(n615) );
  NAND2_X1 U709 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U710 ( .A(KEYINPUT78), .B(n617), .ZN(G156) );
  NAND2_X1 U711 ( .A1(G93), .A2(n641), .ZN(n619) );
  NAND2_X1 U712 ( .A1(G80), .A2(n642), .ZN(n618) );
  NAND2_X1 U713 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U714 ( .A1(G67), .A2(n653), .ZN(n620) );
  XNOR2_X1 U715 ( .A(KEYINPUT79), .B(n620), .ZN(n621) );
  NOR2_X1 U716 ( .A1(n622), .A2(n621), .ZN(n624) );
  NAND2_X1 U717 ( .A1(n649), .A2(G55), .ZN(n623) );
  NAND2_X1 U718 ( .A1(n624), .A2(n623), .ZN(n669) );
  NAND2_X1 U719 ( .A1(n913), .A2(G559), .ZN(n667) );
  XNOR2_X1 U720 ( .A(n688), .B(n667), .ZN(n625) );
  NOR2_X1 U721 ( .A1(G860), .A2(n625), .ZN(n626) );
  XOR2_X1 U722 ( .A(n669), .B(n626), .Z(G145) );
  NAND2_X1 U723 ( .A1(G88), .A2(n641), .ZN(n628) );
  NAND2_X1 U724 ( .A1(G62), .A2(n653), .ZN(n627) );
  NAND2_X1 U725 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U726 ( .A1(n642), .A2(G75), .ZN(n629) );
  XOR2_X1 U727 ( .A(KEYINPUT82), .B(n629), .Z(n630) );
  NOR2_X1 U728 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U729 ( .A1(n649), .A2(G50), .ZN(n632) );
  NAND2_X1 U730 ( .A1(n633), .A2(n632), .ZN(G303) );
  INV_X1 U731 ( .A(G303), .ZN(G166) );
  NAND2_X1 U732 ( .A1(G86), .A2(n641), .ZN(n635) );
  NAND2_X1 U733 ( .A1(G61), .A2(n653), .ZN(n634) );
  NAND2_X1 U734 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U735 ( .A1(n642), .A2(G73), .ZN(n636) );
  XOR2_X1 U736 ( .A(KEYINPUT2), .B(n636), .Z(n637) );
  NOR2_X1 U737 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U738 ( .A1(n649), .A2(G48), .ZN(n639) );
  NAND2_X1 U739 ( .A1(n640), .A2(n639), .ZN(G305) );
  AND2_X1 U740 ( .A1(n653), .A2(G60), .ZN(n646) );
  NAND2_X1 U741 ( .A1(G85), .A2(n641), .ZN(n644) );
  NAND2_X1 U742 ( .A1(G72), .A2(n642), .ZN(n643) );
  NAND2_X1 U743 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U744 ( .A1(n646), .A2(n645), .ZN(n648) );
  NAND2_X1 U745 ( .A1(n649), .A2(G47), .ZN(n647) );
  NAND2_X1 U746 ( .A1(n648), .A2(n647), .ZN(G290) );
  NAND2_X1 U747 ( .A1(G49), .A2(n649), .ZN(n651) );
  NAND2_X1 U748 ( .A1(G74), .A2(G651), .ZN(n650) );
  NAND2_X1 U749 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U750 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U751 ( .A(n654), .B(KEYINPUT80), .ZN(n657) );
  NAND2_X1 U752 ( .A1(G87), .A2(n655), .ZN(n656) );
  NAND2_X1 U753 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U754 ( .A(KEYINPUT81), .B(n658), .Z(G288) );
  XNOR2_X1 U755 ( .A(G166), .B(G305), .ZN(n664) );
  XOR2_X1 U756 ( .A(KEYINPUT84), .B(KEYINPUT19), .Z(n660) );
  XNOR2_X1 U757 ( .A(n976), .B(KEYINPUT83), .ZN(n659) );
  XNOR2_X1 U758 ( .A(n660), .B(n659), .ZN(n661) );
  XOR2_X1 U759 ( .A(n661), .B(G290), .Z(n662) );
  XNOR2_X1 U760 ( .A(n669), .B(n662), .ZN(n663) );
  XNOR2_X1 U761 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U762 ( .A(n665), .B(G288), .ZN(n666) );
  XNOR2_X1 U763 ( .A(n666), .B(n688), .ZN(n912) );
  XNOR2_X1 U764 ( .A(n667), .B(n912), .ZN(n668) );
  NAND2_X1 U765 ( .A1(n668), .A2(G868), .ZN(n672) );
  NAND2_X1 U766 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U767 ( .A1(n672), .A2(n671), .ZN(G295) );
  NAND2_X1 U768 ( .A1(G2084), .A2(G2078), .ZN(n673) );
  XNOR2_X1 U769 ( .A(n673), .B(KEYINPUT20), .ZN(n674) );
  XNOR2_X1 U770 ( .A(n674), .B(KEYINPUT85), .ZN(n675) );
  NAND2_X1 U771 ( .A1(n675), .A2(G2090), .ZN(n676) );
  XNOR2_X1 U772 ( .A(KEYINPUT21), .B(n676), .ZN(n677) );
  NAND2_X1 U773 ( .A1(n677), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U774 ( .A(KEYINPUT86), .B(G44), .ZN(n678) );
  XNOR2_X1 U775 ( .A(n678), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U776 ( .A1(G235), .A2(G236), .ZN(n679) );
  XNOR2_X1 U777 ( .A(n679), .B(KEYINPUT87), .ZN(n680) );
  NOR2_X1 U778 ( .A1(G238), .A2(n680), .ZN(n681) );
  NAND2_X1 U779 ( .A1(G57), .A2(n681), .ZN(n850) );
  NAND2_X1 U780 ( .A1(n850), .A2(G567), .ZN(n686) );
  NOR2_X1 U781 ( .A1(G220), .A2(G219), .ZN(n682) );
  XOR2_X1 U782 ( .A(KEYINPUT22), .B(n682), .Z(n683) );
  NOR2_X1 U783 ( .A1(G218), .A2(n683), .ZN(n684) );
  NAND2_X1 U784 ( .A1(G96), .A2(n684), .ZN(n851) );
  NAND2_X1 U785 ( .A1(n851), .A2(G2106), .ZN(n685) );
  NAND2_X1 U786 ( .A1(n686), .A2(n685), .ZN(n852) );
  NAND2_X1 U787 ( .A1(G483), .A2(G661), .ZN(n687) );
  NOR2_X1 U788 ( .A1(n852), .A2(n687), .ZN(n849) );
  NAND2_X1 U789 ( .A1(n849), .A2(G36), .ZN(G176) );
  INV_X1 U790 ( .A(n688), .ZN(n700) );
  INV_X1 U791 ( .A(n689), .ZN(n691) );
  INV_X1 U792 ( .A(G1384), .ZN(n690) );
  NAND2_X1 U793 ( .A1(n694), .A2(n693), .ZN(n786) );
  NAND2_X1 U794 ( .A1(n703), .A2(G1996), .ZN(n697) );
  INV_X1 U795 ( .A(KEYINPUT26), .ZN(n696) );
  XNOR2_X1 U796 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X1 U797 ( .A1(n698), .A2(n521), .ZN(n699) );
  XNOR2_X1 U798 ( .A(n702), .B(n701), .ZN(n710) );
  NOR2_X1 U799 ( .A1(n710), .A2(n988), .ZN(n708) );
  NAND2_X1 U800 ( .A1(G1348), .A2(n729), .ZN(n705) );
  NAND2_X1 U801 ( .A1(G2067), .A2(n714), .ZN(n704) );
  NAND2_X1 U802 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U803 ( .A(KEYINPUT98), .B(n706), .Z(n707) );
  XNOR2_X1 U804 ( .A(n709), .B(KEYINPUT99), .ZN(n712) );
  NAND2_X1 U805 ( .A1(n710), .A2(n988), .ZN(n711) );
  NAND2_X1 U806 ( .A1(n712), .A2(n711), .ZN(n718) );
  NAND2_X1 U807 ( .A1(n714), .A2(G2072), .ZN(n713) );
  XNOR2_X1 U808 ( .A(n713), .B(KEYINPUT27), .ZN(n716) );
  INV_X1 U809 ( .A(G1956), .ZN(n1006) );
  NOR2_X1 U810 ( .A1(n1006), .A2(n714), .ZN(n715) );
  NOR2_X1 U811 ( .A1(n716), .A2(n715), .ZN(n719) );
  NAND2_X1 U812 ( .A1(n976), .A2(n719), .ZN(n717) );
  NAND2_X1 U813 ( .A1(n718), .A2(n717), .ZN(n722) );
  NOR2_X1 U814 ( .A1(n976), .A2(n719), .ZN(n720) );
  XOR2_X1 U815 ( .A(n720), .B(KEYINPUT28), .Z(n721) );
  NAND2_X1 U816 ( .A1(n722), .A2(n721), .ZN(n724) );
  XNOR2_X1 U817 ( .A(KEYINPUT25), .B(G2078), .ZN(n961) );
  NOR2_X1 U818 ( .A1(n729), .A2(n961), .ZN(n726) );
  AND2_X1 U819 ( .A1(n729), .A2(G1961), .ZN(n725) );
  NOR2_X1 U820 ( .A1(n726), .A2(n725), .ZN(n734) );
  NAND2_X1 U821 ( .A1(G171), .A2(n734), .ZN(n727) );
  NAND2_X1 U822 ( .A1(n728), .A2(n727), .ZN(n739) );
  NOR2_X1 U823 ( .A1(G2084), .A2(n729), .ZN(n744) );
  NOR2_X1 U824 ( .A1(G1966), .A2(n781), .ZN(n740) );
  NOR2_X1 U825 ( .A1(n744), .A2(n740), .ZN(n730) );
  XNOR2_X1 U826 ( .A(KEYINPUT100), .B(n730), .ZN(n731) );
  NAND2_X1 U827 ( .A1(n731), .A2(G8), .ZN(n732) );
  XNOR2_X1 U828 ( .A(KEYINPUT30), .B(n732), .ZN(n733) );
  NOR2_X1 U829 ( .A1(G168), .A2(n733), .ZN(n736) );
  NOR2_X1 U830 ( .A1(G171), .A2(n734), .ZN(n735) );
  NAND2_X1 U831 ( .A1(n739), .A2(n738), .ZN(n750) );
  INV_X1 U832 ( .A(n740), .ZN(n741) );
  XNOR2_X1 U833 ( .A(n743), .B(n742), .ZN(n746) );
  NAND2_X1 U834 ( .A1(G8), .A2(n744), .ZN(n745) );
  NAND2_X1 U835 ( .A1(n746), .A2(n745), .ZN(n756) );
  NOR2_X1 U836 ( .A1(G1971), .A2(n781), .ZN(n748) );
  NOR2_X1 U837 ( .A1(G2090), .A2(n729), .ZN(n747) );
  NOR2_X1 U838 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U839 ( .A1(n749), .A2(G303), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n750), .A2(G286), .ZN(n751) );
  NAND2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U842 ( .A1(G8), .A2(n753), .ZN(n754) );
  XNOR2_X1 U843 ( .A(KEYINPUT32), .B(n754), .ZN(n755) );
  NAND2_X1 U844 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U845 ( .A(n757), .B(KEYINPUT102), .ZN(n779) );
  NOR2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n758) );
  XOR2_X1 U847 ( .A(KEYINPUT103), .B(n758), .Z(n984) );
  NOR2_X1 U848 ( .A1(G1971), .A2(G303), .ZN(n978) );
  XOR2_X1 U849 ( .A(n978), .B(KEYINPUT104), .Z(n759) );
  NAND2_X1 U850 ( .A1(n779), .A2(n761), .ZN(n762) );
  NAND2_X1 U851 ( .A1(G1976), .A2(G288), .ZN(n986) );
  INV_X1 U852 ( .A(n781), .ZN(n765) );
  NAND2_X1 U853 ( .A1(n525), .A2(n764), .ZN(n768) );
  NAND2_X1 U854 ( .A1(n984), .A2(n765), .ZN(n766) );
  NAND2_X1 U855 ( .A1(n766), .A2(KEYINPUT33), .ZN(n767) );
  NAND2_X1 U856 ( .A1(n768), .A2(n767), .ZN(n770) );
  XNOR2_X1 U857 ( .A(n770), .B(n769), .ZN(n772) );
  XNOR2_X1 U858 ( .A(G1981), .B(G305), .ZN(n995) );
  NAND2_X1 U859 ( .A1(n772), .A2(n771), .ZN(n785) );
  NOR2_X1 U860 ( .A1(G1981), .A2(G305), .ZN(n773) );
  XOR2_X1 U861 ( .A(n773), .B(KEYINPUT96), .Z(n774) );
  XNOR2_X1 U862 ( .A(KEYINPUT24), .B(n774), .ZN(n775) );
  NOR2_X1 U863 ( .A1(n781), .A2(n775), .ZN(n776) );
  XNOR2_X1 U864 ( .A(n776), .B(KEYINPUT97), .ZN(n784) );
  NOR2_X1 U865 ( .A1(G2090), .A2(G303), .ZN(n777) );
  NAND2_X1 U866 ( .A1(G8), .A2(n777), .ZN(n778) );
  XNOR2_X1 U867 ( .A(n778), .B(KEYINPUT106), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n782) );
  NAND2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n785), .A2(n524), .ZN(n819) );
  XNOR2_X1 U871 ( .A(G1986), .B(G290), .ZN(n980) );
  NOR2_X1 U872 ( .A1(G164), .A2(G1384), .ZN(n787) );
  NOR2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n830) );
  NAND2_X1 U874 ( .A1(n980), .A2(n830), .ZN(n788) );
  XNOR2_X1 U875 ( .A(n788), .B(KEYINPUT90), .ZN(n808) );
  NAND2_X1 U876 ( .A1(G107), .A2(n893), .ZN(n790) );
  NAND2_X1 U877 ( .A1(G131), .A2(n890), .ZN(n789) );
  NAND2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n794) );
  NAND2_X1 U879 ( .A1(G95), .A2(n889), .ZN(n792) );
  NAND2_X1 U880 ( .A1(G119), .A2(n894), .ZN(n791) );
  NAND2_X1 U881 ( .A1(n792), .A2(n791), .ZN(n793) );
  OR2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n900) );
  NAND2_X1 U883 ( .A1(G1991), .A2(n900), .ZN(n795) );
  XNOR2_X1 U884 ( .A(n795), .B(KEYINPUT92), .ZN(n807) );
  NAND2_X1 U885 ( .A1(G117), .A2(n893), .ZN(n797) );
  NAND2_X1 U886 ( .A1(G129), .A2(n894), .ZN(n796) );
  NAND2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U888 ( .A(KEYINPUT93), .B(n798), .Z(n801) );
  NAND2_X1 U889 ( .A1(n889), .A2(G105), .ZN(n799) );
  XOR2_X1 U890 ( .A(KEYINPUT38), .B(n799), .Z(n800) );
  NOR2_X1 U891 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U892 ( .A(KEYINPUT94), .B(n802), .ZN(n805) );
  NAND2_X1 U893 ( .A1(n890), .A2(G141), .ZN(n803) );
  XOR2_X1 U894 ( .A(KEYINPUT95), .B(n803), .Z(n804) );
  NAND2_X1 U895 ( .A1(n805), .A2(n804), .ZN(n905) );
  NAND2_X1 U896 ( .A1(G1996), .A2(n905), .ZN(n806) );
  NAND2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n938) );
  NAND2_X1 U898 ( .A1(n830), .A2(n938), .ZN(n822) );
  XOR2_X1 U899 ( .A(G2067), .B(KEYINPUT37), .Z(n809) );
  XNOR2_X1 U900 ( .A(KEYINPUT91), .B(n809), .ZN(n828) );
  NAND2_X1 U901 ( .A1(G104), .A2(n889), .ZN(n811) );
  NAND2_X1 U902 ( .A1(G140), .A2(n890), .ZN(n810) );
  NAND2_X1 U903 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U904 ( .A(KEYINPUT34), .B(n812), .ZN(n817) );
  NAND2_X1 U905 ( .A1(G116), .A2(n893), .ZN(n814) );
  NAND2_X1 U906 ( .A1(G128), .A2(n894), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n815) );
  XOR2_X1 U908 ( .A(KEYINPUT35), .B(n815), .Z(n816) );
  NOR2_X1 U909 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U910 ( .A(KEYINPUT36), .B(n818), .ZN(n906) );
  NOR2_X1 U911 ( .A1(n828), .A2(n906), .ZN(n934) );
  NAND2_X1 U912 ( .A1(n830), .A2(n934), .ZN(n827) );
  NAND2_X1 U913 ( .A1(n819), .A2(n520), .ZN(n833) );
  NOR2_X1 U914 ( .A1(G1986), .A2(G290), .ZN(n820) );
  NOR2_X1 U915 ( .A1(G1991), .A2(n900), .ZN(n928) );
  NOR2_X1 U916 ( .A1(n820), .A2(n928), .ZN(n821) );
  XNOR2_X1 U917 ( .A(n821), .B(KEYINPUT107), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n823), .A2(n822), .ZN(n824) );
  OR2_X1 U919 ( .A1(n905), .A2(G1996), .ZN(n929) );
  NAND2_X1 U920 ( .A1(n824), .A2(n929), .ZN(n825) );
  XOR2_X1 U921 ( .A(KEYINPUT39), .B(n825), .Z(n826) );
  NAND2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n828), .A2(n906), .ZN(n949) );
  NAND2_X1 U924 ( .A1(n829), .A2(n949), .ZN(n831) );
  NAND2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U927 ( .A(n834), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U928 ( .A(G1348), .B(G2454), .ZN(n835) );
  XNOR2_X1 U929 ( .A(n835), .B(G2430), .ZN(n836) );
  XNOR2_X1 U930 ( .A(n836), .B(G1341), .ZN(n842) );
  XOR2_X1 U931 ( .A(G2443), .B(G2427), .Z(n838) );
  XNOR2_X1 U932 ( .A(G2438), .B(G2446), .ZN(n837) );
  XNOR2_X1 U933 ( .A(n838), .B(n837), .ZN(n840) );
  XOR2_X1 U934 ( .A(G2451), .B(G2435), .Z(n839) );
  XNOR2_X1 U935 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U936 ( .A(n842), .B(n841), .ZN(n843) );
  NAND2_X1 U937 ( .A1(n843), .A2(G14), .ZN(n918) );
  XOR2_X1 U938 ( .A(KEYINPUT108), .B(n918), .Z(G401) );
  NAND2_X1 U939 ( .A1(G2106), .A2(n844), .ZN(G217) );
  NAND2_X1 U940 ( .A1(G15), .A2(G2), .ZN(n846) );
  INV_X1 U941 ( .A(G661), .ZN(n845) );
  NOR2_X1 U942 ( .A1(n846), .A2(n845), .ZN(n847) );
  XNOR2_X1 U943 ( .A(n847), .B(KEYINPUT109), .ZN(G259) );
  NAND2_X1 U944 ( .A1(G3), .A2(G1), .ZN(n848) );
  NAND2_X1 U945 ( .A1(n849), .A2(n848), .ZN(G188) );
  INV_X1 U947 ( .A(G96), .ZN(G221) );
  NOR2_X1 U948 ( .A1(n851), .A2(n850), .ZN(G325) );
  INV_X1 U949 ( .A(G325), .ZN(G261) );
  INV_X1 U950 ( .A(n852), .ZN(G319) );
  XOR2_X1 U951 ( .A(KEYINPUT111), .B(KEYINPUT110), .Z(n854) );
  XNOR2_X1 U952 ( .A(G2678), .B(KEYINPUT43), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U954 ( .A(KEYINPUT42), .B(G2090), .Z(n856) );
  XNOR2_X1 U955 ( .A(G2067), .B(G2072), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U957 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U958 ( .A(G2096), .B(G2100), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n862) );
  XOR2_X1 U960 ( .A(G2084), .B(G2078), .Z(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(G227) );
  XOR2_X1 U962 ( .A(G1971), .B(G1956), .Z(n864) );
  XNOR2_X1 U963 ( .A(G1986), .B(G1976), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U965 ( .A(n865), .B(KEYINPUT41), .Z(n867) );
  XNOR2_X1 U966 ( .A(G1996), .B(G1991), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n867), .B(n866), .ZN(n871) );
  XOR2_X1 U968 ( .A(G2474), .B(G1961), .Z(n869) );
  XNOR2_X1 U969 ( .A(G1981), .B(G1966), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(G229) );
  NAND2_X1 U972 ( .A1(n889), .A2(G100), .ZN(n878) );
  NAND2_X1 U973 ( .A1(G112), .A2(n893), .ZN(n873) );
  NAND2_X1 U974 ( .A1(G136), .A2(n890), .ZN(n872) );
  NAND2_X1 U975 ( .A1(n873), .A2(n872), .ZN(n876) );
  NAND2_X1 U976 ( .A1(n894), .A2(G124), .ZN(n874) );
  XOR2_X1 U977 ( .A(KEYINPUT44), .B(n874), .Z(n875) );
  NOR2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n877) );
  NAND2_X1 U979 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U980 ( .A(KEYINPUT112), .B(n879), .Z(G162) );
  NAND2_X1 U981 ( .A1(G118), .A2(n893), .ZN(n881) );
  NAND2_X1 U982 ( .A1(G130), .A2(n894), .ZN(n880) );
  NAND2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n886) );
  NAND2_X1 U984 ( .A1(G106), .A2(n889), .ZN(n883) );
  NAND2_X1 U985 ( .A1(G142), .A2(n890), .ZN(n882) );
  NAND2_X1 U986 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U987 ( .A(n884), .B(KEYINPUT45), .Z(n885) );
  NOR2_X1 U988 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U989 ( .A(n887), .B(G162), .ZN(n910) );
  XOR2_X1 U990 ( .A(G164), .B(G160), .Z(n888) );
  XNOR2_X1 U991 ( .A(n925), .B(n888), .ZN(n904) );
  XNOR2_X1 U992 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n902) );
  NAND2_X1 U993 ( .A1(G103), .A2(n889), .ZN(n892) );
  NAND2_X1 U994 ( .A1(G139), .A2(n890), .ZN(n891) );
  NAND2_X1 U995 ( .A1(n892), .A2(n891), .ZN(n899) );
  NAND2_X1 U996 ( .A1(G115), .A2(n893), .ZN(n896) );
  NAND2_X1 U997 ( .A1(G127), .A2(n894), .ZN(n895) );
  NAND2_X1 U998 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U999 ( .A(KEYINPUT47), .B(n897), .Z(n898) );
  NOR2_X1 U1000 ( .A1(n899), .A2(n898), .ZN(n940) );
  XNOR2_X1 U1001 ( .A(n900), .B(n940), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n908) );
  XOR2_X1 U1004 ( .A(n906), .B(n905), .Z(n907) );
  XNOR2_X1 U1005 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1006 ( .A(n910), .B(n909), .Z(n911) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n911), .ZN(G395) );
  XOR2_X1 U1008 ( .A(KEYINPUT113), .B(n912), .Z(n915) );
  XNOR2_X1 U1009 ( .A(n913), .B(G286), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(n915), .B(n914), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(n916), .B(G301), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n917), .ZN(G397) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n918), .ZN(n921) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(n919), .B(KEYINPUT49), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1017 ( .A(KEYINPUT114), .B(n922), .ZN(n924) );
  NOR2_X1 U1018 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1019 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  INV_X1 U1021 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1022 ( .A(G160), .B(G2084), .ZN(n926) );
  NAND2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n936) );
  XNOR2_X1 U1025 ( .A(G162), .B(G2090), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(n931), .B(KEYINPUT115), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(KEYINPUT51), .B(n932), .ZN(n933) );
  NOR2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1031 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1032 ( .A(KEYINPUT116), .B(n939), .Z(n947) );
  XOR2_X1 U1033 ( .A(G2072), .B(n940), .Z(n942) );
  XOR2_X1 U1034 ( .A(G164), .B(G2078), .Z(n941) );
  NOR2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n945) );
  XNOR2_X1 U1036 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(n943), .B(KEYINPUT50), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(n945), .B(n944), .ZN(n946) );
  NOR2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1040 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1041 ( .A(n950), .B(KEYINPUT52), .ZN(n951) );
  XNOR2_X1 U1042 ( .A(KEYINPUT119), .B(n951), .ZN(n952) );
  INV_X1 U1043 ( .A(KEYINPUT55), .ZN(n971) );
  NAND2_X1 U1044 ( .A1(n952), .A2(n971), .ZN(n953) );
  NAND2_X1 U1045 ( .A1(n953), .A2(G29), .ZN(n1036) );
  XNOR2_X1 U1046 ( .A(G2090), .B(G35), .ZN(n966) );
  XNOR2_X1 U1047 ( .A(G1996), .B(G32), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(G33), .B(G2072), .ZN(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n960) );
  XOR2_X1 U1050 ( .A(G1991), .B(G25), .Z(n956) );
  NAND2_X1 U1051 ( .A1(n956), .A2(G28), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(G26), .B(G2067), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n963) );
  XOR2_X1 U1055 ( .A(G27), .B(n961), .Z(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(KEYINPUT53), .B(n964), .ZN(n965) );
  NOR2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n969) );
  XOR2_X1 U1059 ( .A(G2084), .B(G34), .Z(n967) );
  XNOR2_X1 U1060 ( .A(KEYINPUT54), .B(n967), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(n971), .B(n970), .ZN(n973) );
  INV_X1 U1063 ( .A(G29), .ZN(n972) );
  NAND2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1065 ( .A1(G11), .A2(n974), .ZN(n1034) );
  INV_X1 U1066 ( .A(G16), .ZN(n1030) );
  XOR2_X1 U1067 ( .A(KEYINPUT56), .B(KEYINPUT120), .Z(n975) );
  XNOR2_X1 U1068 ( .A(n1030), .B(n975), .ZN(n1003) );
  XNOR2_X1 U1069 ( .A(G171), .B(G1961), .ZN(n1001) );
  XNOR2_X1 U1070 ( .A(n976), .B(n1006), .ZN(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n982) );
  AND2_X1 U1072 ( .A1(G303), .A2(G1971), .ZN(n979) );
  NOR2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1077 ( .A(n987), .B(KEYINPUT123), .ZN(n993) );
  XNOR2_X1 U1078 ( .A(G1348), .B(KEYINPUT122), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(n989), .B(n988), .ZN(n991) );
  XNOR2_X1 U1080 ( .A(G1341), .B(n688), .ZN(n990) );
  NOR2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n999) );
  XOR2_X1 U1083 ( .A(G1966), .B(G168), .Z(n994) );
  NOR2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1085 ( .A(KEYINPUT121), .B(n996), .Z(n997) );
  XNOR2_X1 U1086 ( .A(n997), .B(KEYINPUT57), .ZN(n998) );
  NOR2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1089 ( .A1(n1003), .A2(n1002), .ZN(n1032) );
  XOR2_X1 U1090 ( .A(KEYINPUT124), .B(G4), .Z(n1005) );
  XNOR2_X1 U1091 ( .A(G1348), .B(KEYINPUT59), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(n1005), .B(n1004), .ZN(n1012) );
  XNOR2_X1 U1093 ( .A(G20), .B(n1006), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(G1981), .B(G6), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(G1341), .B(G19), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1099 ( .A(KEYINPUT60), .B(n1013), .Z(n1014) );
  XNOR2_X1 U1100 ( .A(KEYINPUT125), .B(n1014), .ZN(n1018) );
  XNOR2_X1 U1101 ( .A(G1966), .B(G21), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(G1961), .B(G5), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(KEYINPUT126), .B(n1019), .ZN(n1027) );
  XOR2_X1 U1106 ( .A(G1986), .B(G24), .Z(n1023) );
  XNOR2_X1 U1107 ( .A(G1976), .B(G23), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(G1971), .B(G22), .ZN(n1020) );
  NOR2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1111 ( .A(KEYINPUT127), .B(n1024), .Z(n1025) );
  XNOR2_X1 U1112 ( .A(KEYINPUT58), .B(n1025), .ZN(n1026) );
  NOR2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1114 ( .A(KEYINPUT61), .B(n1028), .ZN(n1029) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1117 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1118 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XOR2_X1 U1119 ( .A(KEYINPUT62), .B(n1037), .Z(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

