//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n210), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(KEYINPUT64), .B(G68), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G58), .A2(G232), .ZN(new_n229));
  NAND4_X1  g0029(.A1(new_n226), .A2(new_n227), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n212), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n215), .B(new_n221), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT65), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n237), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n202), .A2(G68), .ZN(new_n246));
  INV_X1    g0046(.A(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n245), .B(new_n251), .Z(G351));
  NAND2_X1  g0052(.A1(G20), .A2(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT15), .B(G87), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n210), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT8), .B(G58), .ZN(new_n258));
  OAI221_X1 g0058(.A(new_n253), .B1(new_n254), .B2(new_n255), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n219), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G13), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G1), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G77), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n261), .B1(new_n209), .B2(G20), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n268), .B1(new_n270), .B2(new_n267), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n262), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(G232), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(G238), .A3(G1698), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT3), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G107), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n276), .A2(new_n277), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT71), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n276), .A2(new_n277), .A3(KEYINPUT71), .A4(new_n283), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G274), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n287), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(KEYINPUT67), .ZN(new_n294));
  INV_X1    g0094(.A(G41), .ZN(new_n295));
  OAI211_X1 g0095(.A(G1), .B(G13), .C1(new_n278), .C2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT67), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n297), .B(new_n209), .C1(G41), .C2(G45), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n294), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n299), .A2(KEYINPUT68), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT68), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n294), .A2(new_n301), .A3(new_n296), .A4(new_n298), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(G244), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n289), .A2(new_n293), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n273), .B1(new_n305), .B2(G200), .ZN(new_n306));
  INV_X1    g0106(.A(G190), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n306), .B1(new_n307), .B2(new_n305), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n305), .A2(G179), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n272), .B1(new_n305), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT72), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n309), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  AOI211_X1 g0113(.A(KEYINPUT72), .B(new_n272), .C1(new_n305), .C2(new_n310), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n308), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT73), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n274), .A2(G232), .A3(G1698), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n274), .A2(G226), .A3(new_n275), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G33), .A2(G97), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n292), .B1(new_n321), .B2(new_n287), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n299), .A2(KEYINPUT68), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n224), .B1(new_n324), .B2(new_n302), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT13), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(G238), .B1(new_n300), .B2(new_n303), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT13), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n322), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n326), .A2(G190), .A3(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n222), .A2(new_n210), .ZN(new_n331));
  OAI22_X1  g0131(.A1(new_n257), .A2(new_n202), .B1(new_n255), .B2(new_n267), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n261), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT76), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT76), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n335), .B(new_n261), .C1(new_n331), .C2(new_n332), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT11), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT11), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n334), .A2(new_n339), .A3(new_n336), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n331), .A2(KEYINPUT12), .A3(new_n264), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(KEYINPUT12), .B2(new_n266), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n247), .B1(new_n270), .B2(KEYINPUT12), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n338), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n330), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G200), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(new_n326), .B2(new_n329), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  AND3_X1   g0149(.A1(new_n327), .A2(new_n328), .A3(new_n322), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n328), .B1(new_n327), .B2(new_n322), .ZN(new_n351));
  OAI21_X1  g0151(.A(G169), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT14), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n326), .A2(G179), .A3(new_n329), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT14), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n355), .B(G169), .C1(new_n350), .C2(new_n351), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n353), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n345), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n349), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n308), .B(KEYINPUT73), .C1(new_n313), .C2(new_n314), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n317), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n261), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT16), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n201), .B1(new_n222), .B2(G58), .ZN(new_n364));
  INV_X1    g0164(.A(G159), .ZN(new_n365));
  OAI22_X1  g0165(.A1(new_n364), .A2(new_n210), .B1(new_n365), .B2(new_n257), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT7), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n274), .B2(G20), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n282), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n223), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n363), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT79), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n274), .A2(new_n367), .A3(G20), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT7), .B1(new_n282), .B2(new_n210), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n222), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AND2_X1   g0176(.A1(KEYINPUT64), .A2(G68), .ZN(new_n377));
  NOR2_X1   g0177(.A1(KEYINPUT64), .A2(G68), .ZN(new_n378));
  OAI21_X1  g0178(.A(G58), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n210), .B1(new_n379), .B2(new_n216), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n257), .A2(new_n365), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n383), .A2(KEYINPUT79), .A3(new_n363), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n362), .B1(new_n373), .B2(new_n384), .ZN(new_n385));
  NOR3_X1   g0185(.A1(new_n380), .A2(new_n363), .A3(new_n381), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n280), .A2(G33), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n278), .A2(KEYINPUT3), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT77), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT77), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n279), .A2(new_n281), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(new_n210), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n374), .B1(new_n392), .B2(new_n367), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n386), .B1(new_n393), .B2(new_n247), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT78), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(KEYINPUT78), .B(new_n386), .C1(new_n393), .C2(new_n247), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n385), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(KEYINPUT69), .A2(G58), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n400), .B(KEYINPUT8), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n266), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(new_n401), .B2(new_n270), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT80), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n294), .A2(new_n296), .A3(new_n298), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n292), .B1(new_n406), .B2(G232), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n279), .A2(new_n281), .A3(G226), .A4(G1698), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n279), .A2(new_n281), .A3(G223), .A4(new_n275), .ZN(new_n409));
  INV_X1    g0209(.A(G87), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n408), .B(new_n409), .C1(new_n278), .C2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n287), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n407), .A2(new_n307), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(G200), .B1(new_n407), .B2(new_n412), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n405), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n407), .A2(new_n412), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n347), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n407), .A2(new_n307), .A3(new_n412), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(KEYINPUT80), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  AND4_X1   g0220(.A1(KEYINPUT17), .A2(new_n399), .A3(new_n404), .A4(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n403), .B1(new_n385), .B2(new_n398), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT17), .B1(new_n422), .B2(new_n420), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n396), .A2(new_n397), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT79), .B1(new_n383), .B2(new_n363), .ZN(new_n426));
  AOI211_X1 g0226(.A(new_n372), .B(KEYINPUT16), .C1(new_n376), .C2(new_n382), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n261), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n404), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(G179), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n416), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(G169), .B2(new_n416), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n429), .A2(KEYINPUT18), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT18), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n422), .B2(new_n432), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n424), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n274), .A2(G222), .A3(new_n275), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n274), .A2(G1698), .ZN(new_n441));
  INV_X1    g0241(.A(G223), .ZN(new_n442));
  OAI221_X1 g0242(.A(new_n440), .B1(new_n267), .B2(new_n274), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n292), .B1(new_n443), .B2(new_n287), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT66), .B(G226), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n300), .B2(new_n303), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n255), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n401), .A2(new_n449), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n256), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n261), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n265), .A2(G50), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n454), .B1(G50), .B2(new_n269), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n448), .A2(new_n310), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n444), .A2(new_n430), .A3(new_n447), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(KEYINPUT70), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT70), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n460), .B1(new_n456), .B2(new_n457), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n453), .A2(KEYINPUT9), .A3(new_n455), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT9), .B1(new_n453), .B2(new_n455), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT10), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n444), .A2(G190), .A3(new_n447), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT75), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT74), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n448), .A2(new_n471), .A3(G200), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n448), .A2(G200), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT74), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n469), .A2(new_n470), .A3(new_n472), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n472), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT75), .B1(new_n476), .B2(new_n468), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n473), .A2(new_n465), .A3(new_n467), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT10), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n462), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n361), .A2(new_n439), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n274), .A2(G257), .A3(new_n275), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n282), .A2(G303), .ZN(new_n484));
  INV_X1    g0284(.A(G264), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n483), .B(new_n484), .C1(new_n441), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n287), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT5), .B(G41), .ZN(new_n488));
  INV_X1    g0288(.A(G45), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(G1), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(G270), .A3(new_n296), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n488), .A2(new_n296), .A3(G274), .A4(new_n490), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n492), .A2(KEYINPUT86), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(KEYINPUT86), .B1(new_n492), .B2(new_n493), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n487), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(G20), .B1(G33), .B2(G283), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(G33), .B2(new_n205), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT87), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT87), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n497), .B(new_n500), .C1(G33), .C2(new_n205), .ZN(new_n501));
  INV_X1    g0301(.A(G116), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G20), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n499), .A2(new_n261), .A3(new_n501), .A4(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT20), .ZN(new_n505));
  OR2_X1    g0305(.A1(new_n505), .A2(KEYINPUT88), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(KEYINPUT88), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n265), .A2(G116), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n209), .A2(G33), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n362), .A2(new_n265), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n509), .B1(new_n512), .B2(G116), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n261), .A2(new_n503), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(KEYINPUT87), .B2(new_n498), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n515), .A2(KEYINPUT88), .A3(new_n505), .A4(new_n501), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n508), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n496), .A2(new_n517), .A3(KEYINPUT21), .A4(G169), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n492), .A2(new_n493), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT86), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n492), .A2(KEYINPUT86), .A3(new_n493), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n517), .A2(new_n523), .A3(G179), .A4(new_n487), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n517), .B1(new_n496), .B2(G200), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n307), .B2(new_n496), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n496), .A2(new_n517), .A3(G169), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT21), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n525), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n266), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(KEYINPUT25), .B1(new_n266), .B2(new_n206), .ZN(new_n534));
  OAI22_X1  g0334(.A1(new_n533), .A2(new_n534), .B1(new_n511), .B2(new_n206), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n491), .A2(G264), .A3(new_n296), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT90), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n287), .B1(new_n490), .B2(new_n488), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT90), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n539), .A2(new_n540), .A3(G264), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n274), .A2(G257), .A3(G1698), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n274), .A2(G250), .A3(new_n275), .ZN(new_n544));
  INV_X1    g0344(.A(G294), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n543), .B(new_n544), .C1(new_n278), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n287), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n542), .A2(new_n493), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n347), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n538), .A2(new_n541), .B1(new_n546), .B2(new_n287), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n550), .A2(new_n307), .A3(new_n493), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT89), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n274), .A2(new_n210), .A3(G87), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT22), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT22), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n274), .A2(new_n556), .A3(new_n210), .A4(G87), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT23), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n210), .B2(G107), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n278), .A2(new_n502), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n210), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n558), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT24), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT24), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n558), .A2(new_n569), .A3(new_n566), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n553), .B1(new_n571), .B2(new_n261), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n569), .B1(new_n558), .B2(new_n566), .ZN(new_n573));
  AOI211_X1 g0373(.A(KEYINPUT24), .B(new_n565), .C1(new_n555), .C2(new_n557), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n553), .B(new_n261), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n536), .B(new_n552), .C1(new_n572), .C2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n261), .B1(new_n573), .B2(new_n574), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT89), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n535), .B1(new_n579), .B2(new_n575), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n548), .A2(new_n310), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(G179), .B2(new_n548), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n577), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT6), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n584), .A2(new_n205), .A3(G107), .ZN(new_n585));
  XNOR2_X1  g0385(.A(G97), .B(G107), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n585), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  OAI22_X1  g0387(.A1(new_n587), .A2(new_n210), .B1(new_n267), .B2(new_n257), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n206), .B1(new_n368), .B2(new_n369), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n261), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n265), .A2(G97), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n512), .B2(G97), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT81), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n590), .A2(KEYINPUT81), .A3(new_n592), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n539), .A2(G257), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n493), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n282), .A2(new_n275), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n599), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n279), .A2(new_n281), .A3(G244), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n601), .A2(KEYINPUT82), .A3(KEYINPUT4), .A4(new_n275), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n274), .A2(KEYINPUT4), .A3(G244), .A4(new_n275), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT82), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n274), .A2(G244), .A3(new_n275), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT4), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n600), .A2(new_n602), .A3(new_n605), .A4(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n598), .B1(new_n609), .B2(new_n287), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n610), .A2(G200), .ZN(new_n611));
  AOI211_X1 g0411(.A(G190), .B(new_n598), .C1(new_n609), .C2(new_n287), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n595), .B(new_n596), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n274), .A2(G244), .A3(G1698), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n274), .A2(G238), .A3(new_n275), .ZN(new_n615));
  INV_X1    g0415(.A(new_n563), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n287), .ZN(new_n618));
  INV_X1    g0418(.A(new_n490), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n296), .A2(new_n619), .A3(G250), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n296), .A2(G274), .A3(new_n490), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT83), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n622), .B1(new_n620), .B2(new_n621), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n618), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(G200), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n274), .A2(new_n210), .A3(G68), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT19), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n210), .B1(new_n320), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(G87), .B2(new_n207), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n210), .A2(G33), .A3(G97), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n632), .A2(KEYINPUT84), .A3(new_n629), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT84), .B1(new_n632), .B2(new_n629), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n628), .B(new_n631), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n261), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n266), .A2(new_n254), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n512), .A2(G87), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n618), .B(G190), .C1(new_n624), .C2(new_n625), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n627), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n637), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n635), .B2(new_n261), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n254), .B(KEYINPUT85), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n512), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n618), .B(new_n430), .C1(new_n624), .C2(new_n625), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n620), .A2(new_n621), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(KEYINPUT83), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n649), .A2(new_n623), .B1(new_n287), .B2(new_n617), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n646), .B(new_n647), .C1(G169), .C2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n641), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n609), .A2(new_n287), .ZN(new_n653));
  INV_X1    g0453(.A(new_n598), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n310), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AOI211_X1 g0455(.A(new_n430), .B(new_n598), .C1(new_n609), .C2(new_n287), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n593), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n613), .A2(new_n652), .A3(new_n657), .ZN(new_n658));
  NOR4_X1   g0458(.A1(new_n482), .A2(new_n531), .A3(new_n583), .A4(new_n658), .ZN(G372));
  NAND2_X1  g0459(.A1(new_n356), .A2(new_n354), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n326), .A2(new_n329), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n355), .B1(new_n661), .B2(G169), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n358), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n311), .A2(new_n312), .ZN(new_n664));
  INV_X1    g0464(.A(new_n314), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(new_n665), .A3(new_n309), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n663), .B1(new_n666), .B2(new_n349), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n667), .A2(new_n424), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT92), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n429), .A2(new_n669), .A3(new_n433), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT92), .B1(new_n422), .B2(new_n432), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n670), .A2(KEYINPUT18), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT18), .B1(new_n670), .B2(new_n671), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n478), .A2(new_n480), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n462), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT91), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n643), .A2(new_n678), .A3(new_n638), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n678), .B1(new_n643), .B2(new_n638), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n627), .B(new_n640), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n613), .A2(new_n657), .A3(new_n681), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n525), .B(new_n530), .C1(new_n580), .C2(new_n582), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(new_n577), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n610), .A2(G179), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n310), .B2(new_n610), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n595), .A2(new_n596), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n686), .A2(new_n681), .A3(new_n687), .A4(new_n651), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT26), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n652), .A2(KEYINPUT26), .A3(new_n593), .A4(new_n686), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n684), .A2(new_n692), .A3(new_n651), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n677), .B1(new_n482), .B2(new_n694), .ZN(G369));
  NOR2_X1   g0495(.A1(new_n580), .A2(new_n582), .ZN(new_n696));
  AOI221_X4 g0496(.A(new_n535), .B1(new_n549), .B2(new_n551), .C1(new_n579), .C2(new_n575), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n264), .A2(new_n210), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT27), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT27), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n264), .A2(new_n701), .A3(new_n210), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n700), .A2(G213), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G343), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT93), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n698), .B1(new_n580), .B2(new_n706), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(KEYINPUT94), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(KEYINPUT94), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n708), .A2(new_n709), .B1(new_n696), .B2(new_n705), .ZN(new_n710));
  INV_X1    g0510(.A(new_n531), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n705), .A2(new_n517), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n525), .A2(new_n530), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n713), .B1(new_n715), .B2(new_n712), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G330), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n710), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n715), .A2(new_n705), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n708), .A2(new_n709), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n696), .A2(new_n706), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n719), .A2(new_n724), .ZN(G399));
  INV_X1    g0525(.A(new_n213), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G41), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(G1), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n217), .B2(new_n728), .ZN(new_n731));
  XOR2_X1   g0531(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n732));
  XNOR2_X1  g0532(.A(new_n731), .B(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(G330), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n653), .A2(new_n550), .A3(new_n654), .A4(new_n650), .ZN(new_n736));
  OAI211_X1 g0536(.A(G179), .B(new_n487), .C1(new_n494), .C2(new_n495), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n550), .A2(new_n650), .ZN(new_n739));
  INV_X1    g0539(.A(new_n737), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n739), .A2(new_n740), .A3(KEYINPUT30), .A4(new_n610), .ZN(new_n741));
  INV_X1    g0541(.A(new_n610), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n650), .A2(G179), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n742), .A2(new_n743), .A3(new_n496), .A4(new_n548), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n738), .A2(new_n741), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n705), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT31), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n745), .A2(KEYINPUT31), .A3(new_n705), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n658), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n698), .A2(new_n711), .A3(new_n751), .A4(new_n706), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n734), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n641), .A2(new_n651), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n689), .B1(new_n657), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(new_n688), .B2(new_n689), .ZN(new_n756));
  INV_X1    g0556(.A(new_n683), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n577), .A2(new_n657), .A3(new_n613), .A4(new_n681), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n756), .B(new_n651), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(KEYINPUT29), .A3(new_n706), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(KEYINPUT96), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT96), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n759), .A2(new_n762), .A3(KEYINPUT29), .A4(new_n706), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(KEYINPUT29), .B1(new_n693), .B2(new_n706), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n753), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n733), .B1(new_n767), .B2(G1), .ZN(G364));
  INV_X1    g0568(.A(new_n717), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n263), .A2(G20), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n209), .B1(new_n770), .B2(G45), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n727), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(G330), .B2(new_n716), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n219), .B1(G20), .B2(new_n310), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(G20), .A2(G179), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G190), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n274), .B1(new_n781), .B2(new_n267), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n779), .A2(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G190), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n210), .A2(G179), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n786), .A2(new_n307), .A3(G200), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n785), .A2(new_n247), .B1(new_n206), .B2(new_n787), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n778), .A2(new_n307), .A3(G200), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n782), .B(new_n788), .C1(G58), .C2(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n786), .A2(G190), .A3(G200), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT100), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G87), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n786), .A2(new_n780), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n365), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT99), .B(KEYINPUT32), .Z(new_n801));
  NOR3_X1   g0601(.A1(new_n307), .A2(G179), .A3(G200), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n210), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n800), .A2(new_n801), .B1(new_n804), .B2(G97), .ZN(new_n805));
  INV_X1    g0605(.A(new_n801), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n783), .A2(new_n307), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n799), .A2(new_n806), .B1(new_n807), .B2(G50), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n790), .A2(new_n797), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n789), .ZN(new_n810));
  INV_X1    g0610(.A(G322), .ZN(new_n811));
  INV_X1    g0611(.A(G311), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n810), .A2(new_n811), .B1(new_n781), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n798), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n274), .B(new_n813), .C1(G329), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n796), .A2(G303), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n804), .A2(G294), .B1(new_n807), .B2(G326), .ZN(new_n817));
  XNOR2_X1  g0617(.A(KEYINPUT33), .B(G317), .ZN(new_n818));
  INV_X1    g0618(.A(new_n787), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n784), .A2(new_n818), .B1(new_n819), .B2(G283), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n815), .A2(new_n816), .A3(new_n817), .A4(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n777), .B1(new_n809), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(G13), .A2(G33), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(G20), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(new_n776), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT98), .Z(new_n827));
  NAND2_X1  g0627(.A1(new_n389), .A2(new_n391), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n213), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT97), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n218), .A2(new_n489), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n831), .B(new_n832), .C1(new_n489), .C2(new_n251), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n726), .A2(new_n282), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n834), .A2(G355), .B1(new_n502), .B2(new_n726), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n827), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n773), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n822), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n825), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n838), .B1(new_n716), .B2(new_n839), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n775), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G396));
  NAND2_X1  g0642(.A1(new_n693), .A2(new_n706), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n705), .A2(new_n273), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT102), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n666), .A2(new_n308), .A3(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n844), .B(KEYINPUT102), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n315), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n843), .B(new_n850), .Z(new_n851));
  INV_X1    g0651(.A(new_n753), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n773), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n852), .B2(new_n851), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n776), .A2(new_n823), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n837), .B1(new_n267), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n781), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n857), .A2(G159), .B1(G143), .B2(new_n789), .ZN(new_n858));
  INV_X1    g0658(.A(new_n807), .ZN(new_n859));
  INV_X1    g0659(.A(G137), .ZN(new_n860));
  INV_X1    g0660(.A(G150), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n858), .B1(new_n859), .B2(new_n860), .C1(new_n861), .C2(new_n785), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT34), .ZN(new_n863));
  INV_X1    g0663(.A(G132), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n828), .B1(new_n864), .B2(new_n798), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n819), .A2(G68), .ZN(new_n866));
  INV_X1    g0666(.A(G58), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n866), .B1(new_n867), .B2(new_n803), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n865), .B(new_n868), .C1(new_n796), .C2(G50), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n282), .B1(new_n795), .B2(new_n206), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT101), .ZN(new_n871));
  AOI22_X1  g0671(.A1(G311), .A2(new_n814), .B1(new_n857), .B2(G116), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n545), .B2(new_n810), .ZN(new_n873));
  INV_X1    g0673(.A(G283), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n785), .A2(new_n874), .B1(new_n205), .B2(new_n803), .ZN(new_n875));
  INV_X1    g0675(.A(G303), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n859), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n787), .A2(new_n410), .ZN(new_n878));
  NOR4_X1   g0678(.A1(new_n873), .A2(new_n875), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n863), .A2(new_n869), .B1(new_n871), .B2(new_n879), .ZN(new_n880));
  OAI221_X1 g0680(.A(new_n856), .B1(new_n777), .B2(new_n880), .C1(new_n850), .C2(new_n824), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n854), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(G384));
  INV_X1    g0683(.A(new_n587), .ZN(new_n884));
  OR2_X1    g0684(.A1(new_n884), .A2(KEYINPUT35), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(KEYINPUT35), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n885), .A2(G116), .A3(new_n220), .A4(new_n886), .ZN(new_n887));
  XNOR2_X1  g0687(.A(KEYINPUT103), .B(KEYINPUT36), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n887), .B(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n218), .A2(G77), .A3(new_n379), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n246), .B(KEYINPUT104), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n209), .B(G13), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n349), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n358), .A2(new_n705), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n663), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n358), .B(new_n705), .C1(new_n357), .C2(new_n349), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR4_X1   g0698(.A1(new_n583), .A2(new_n658), .A3(new_n531), .A4(new_n705), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n748), .A2(new_n749), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n898), .B(new_n850), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT105), .B1(new_n429), .B2(new_n703), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT105), .ZN(new_n905));
  INV_X1    g0705(.A(new_n703), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n422), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT106), .B1(new_n421), .B2(new_n423), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n399), .A2(new_n404), .A3(new_n420), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT17), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT106), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n422), .A2(KEYINPUT17), .A3(new_n420), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n909), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n908), .B1(new_n674), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n669), .B1(new_n429), .B2(new_n433), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n422), .A2(KEYINPUT92), .A3(new_n432), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n910), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT37), .B1(new_n920), .B2(new_n908), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n429), .A2(new_n433), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT37), .B1(new_n422), .B2(new_n420), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n922), .B(new_n923), .C1(new_n904), .C2(new_n907), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT38), .B1(new_n917), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n923), .A2(new_n922), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n429), .A2(KEYINPUT105), .A3(new_n703), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n905), .B1(new_n422), .B2(new_n906), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n382), .B1(new_n393), .B2(new_n247), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n362), .B1(new_n931), .B2(new_n363), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n398), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n404), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n703), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n433), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n935), .A2(new_n936), .A3(new_n910), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n927), .A2(new_n930), .B1(new_n937), .B2(KEYINPUT37), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n935), .B1(new_n424), .B2(new_n437), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT38), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n903), .B1(new_n926), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n901), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n403), .B1(new_n398), .B2(new_n932), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n910), .B1(new_n432), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n944), .A2(new_n906), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT37), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n924), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT18), .B1(new_n429), .B2(new_n433), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n422), .A2(new_n435), .A3(new_n432), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n912), .A2(new_n914), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n946), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT38), .B1(new_n948), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n943), .B1(new_n941), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n902), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n942), .A2(new_n956), .A3(G330), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n852), .A2(new_n482), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT109), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n942), .A2(new_n956), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n482), .B1(new_n752), .B2(new_n750), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT107), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n357), .A2(new_n358), .A3(new_n706), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n438), .A2(new_n946), .B1(new_n924), .B2(new_n947), .ZN(new_n966));
  AOI21_X1  g0766(.A(KEYINPUT39), .B1(new_n966), .B2(KEYINPUT38), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n909), .B(new_n915), .C1(new_n672), .C2(new_n673), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n968), .A2(new_n908), .B1(new_n921), .B2(new_n924), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n967), .B1(new_n969), .B2(KEYINPUT38), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n940), .B1(new_n938), .B2(new_n939), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n948), .A2(new_n953), .A3(KEYINPUT38), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(KEYINPUT39), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n965), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n898), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n693), .A2(new_n706), .A3(new_n850), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n666), .A2(new_n705), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n976), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n973), .A2(new_n980), .B1(new_n674), .B2(new_n906), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n964), .B1(new_n975), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n916), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n670), .A2(new_n671), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n435), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n670), .A2(new_n671), .A3(KEYINPUT18), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n930), .B1(new_n984), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n985), .A2(new_n930), .A3(new_n910), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n990), .A2(KEYINPUT37), .B1(new_n930), .B2(new_n927), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n940), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n992), .A2(new_n967), .B1(new_n973), .B2(KEYINPUT39), .ZN(new_n993));
  OAI211_X1 g0793(.A(KEYINPUT107), .B(new_n981), .C1(new_n993), .C2(new_n965), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n983), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n482), .A2(new_n765), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n764), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(KEYINPUT108), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT108), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n764), .A2(new_n996), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n677), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n995), .B(new_n1002), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n963), .A2(new_n1003), .B1(new_n209), .B2(new_n770), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n963), .A2(new_n1003), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n893), .B1(new_n1004), .B2(new_n1005), .ZN(G367));
  NAND2_X1  g0806(.A1(new_n681), .A2(new_n651), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n706), .A2(new_n679), .A3(new_n680), .ZN(new_n1008));
  MUX2_X1   g0808(.A(new_n1007), .B(new_n651), .S(new_n1008), .Z(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT110), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(KEYINPUT43), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT112), .Z(new_n1012));
  NAND2_X1  g0812(.A1(new_n687), .A2(new_n705), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n613), .A2(new_n1013), .A3(new_n657), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n686), .A2(new_n687), .A3(new_n705), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(KEYINPUT42), .B1(new_n721), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n657), .B2(new_n705), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1017), .B1(KEYINPUT42), .B2(new_n722), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n723), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1012), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1022), .A2(new_n718), .A3(new_n1016), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT111), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1024), .A2(KEYINPUT43), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(KEYINPUT43), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1010), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1012), .B1(new_n719), .B2(new_n1017), .C1(new_n1019), .C2(new_n1021), .ZN(new_n1028));
  AND3_X1   g0828(.A1(new_n1023), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1027), .B1(new_n1023), .B2(new_n1028), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n727), .B(KEYINPUT41), .Z(new_n1032));
  INV_X1    g0832(.A(KEYINPUT45), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n723), .B2(new_n1017), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  NOR3_X1   g0835(.A1(new_n723), .A2(new_n1033), .A3(new_n1017), .ZN(new_n1036));
  AOI21_X1  g0836(.A(KEYINPUT44), .B1(new_n723), .B2(new_n1017), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT44), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1038), .B(new_n1016), .C1(new_n721), .C2(new_n722), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n1035), .A2(new_n1036), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n718), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n724), .A2(KEYINPUT45), .A3(new_n1016), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n1034), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1042), .A2(new_n719), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT113), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n720), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n710), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n721), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1046), .B1(new_n710), .B2(new_n1047), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n769), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1050), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1052), .A2(new_n717), .A3(new_n721), .A4(new_n1048), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1041), .A2(new_n767), .A3(new_n1045), .A4(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1032), .B1(new_n1055), .B2(new_n767), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1031), .B1(new_n1056), .B2(new_n772), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n827), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n831), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1058), .B1(new_n213), .B2(new_n254), .C1(new_n1059), .C2(new_n237), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1060), .A2(new_n773), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n810), .A2(new_n861), .B1(new_n781), .B2(new_n202), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n282), .B(new_n1062), .C1(G137), .C2(new_n814), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n796), .A2(G58), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G143), .A2(new_n807), .B1(new_n819), .B2(G77), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n804), .A2(G68), .B1(new_n784), .B2(G159), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n796), .A2(G116), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT46), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1068), .A2(new_n1069), .B1(G294), .B2(new_n784), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n1069), .B2(new_n1068), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT114), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n814), .A2(G317), .B1(new_n789), .B2(G303), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n874), .B2(new_n781), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n859), .A2(new_n812), .B1(new_n206), .B2(new_n803), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n787), .A2(new_n205), .ZN(new_n1077));
  NOR4_X1   g0877(.A1(new_n1075), .A2(new_n1076), .A3(new_n828), .A4(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1067), .B1(new_n1073), .B2(new_n1079), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT47), .Z(new_n1081));
  OAI221_X1 g0881(.A(new_n1061), .B1(new_n1081), .B2(new_n777), .C1(new_n1010), .C2(new_n839), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1057), .A2(new_n1082), .ZN(G387));
  AOI22_X1  g0883(.A1(new_n857), .A2(G303), .B1(G317), .B2(new_n789), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1084), .B1(new_n859), .B2(new_n811), .C1(new_n812), .C2(new_n785), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT48), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n796), .A2(G294), .B1(G283), .B2(new_n804), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT49), .Z(new_n1091));
  AOI21_X1  g0891(.A(new_n828), .B1(G326), .B2(new_n814), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n502), .B2(new_n787), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n644), .A2(new_n804), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n814), .A2(G150), .B1(new_n789), .B2(G50), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(new_n247), .C2(new_n781), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n795), .A2(new_n267), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n828), .B1(new_n205), .B2(new_n787), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n401), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1100), .A2(new_n785), .B1(new_n859), .B2(new_n365), .ZN(new_n1101));
  NOR4_X1   g0901(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .A4(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n776), .B1(new_n1094), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n729), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n834), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(G107), .B2(new_n213), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n241), .A2(G45), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT115), .Z(new_n1108));
  NOR2_X1   g0908(.A1(new_n258), .A2(G50), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT50), .ZN(new_n1110));
  AOI211_X1 g0910(.A(G45), .B(new_n1104), .C1(G68), .C2(G77), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1059), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1106), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1103), .B(new_n773), .C1(new_n827), .C2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT116), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n710), .B2(new_n825), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n1054), .B2(new_n772), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1054), .A2(new_n767), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n727), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1054), .A2(new_n767), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1117), .B1(new_n1119), .B2(new_n1120), .ZN(G393));
  NOR2_X1   g0921(.A1(new_n1040), .A2(new_n718), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n719), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1017), .A2(new_n825), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n804), .A2(G116), .B1(G294), .B2(new_n857), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n876), .B2(new_n785), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1127), .B(KEYINPUT117), .Z(new_n1128));
  AOI22_X1  g0928(.A1(new_n807), .A2(G317), .B1(G311), .B2(new_n789), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT52), .Z(new_n1130));
  OAI221_X1 g0930(.A(new_n282), .B1(new_n798), .B2(new_n811), .C1(new_n206), .C2(new_n787), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n796), .B2(G283), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1128), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n807), .A2(G150), .B1(G159), .B2(new_n789), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT51), .Z(new_n1135));
  NOR2_X1   g0935(.A1(new_n803), .A2(new_n267), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n878), .B(new_n1136), .C1(G50), .C2(new_n784), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n796), .A2(new_n222), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n781), .A2(new_n258), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1139), .B(new_n829), .C1(G143), .C2(new_n814), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1135), .A2(new_n1137), .A3(new_n1138), .A4(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n777), .B1(new_n1133), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n831), .A2(new_n245), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n827), .B1(G97), .B2(new_n726), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n837), .B(new_n1142), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1124), .A2(new_n772), .B1(new_n1125), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1118), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1147), .A2(new_n727), .A3(new_n1055), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(G390));
  INV_X1    g0949(.A(new_n965), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n970), .B(new_n974), .C1(new_n1150), .C2(new_n980), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n965), .B(KEYINPUT118), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n759), .A2(new_n706), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n978), .B1(new_n1153), .B2(new_n850), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1152), .B1(new_n1154), .B2(new_n976), .C1(new_n926), .C2(new_n941), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n753), .A2(new_n850), .A3(new_n898), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1151), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(new_n772), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n993), .A2(new_n823), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n837), .B1(new_n1100), .B2(new_n855), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n796), .A2(G150), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT53), .ZN(new_n1165));
  INV_X1    g0965(.A(G128), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n859), .A2(new_n1166), .B1(new_n202), .B2(new_n787), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G159), .B2(new_n804), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT54), .B(G143), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n785), .A2(new_n860), .B1(new_n781), .B2(new_n1169), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n1170), .A2(KEYINPUT120), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n274), .B1(new_n810), .B2(new_n864), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G125), .B2(new_n814), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1170), .A2(KEYINPUT120), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1168), .A2(new_n1171), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1165), .A2(new_n1175), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n282), .B1(new_n781), .B2(new_n205), .C1(new_n545), .C2(new_n798), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n866), .B1(new_n859), .B2(new_n874), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(G107), .C2(new_n784), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n803), .A2(new_n267), .B1(new_n810), .B2(new_n502), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1180), .A2(KEYINPUT121), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(KEYINPUT121), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n797), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1176), .B1(new_n1179), .B2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1162), .B(new_n1163), .C1(new_n777), .C2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1161), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT122), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n850), .B(G330), .C1(new_n899), .C2(new_n900), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n976), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1157), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT119), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n977), .A2(new_n979), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1154), .A2(new_n1157), .A3(new_n1190), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1192), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n764), .A2(new_n996), .A3(new_n999), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n999), .B1(new_n764), .B2(new_n996), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n677), .B(new_n958), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1159), .A2(new_n1198), .A3(new_n1202), .A4(new_n1160), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n1151), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1157), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n1204), .A2(new_n1205), .B1(new_n1206), .B2(new_n1201), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1203), .A2(new_n1207), .A3(new_n727), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1161), .A2(KEYINPUT122), .A3(new_n1185), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1188), .A2(new_n1208), .A3(new_n1209), .ZN(G378));
  INV_X1    g1010(.A(KEYINPUT125), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1201), .A2(new_n1211), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1001), .A2(KEYINPUT125), .A3(new_n677), .A4(new_n958), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1203), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n676), .A2(new_n458), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n453), .A2(new_n455), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n703), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT55), .Z(new_n1219));
  NAND2_X1  g1019(.A1(new_n1216), .A2(new_n1219), .ZN(new_n1220));
  XOR2_X1   g1020(.A(KEYINPUT124), .B(KEYINPUT56), .Z(new_n1221));
  INV_X1    g1021(.A(new_n1219), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n676), .A2(new_n458), .A3(new_n1222), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1220), .A2(new_n1221), .A3(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1221), .B1(new_n1220), .B2(new_n1223), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n957), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1226), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1228), .A2(new_n942), .A3(G330), .A4(new_n956), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n995), .A2(new_n1230), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n983), .A2(new_n1227), .A3(new_n994), .A4(new_n1229), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1215), .A2(new_n1233), .A3(KEYINPUT57), .ZN(new_n1234));
  AND4_X1   g1034(.A1(new_n983), .A2(new_n1227), .A3(new_n994), .A4(new_n1229), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n983), .A2(new_n994), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1206), .A2(new_n1201), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1238), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1237), .A2(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n727), .B(new_n1234), .C1(new_n1242), .C2(KEYINPUT57), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n295), .B1(new_n798), .B2(new_n874), .C1(new_n810), .C2(new_n206), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n828), .B(new_n1244), .C1(G68), .C2(new_n804), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n644), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1245), .B1(new_n1246), .B2(new_n781), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(G116), .A2(new_n807), .B1(new_n819), .B2(G58), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n205), .B2(new_n785), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1247), .A2(new_n1098), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT58), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n295), .B1(new_n829), .B2(new_n278), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n202), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n807), .A2(G125), .B1(G128), .B2(new_n789), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n861), .B2(new_n803), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n784), .A2(G132), .B1(new_n857), .B2(G137), .ZN(new_n1257));
  XOR2_X1   g1057(.A(new_n1257), .B(KEYINPUT123), .Z(new_n1258));
  INV_X1    g1058(.A(new_n1169), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n1256), .B(new_n1258), .C1(new_n796), .C2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(KEYINPUT59), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n819), .A2(G159), .ZN(new_n1263));
  AOI211_X1 g1063(.A(G33), .B(G41), .C1(new_n814), .C2(G124), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1261), .A2(KEYINPUT59), .ZN(new_n1266));
  OAI221_X1 g1066(.A(new_n1254), .B1(KEYINPUT58), .B2(new_n1250), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n776), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n837), .B1(new_n202), .B2(new_n855), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1268), .B(new_n1269), .C1(new_n1226), .C2(new_n824), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(new_n1233), .B2(new_n772), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1243), .A2(new_n1272), .ZN(G375));
  OAI22_X1  g1073(.A1(new_n859), .A2(new_n864), .B1(new_n202), .B2(new_n803), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(new_n784), .B2(new_n1259), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n796), .A2(G159), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n798), .A2(new_n1166), .B1(new_n781), .B2(new_n861), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(G137), .B2(new_n789), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n829), .B1(G58), .B2(new_n819), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1275), .A2(new_n1276), .A3(new_n1278), .A4(new_n1279), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n859), .A2(new_n545), .B1(new_n267), .B2(new_n787), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(G116), .B2(new_n784), .ZN(new_n1282));
  OAI22_X1  g1082(.A1(new_n810), .A2(new_n874), .B1(new_n781), .B2(new_n206), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n274), .B(new_n1283), .C1(G303), .C2(new_n814), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1282), .A2(new_n1284), .A3(new_n1095), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n795), .A2(new_n205), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1280), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n776), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n837), .B1(new_n247), .B2(new_n855), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1288), .B(new_n1289), .C1(new_n898), .C2(new_n824), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1290), .B1(new_n1206), .B2(new_n771), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1240), .A2(new_n1032), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1206), .A2(new_n1201), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1291), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(G381));
  NOR4_X1   g1095(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1057), .A2(new_n1082), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1208), .A2(new_n1161), .A3(new_n1185), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1296), .A2(new_n1297), .A3(new_n1294), .A4(new_n1298), .ZN(new_n1299));
  OR2_X1    g1099(.A1(new_n1299), .A2(G375), .ZN(G407));
  INV_X1    g1100(.A(G343), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(G213), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1243), .A2(new_n1272), .A3(new_n1298), .A4(new_n1303), .ZN(new_n1304));
  OAI211_X1 g1104(.A(G213), .B(new_n1304), .C1(new_n1299), .C2(G375), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT126), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1305), .B(new_n1306), .ZN(G409));
  XNOR2_X1  g1107(.A(G393), .B(new_n841), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1057), .A2(new_n1082), .A3(G390), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G390), .B1(new_n1057), .B2(new_n1082), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1309), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(G390), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(G387), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1057), .A2(G390), .A3(new_n1082), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1314), .A2(new_n1308), .A3(new_n1315), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1312), .A2(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(KEYINPUT57), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n727), .B1(new_n1318), .B2(new_n1241), .ZN(new_n1319));
  AOI21_X1  g1119(.A(KEYINPUT57), .B1(new_n1215), .B2(new_n1233), .ZN(new_n1320));
  OAI211_X1 g1120(.A(G378), .B(new_n1272), .C1(new_n1319), .C2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1032), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1215), .A2(new_n1233), .A3(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1270), .B1(new_n1237), .B2(new_n771), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1298), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1321), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1302), .ZN(new_n1327));
  OAI21_X1  g1127(.A(KEYINPUT60), .B1(new_n1206), .B2(new_n1201), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(new_n1293), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1206), .A2(KEYINPUT60), .A3(new_n1201), .ZN(new_n1330));
  AND3_X1   g1130(.A1(new_n1329), .A2(new_n727), .A3(new_n1330), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n882), .B1(new_n1331), .B2(new_n1291), .ZN(new_n1332));
  AND2_X1   g1132(.A1(new_n1330), .A2(new_n727), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1291), .B1(new_n1333), .B2(new_n1329), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(G384), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1303), .A2(G2897), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1332), .A2(new_n1335), .A3(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1336), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1334), .A2(G384), .ZN(new_n1339));
  AOI211_X1 g1139(.A(new_n882), .B(new_n1291), .C1(new_n1333), .C2(new_n1329), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1338), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  AND2_X1   g1141(.A1(new_n1337), .A2(new_n1341), .ZN(new_n1342));
  AOI21_X1  g1142(.A(KEYINPUT61), .B1(new_n1327), .B2(new_n1342), .ZN(new_n1343));
  XNOR2_X1  g1143(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1344), .B1(new_n1327), .B2(new_n1346), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1303), .B1(new_n1321), .B2(new_n1325), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1348), .A2(KEYINPUT63), .A3(new_n1345), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1317), .A2(new_n1343), .A3(new_n1347), .A4(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT62), .ZN(new_n1351));
  AND3_X1   g1151(.A1(new_n1348), .A2(new_n1351), .A3(new_n1345), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT61), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1337), .A2(new_n1341), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1353), .B1(new_n1348), .B2(new_n1354), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1351), .B1(new_n1348), .B2(new_n1345), .ZN(new_n1356));
  NOR3_X1   g1156(.A1(new_n1352), .A2(new_n1355), .A3(new_n1356), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1350), .B1(new_n1357), .B2(new_n1317), .ZN(G405));
  NAND2_X1  g1158(.A1(G375), .A2(new_n1298), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1359), .A2(new_n1321), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1360), .A2(new_n1345), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1359), .A2(new_n1346), .A3(new_n1321), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(new_n1317), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1363), .A2(new_n1364), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1317), .A2(new_n1361), .A3(new_n1362), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1365), .A2(new_n1366), .ZN(G402));
endmodule


