//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0 1 1 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1329,
    new_n1330, new_n1331, new_n1332;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  INV_X1    g0003(.A(G87), .ZN(new_n204));
  INV_X1    g0004(.A(G250), .ZN(new_n205));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G257), .ZN(new_n207));
  OAI22_X1  g0007(.A1(new_n204), .A2(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  AOI21_X1  g0008(.A(new_n208), .B1(G68), .B2(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G107), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n203), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n203), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT0), .Z(new_n226));
  NOR2_X1   g0026(.A1(G58), .A2(G68), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n223), .A2(new_n226), .A3(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n220), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n211), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G270), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT64), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n253));
  AND2_X1   g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G222), .ZN(new_n256));
  INV_X1    g0056(.A(G223), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n254), .B(new_n256), .C1(new_n257), .C2(new_n255), .ZN(new_n258));
  INV_X1    g0058(.A(new_n231), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n258), .B(new_n262), .C1(G77), .C2(new_n254), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n265));
  INV_X1    g0065(.A(G274), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n231), .B1(KEYINPUT65), .B2(new_n260), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT65), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G33), .A3(G41), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n265), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n263), .B(new_n268), .C1(new_n215), .C2(new_n273), .ZN(new_n274));
  OR2_X1    g0074(.A1(new_n274), .A2(G179), .ZN(new_n275));
  OAI21_X1  g0075(.A(G20), .B1(new_n228), .B2(G50), .ZN(new_n276));
  INV_X1    g0076(.A(G150), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n252), .A2(G20), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  OAI221_X1 g0082(.A(new_n276), .B1(new_n277), .B2(new_n279), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n231), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n285), .B1(new_n264), .B2(G20), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n283), .A2(new_n285), .B1(G50), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G13), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(G1), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G20), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n287), .B1(G50), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G169), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n274), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n275), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n274), .A2(G200), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT9), .ZN(new_n298));
  OAI221_X1 g0098(.A(new_n296), .B1(new_n297), .B2(new_n274), .C1(new_n298), .C2(new_n291), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(new_n298), .B2(new_n291), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT10), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n301), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n295), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT75), .B1(new_n250), .B2(G33), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT75), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(new_n252), .A3(KEYINPUT3), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n305), .A2(new_n307), .B1(new_n250), .B2(G33), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n257), .A2(new_n255), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n215), .A2(G1698), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G87), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n261), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n268), .B1(new_n273), .B2(new_n220), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT78), .ZN(new_n315));
  NOR4_X1   g0115(.A1(new_n313), .A2(new_n314), .A3(new_n315), .A4(G179), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n292), .B1(new_n313), .B2(new_n314), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT78), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n313), .A2(new_n314), .ZN(new_n319));
  INV_X1    g0119(.A(G179), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n316), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n305), .A2(new_n307), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n251), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT7), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(new_n325), .A3(new_n230), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT7), .B1(new_n308), .B2(G20), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n327), .A3(G68), .ZN(new_n328));
  XNOR2_X1  g0128(.A(G58), .B(G68), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n329), .A2(G20), .B1(G159), .B2(new_n278), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(KEYINPUT16), .A3(new_n330), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G68), .ZN(new_n334));
  NAND2_X1  g0134(.A1(KEYINPUT77), .A2(KEYINPUT7), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n254), .B2(G20), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n251), .A2(new_n253), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT77), .B(KEYINPUT7), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(new_n338), .A3(new_n230), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n334), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n330), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n333), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n331), .A2(new_n342), .A3(new_n285), .ZN(new_n343));
  INV_X1    g0143(.A(new_n282), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(new_n290), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(new_n286), .B2(new_n344), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n322), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT79), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT18), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(KEYINPUT79), .A2(KEYINPUT18), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n348), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n322), .A2(new_n349), .A3(new_n350), .A4(new_n347), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(G200), .B1(new_n313), .B2(new_n314), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n319), .A2(G190), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n343), .A2(new_n356), .A3(new_n357), .A4(new_n346), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT17), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT80), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT80), .ZN(new_n361));
  INV_X1    g0161(.A(new_n358), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n362), .A2(KEYINPUT17), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT17), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n358), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n361), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n355), .B1(new_n360), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G200), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n337), .A2(new_n220), .A3(G1698), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n369), .B(KEYINPUT66), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n337), .A2(G107), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n254), .A2(G238), .A3(G1698), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT67), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT67), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n370), .A2(new_n375), .A3(new_n371), .A4(new_n372), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n262), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n273), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n267), .B1(new_n378), .B2(G244), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n368), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n285), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n282), .B(KEYINPUT68), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n278), .ZN(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT15), .B(G87), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n385), .A2(new_n280), .B1(G20), .B2(G77), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n381), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n286), .A2(G77), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n290), .A2(G77), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n377), .A2(new_n379), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n390), .B1(new_n391), .B2(new_n297), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n304), .B(new_n367), .C1(new_n380), .C2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G41), .ZN(new_n394));
  AND2_X1   g0194(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n395));
  NOR2_X1   g0195(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n394), .A2(KEYINPUT5), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G45), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n401), .A2(G1), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n272), .B(G270), .C1(new_n400), .C2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT87), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n397), .A2(new_n399), .B1(new_n269), .B2(new_n271), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n402), .B1(new_n269), .B2(new_n271), .ZN(new_n408));
  OAI211_X1 g0208(.A(KEYINPUT87), .B(G270), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n207), .A2(new_n255), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n211), .A2(G1698), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n323), .A2(new_n251), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n337), .A2(G303), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n402), .A2(G274), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n400), .B2(KEYINPUT83), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT83), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n397), .A2(new_n418), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n262), .A2(new_n415), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n410), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G33), .A2(G283), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n422), .B(new_n230), .C1(G33), .C2(new_n206), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n423), .B(new_n285), .C1(new_n230), .C2(G116), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT20), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT88), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n230), .A2(G116), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n381), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT88), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n428), .A2(new_n429), .A3(KEYINPUT20), .A4(new_n423), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n424), .A2(new_n425), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n426), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n289), .A2(new_n427), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n264), .A2(G33), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n381), .A2(new_n290), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G116), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n432), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n421), .A2(G169), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT21), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n421), .A2(KEYINPUT21), .A3(new_n438), .A4(G169), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n438), .A2(G179), .A3(new_n420), .A4(new_n410), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n438), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n410), .A2(G190), .A3(new_n420), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n368), .B1(new_n410), .B2(new_n420), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT89), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n448), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT89), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n450), .A2(new_n451), .A3(new_n445), .A4(new_n446), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n444), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT92), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n260), .A2(KEYINPUT65), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n455), .A2(new_n271), .A3(new_n259), .ZN(new_n456));
  XNOR2_X1  g0256(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n398), .B1(new_n457), .B2(new_n394), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n456), .B1(new_n458), .B2(new_n402), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G257), .A2(G1698), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(new_n205), .B2(G1698), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n306), .B1(KEYINPUT3), .B2(new_n252), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n250), .A2(KEYINPUT75), .A3(G33), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n251), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G294), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n459), .A2(G264), .B1(new_n466), .B2(new_n262), .ZN(new_n467));
  INV_X1    g0267(.A(new_n416), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n419), .B(new_n468), .C1(new_n458), .C2(new_n418), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n454), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n466), .A2(new_n262), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n272), .B(G264), .C1(new_n400), .C2(new_n403), .ZN(new_n472));
  AND4_X1   g0272(.A1(new_n454), .A2(new_n471), .A3(new_n472), .A4(new_n469), .ZN(new_n473));
  OAI21_X1  g0273(.A(G169), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n471), .A2(new_n472), .A3(new_n469), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(new_n320), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n289), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n210), .A2(G20), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT25), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT25), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n289), .A2(new_n481), .A3(G20), .A4(new_n210), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n480), .B(new_n482), .C1(new_n435), .C2(new_n210), .ZN(new_n483));
  XNOR2_X1  g0283(.A(new_n483), .B(KEYINPUT91), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT22), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(new_n204), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n323), .A2(new_n230), .A3(new_n251), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n230), .A2(G87), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n485), .B1(new_n337), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT23), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n479), .B(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n230), .A2(G33), .A3(G116), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT90), .ZN(new_n494));
  XNOR2_X1  g0294(.A(new_n493), .B(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n490), .A2(KEYINPUT24), .A3(new_n492), .A4(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n487), .A2(new_n495), .A3(new_n492), .A4(new_n489), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT24), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n496), .A2(new_n285), .A3(new_n499), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n474), .A2(new_n477), .B1(new_n484), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n484), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n467), .A2(new_n454), .A3(new_n469), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n475), .A2(KEYINPUT92), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n503), .A2(new_n504), .A3(new_n297), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n475), .A2(new_n368), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT93), .B1(new_n501), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n505), .A2(new_n506), .ZN(new_n509));
  INV_X1    g0309(.A(new_n502), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT93), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n292), .B1(new_n503), .B2(new_n504), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n502), .B1(new_n513), .B2(new_n476), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n511), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n217), .A2(G1698), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n323), .A2(new_n251), .A3(new_n516), .ZN(new_n517));
  XOR2_X1   g0317(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n516), .A2(KEYINPUT4), .B1(G250), .B2(G1698), .ZN(new_n520));
  OR2_X1    g0320(.A1(new_n520), .A2(new_n337), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n521), .A3(new_n422), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n262), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n272), .B(G257), .C1(new_n400), .C2(new_n403), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n469), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n523), .A2(new_n526), .A3(new_n320), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT85), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n523), .A2(new_n526), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n292), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n210), .B1(new_n336), .B2(new_n339), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT6), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n533), .A2(new_n206), .A3(G107), .ZN(new_n534));
  XNOR2_X1  g0334(.A(G97), .B(G107), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n534), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n536), .A2(new_n230), .B1(new_n216), .B2(new_n279), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n285), .B1(new_n532), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n436), .A2(G97), .ZN(new_n539));
  INV_X1    g0339(.A(new_n290), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n206), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n523), .A2(new_n526), .A3(KEYINPUT85), .A4(new_n320), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n529), .A2(new_n531), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n422), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n545), .B1(new_n517), .B2(new_n518), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n261), .B1(new_n546), .B2(new_n521), .ZN(new_n547));
  OAI21_X1  g0347(.A(G200), .B1(new_n547), .B2(new_n525), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT84), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n523), .A2(new_n526), .A3(G190), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT84), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n552), .B(G200), .C1(new_n547), .C2(new_n525), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n549), .A2(new_n550), .A3(new_n551), .A4(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n308), .A2(new_n230), .A3(G68), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT19), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n280), .A2(new_n556), .A3(G97), .ZN(new_n557));
  NOR2_X1   g0357(.A1(G97), .A2(G107), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G33), .A2(G97), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n558), .A2(new_n204), .B1(new_n559), .B2(new_n230), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n557), .B1(new_n560), .B2(new_n556), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n285), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n540), .A2(new_n384), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n436), .A2(new_n385), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n468), .B1(new_n408), .B2(G250), .ZN(new_n567));
  NOR2_X1   g0367(.A1(G238), .A2(G1698), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n568), .B1(new_n217), .B2(G1698), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n308), .A2(new_n569), .B1(G33), .B2(G116), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n567), .B1(new_n570), .B2(new_n261), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n292), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n567), .B(new_n320), .C1(new_n570), .C2(new_n261), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n566), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n571), .A2(G200), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n562), .A2(new_n285), .B1(new_n540), .B2(new_n384), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n567), .B(G190), .C1(new_n570), .C2(new_n261), .ZN(new_n577));
  OR3_X1    g0377(.A1(new_n435), .A2(KEYINPUT86), .A3(new_n204), .ZN(new_n578));
  OAI21_X1  g0378(.A(KEYINPUT86), .B1(new_n435), .B2(new_n204), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n575), .A2(new_n576), .A3(new_n577), .A4(new_n580), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n574), .A2(new_n581), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n544), .A2(new_n554), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n453), .A2(new_n508), .A3(new_n515), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(KEYINPUT74), .A2(KEYINPUT14), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n215), .A2(new_n255), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n220), .A2(G1698), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n251), .A2(new_n586), .A3(new_n253), .A4(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT69), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n588), .A2(new_n589), .A3(new_n559), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n589), .B1(new_n588), .B2(new_n559), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n590), .A2(new_n591), .A3(new_n261), .ZN(new_n592));
  INV_X1    g0392(.A(G238), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n268), .B1(new_n273), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(KEYINPUT13), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT71), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n594), .ZN(new_n598));
  INV_X1    g0398(.A(new_n591), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n588), .A2(new_n589), .A3(new_n559), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n262), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT13), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n598), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT70), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n598), .A2(new_n601), .A3(KEYINPUT70), .A4(new_n602), .ZN(new_n606));
  OAI211_X1 g0406(.A(KEYINPUT71), .B(KEYINPUT13), .C1(new_n592), .C2(new_n594), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n597), .A2(new_n605), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n585), .B1(new_n608), .B2(G169), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n595), .A2(new_n603), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(G179), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n608), .A2(G169), .A3(new_n585), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n280), .A2(G77), .B1(new_n278), .B2(G50), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n230), .B2(G68), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n285), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT11), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n617), .A2(new_n618), .B1(G68), .B2(new_n286), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n618), .B2(new_n617), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT73), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n540), .A2(new_n621), .A3(new_n334), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT12), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n621), .B1(new_n540), .B2(new_n334), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n623), .B(new_n624), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n614), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n608), .A2(G200), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n595), .A2(new_n603), .A3(G190), .ZN(new_n629));
  XNOR2_X1  g0429(.A(new_n629), .B(KEYINPUT72), .ZN(new_n630));
  OR3_X1    g0430(.A1(new_n628), .A2(new_n630), .A3(new_n626), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n391), .A2(G179), .ZN(new_n632));
  AOI21_X1  g0432(.A(G169), .B1(new_n377), .B2(new_n379), .ZN(new_n633));
  OR3_X1    g0433(.A1(new_n632), .A2(new_n390), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n627), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n393), .A2(new_n584), .A3(new_n635), .ZN(G372));
  INV_X1    g0436(.A(KEYINPUT95), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n322), .A2(new_n637), .A3(new_n347), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n637), .B1(new_n322), .B2(new_n347), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n350), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n348), .A2(KEYINPUT95), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n322), .A2(new_n637), .A3(new_n347), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(KEYINPUT18), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n628), .A2(new_n630), .A3(new_n626), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n627), .B1(new_n645), .B2(new_n634), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n360), .A2(new_n366), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n644), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n302), .A2(new_n303), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n294), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n393), .A2(new_n635), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT94), .ZN(new_n654));
  OR3_X1    g0454(.A1(new_n570), .A2(new_n654), .A3(new_n261), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n654), .B1(new_n570), .B2(new_n261), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n567), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(G200), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n576), .A2(new_n580), .ZN(new_n660));
  INV_X1    g0460(.A(new_n571), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n660), .B1(G190), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n511), .B(new_n554), .C1(new_n444), .C2(new_n501), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n665), .B1(new_n666), .B2(new_n544), .ZN(new_n667));
  INV_X1    g0467(.A(new_n582), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT26), .B1(new_n668), .B2(new_n544), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n658), .A2(new_n292), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n670), .A2(new_n573), .A3(new_n566), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n653), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n652), .A2(new_n674), .ZN(G369));
  NAND2_X1  g0475(.A1(new_n508), .A2(new_n515), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  OR3_X1    g0477(.A1(new_n478), .A2(KEYINPUT27), .A3(G20), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT27), .B1(new_n478), .B2(G20), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n677), .B1(new_n510), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n501), .A2(new_n682), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n445), .A2(new_n683), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n444), .A2(new_n687), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n449), .A2(new_n452), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n688), .B1(new_n691), .B2(new_n687), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT96), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n692), .A2(new_n693), .A3(G330), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n693), .B1(new_n692), .B2(G330), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n686), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n508), .A2(new_n515), .A3(new_n444), .A4(new_n683), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n501), .A2(new_n683), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n696), .A2(new_n700), .ZN(G399));
  INV_X1    g0501(.A(new_n224), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G41), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G1), .ZN(new_n705));
  INV_X1    g0505(.A(G116), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n558), .A2(new_n204), .A3(new_n706), .ZN(new_n707));
  OAI22_X1  g0507(.A1(new_n705), .A2(new_n707), .B1(new_n229), .B2(new_n704), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT97), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT28), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n664), .B1(new_n668), .B2(new_n544), .ZN(new_n711));
  INV_X1    g0511(.A(new_n544), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT26), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n671), .A2(new_n663), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n711), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  XOR2_X1   g0515(.A(new_n671), .B(KEYINPUT100), .Z(new_n716));
  NAND2_X1  g0516(.A1(new_n689), .A2(new_n514), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n671), .A2(new_n663), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n717), .A2(new_n511), .A3(new_n554), .A4(new_n718), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n715), .B(new_n716), .C1(new_n719), .C2(new_n712), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT29), .B1(new_n721), .B2(new_n682), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n410), .A2(new_n420), .A3(G179), .A4(new_n467), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n661), .A2(new_n523), .A3(new_n526), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT98), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI211_X1 g0528(.A(KEYINPUT98), .B(new_n723), .C1(new_n724), .C2(new_n725), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(G179), .B1(new_n657), .B2(new_n567), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(new_n475), .A3(new_n530), .A4(new_n421), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n724), .A2(new_n725), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT30), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n682), .B1(new_n730), .B2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT31), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n726), .ZN(new_n739));
  OAI211_X1 g0539(.A(KEYINPUT31), .B(new_n682), .C1(new_n735), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(KEYINPUT99), .B1(new_n584), .B2(new_n682), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n583), .A2(new_n689), .A3(new_n690), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT99), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n677), .A2(new_n743), .A3(new_n744), .A4(new_n683), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n741), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G330), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n673), .A2(new_n683), .ZN(new_n748));
  OAI221_X1 g0548(.A(new_n722), .B1(new_n746), .B2(new_n747), .C1(KEYINPUT29), .C2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n710), .B1(new_n750), .B2(G1), .ZN(G364));
  NOR2_X1   g0551(.A1(new_n694), .A2(new_n695), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n288), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n705), .B1(G45), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n752), .B(new_n755), .C1(G330), .C2(new_n692), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n692), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n702), .A2(new_n337), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G355), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n248), .A2(new_n401), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n308), .A2(new_n702), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(G45), .B2(new_n229), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n763), .B1(G116), .B2(new_n224), .C1(new_n764), .C2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n231), .B1(G20), .B2(new_n292), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n759), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n320), .A2(new_n368), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n230), .A2(new_n297), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n214), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G179), .A2(G200), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G190), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n206), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n320), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n772), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n337), .B(new_n779), .C1(G58), .C2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n368), .A2(G179), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n772), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G87), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n230), .A2(G190), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n784), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n210), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n788), .A2(new_n780), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n790), .B1(G77), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n788), .A2(new_n775), .ZN(new_n794));
  INV_X1    g0594(.A(G159), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT32), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n783), .A2(new_n787), .A3(new_n793), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n771), .A2(new_n788), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n774), .B(new_n798), .C1(G68), .C2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G317), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(KEYINPUT33), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n802), .A2(KEYINPUT33), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n800), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n794), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G329), .ZN(new_n807));
  INV_X1    g0607(.A(G283), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n805), .B(new_n807), .C1(new_n808), .C2(new_n789), .ZN(new_n809));
  INV_X1    g0609(.A(new_n773), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(G326), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n786), .A2(G303), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n254), .B1(new_n782), .B2(G322), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n777), .A2(G294), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n811), .A2(new_n812), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(G311), .B2(new_n792), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n768), .B1(new_n801), .B2(new_n816), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n761), .A2(new_n770), .A3(new_n754), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n756), .A2(new_n818), .ZN(G396));
  NOR4_X1   g0619(.A1(new_n632), .A2(new_n633), .A3(new_n390), .A4(new_n682), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n392), .A2(new_n380), .B1(new_n390), .B2(new_n683), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n820), .B1(new_n634), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n748), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n822), .B(new_n683), .C1(new_n672), .C2(new_n667), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n742), .A2(new_n745), .ZN(new_n827));
  INV_X1    g0627(.A(new_n741), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n747), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n826), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n755), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n768), .A2(new_n757), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n755), .B1(new_n216), .B2(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT101), .Z(new_n834));
  AOI21_X1  g0634(.A(new_n779), .B1(G303), .B2(new_n810), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n706), .B2(new_n791), .ZN(new_n836));
  INV_X1    g0636(.A(new_n789), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G87), .A2(new_n837), .B1(new_n806), .B2(G311), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n808), .B2(new_n799), .ZN(new_n839));
  NOR3_X1   g0639(.A1(new_n836), .A2(new_n254), .A3(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(G294), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n840), .B1(new_n210), .B2(new_n785), .C1(new_n841), .C2(new_n781), .ZN(new_n842));
  AOI22_X1  g0642(.A1(G143), .A2(new_n782), .B1(new_n792), .B2(G159), .ZN(new_n843));
  INV_X1    g0643(.A(G137), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n843), .B1(new_n844), .B2(new_n773), .C1(new_n277), .C2(new_n799), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT34), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n777), .A2(G58), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n837), .A2(G68), .ZN(new_n849));
  INV_X1    g0649(.A(G132), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n785), .A2(new_n214), .B1(new_n794), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n851), .A2(new_n324), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n847), .A2(new_n848), .A3(new_n849), .A4(new_n852), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n845), .A2(new_n846), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n842), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT102), .ZN(new_n856));
  INV_X1    g0656(.A(new_n768), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n834), .B1(new_n856), .B2(new_n857), .C1(new_n822), .C2(new_n758), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n831), .A2(new_n858), .ZN(G384));
  XNOR2_X1  g0659(.A(new_n736), .B(new_n737), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n745), .B2(new_n742), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n626), .A2(new_n682), .ZN(new_n862));
  INV_X1    g0662(.A(new_n613), .ZN(new_n863));
  INV_X1    g0663(.A(new_n612), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n863), .A2(new_n609), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n626), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n631), .B(new_n862), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n626), .B(new_n682), .C1(new_n614), .C2(new_n645), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR4_X1   g0669(.A1(new_n861), .A2(new_n869), .A3(KEYINPUT40), .A4(new_n823), .ZN(new_n870));
  INV_X1    g0670(.A(new_n680), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n347), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n873), .A2(KEYINPUT37), .A3(new_n362), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n348), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n331), .A2(new_n285), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n332), .B1(new_n328), .B2(new_n330), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n346), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n322), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n871), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(new_n880), .A3(new_n358), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n875), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n367), .B2(new_n880), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(KEYINPUT38), .B(new_n883), .C1(new_n367), .C2(new_n880), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n640), .A2(new_n643), .A3(new_n359), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n641), .A2(new_n358), .A3(new_n642), .A4(new_n872), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n889), .A2(new_n873), .B1(new_n891), .B2(new_n875), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n887), .B1(new_n892), .B2(KEYINPUT38), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n736), .B(KEYINPUT31), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n583), .A2(new_n689), .A3(new_n690), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n895), .A2(new_n676), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n744), .B1(new_n896), .B2(new_n683), .ZN(new_n897));
  NOR4_X1   g0697(.A1(new_n895), .A2(new_n676), .A3(KEYINPUT99), .A4(new_n682), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n867), .A2(new_n868), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n893), .A2(new_n899), .A3(new_n822), .A4(new_n900), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n870), .A2(new_n888), .B1(new_n901), .B2(KEYINPUT40), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n861), .A2(new_n393), .A3(new_n635), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n902), .B(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(G330), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n722), .B1(new_n748), .B2(KEYINPUT29), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT104), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(new_n907), .A3(new_n653), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n907), .B1(new_n906), .B2(new_n653), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n652), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n905), .B(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n820), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n869), .B1(new_n825), .B2(new_n913), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n914), .A2(new_n888), .B1(new_n644), .B2(new_n680), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n893), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n627), .A2(new_n682), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n886), .A2(KEYINPUT39), .A3(new_n887), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n912), .B(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n264), .B2(new_n753), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT35), .ZN(new_n924));
  AOI211_X1 g0724(.A(new_n230), .B(new_n231), .C1(new_n536), .C2(new_n924), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n925), .B(G116), .C1(new_n924), .C2(new_n536), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT36), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT103), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n334), .B2(G50), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n214), .A2(KEYINPUT103), .A3(G68), .ZN(new_n930));
  OAI21_X1  g0730(.A(G77), .B1(new_n219), .B2(new_n334), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n929), .B(new_n930), .C1(new_n229), .C2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(G1), .A3(new_n288), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n923), .A2(new_n927), .A3(new_n933), .ZN(G367));
  NAND3_X1  g0734(.A1(new_n712), .A2(KEYINPUT105), .A3(new_n682), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT105), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n544), .B2(new_n683), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n544), .B(new_n554), .C1(new_n551), .C2(new_n683), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OR3_X1    g0741(.A1(new_n941), .A2(new_n697), .A3(KEYINPUT42), .ZN(new_n942));
  OAI21_X1  g0742(.A(KEYINPUT42), .B1(new_n941), .B2(new_n697), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n712), .B1(new_n940), .B2(new_n501), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n942), .B(new_n943), .C1(new_n682), .C2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n660), .A2(new_n682), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n718), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n671), .B2(new_n946), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n945), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n696), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n940), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n950), .B(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n703), .B(KEYINPUT41), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n960));
  NAND3_X1  g0760(.A1(new_n700), .A2(new_n940), .A3(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n960), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n941), .B2(new_n699), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(KEYINPUT44), .B1(new_n700), .B2(new_n940), .ZN(new_n965));
  OR3_X1    g0765(.A1(new_n700), .A2(KEYINPUT44), .A3(new_n940), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n951), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n964), .A2(new_n696), .A3(new_n965), .A4(new_n966), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n684), .B(new_n685), .C1(new_n689), .C2(new_n682), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n697), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n694), .B2(new_n695), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n752), .A2(new_n972), .A3(new_n697), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n971), .A2(KEYINPUT107), .A3(new_n750), .A4(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT107), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n750), .A2(new_n976), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n978), .B1(new_n979), .B2(new_n970), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n959), .B1(new_n981), .B2(new_n750), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n264), .B1(new_n753), .B2(G45), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n957), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G58), .A2(new_n786), .B1(new_n837), .B2(G77), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n214), .B2(new_n791), .C1(new_n844), .C2(new_n794), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n799), .A2(new_n795), .ZN(new_n988));
  INV_X1    g0788(.A(G143), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n254), .B1(new_n781), .B2(new_n277), .C1(new_n989), .C2(new_n773), .ZN(new_n990));
  OR3_X1    g0790(.A1(new_n987), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n778), .A2(new_n334), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n778), .A2(new_n210), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n324), .B1(new_n206), .B2(new_n789), .C1(new_n841), .C2(new_n799), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(G303), .B2(new_n782), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n806), .A2(G317), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n792), .A2(G283), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n785), .A2(new_n706), .ZN(new_n998));
  INV_X1    g0798(.A(G311), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n998), .A2(KEYINPUT46), .B1(new_n999), .B2(new_n773), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(KEYINPUT46), .B2(new_n998), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n995), .A2(new_n996), .A3(new_n997), .A4(new_n1001), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n991), .A2(new_n992), .B1(new_n993), .B2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT47), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n768), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n765), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n769), .B1(new_n224), .B2(new_n384), .C1(new_n240), .C2(new_n1006), .ZN(new_n1007));
  AND3_X1   g0807(.A1(new_n1005), .A2(new_n754), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n760), .B2(new_n948), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n985), .A2(new_n1009), .ZN(G387));
  NAND3_X1  g0810(.A1(new_n749), .A2(new_n975), .A3(new_n974), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n979), .A2(new_n1011), .A3(new_n703), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n778), .A2(new_n384), .B1(new_n773), .B2(new_n795), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n789), .A2(new_n206), .B1(new_n794), .B2(new_n277), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n324), .B(new_n1014), .C1(G77), .C2(new_n786), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT109), .Z(new_n1016));
  AOI211_X1 g0816(.A(new_n1013), .B(new_n1016), .C1(G50), .C2(new_n782), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(new_n334), .B2(new_n791), .C1(new_n282), .C2(new_n799), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G322), .A2(new_n810), .B1(new_n800), .B2(G311), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n792), .A2(G303), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1019), .B(new_n1020), .C1(new_n802), .C2(new_n781), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT48), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n808), .B2(new_n778), .C1(new_n841), .C2(new_n785), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT49), .Z(new_n1024));
  NAND2_X1  g0824(.A1(new_n806), .A2(G326), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1025), .B(new_n324), .C1(new_n706), .C2(new_n789), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1018), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n768), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1028), .B(new_n754), .C1(new_n686), .C2(new_n760), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n382), .A2(new_n214), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT108), .Z(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT50), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n334), .A2(new_n216), .ZN(new_n1033));
  NOR4_X1   g0833(.A1(new_n1032), .A2(G45), .A3(new_n1033), .A4(new_n707), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1006), .B1(new_n237), .B2(G45), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n707), .B2(new_n762), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n1034), .A2(new_n1036), .B1(G107), .B2(new_n224), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1029), .B1(new_n769), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n984), .B2(new_n976), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1012), .A2(new_n1039), .ZN(G393));
  NOR2_X1   g0840(.A1(new_n970), .A2(new_n983), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n941), .A2(new_n759), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n773), .A2(new_n277), .B1(new_n781), .B2(new_n795), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT51), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n204), .B2(new_n789), .C1(new_n989), .C2(new_n794), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n382), .A2(new_n792), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n777), .A2(G77), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n324), .B1(G68), .B2(new_n786), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n800), .A2(G50), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n785), .A2(new_n808), .B1(new_n791), .B2(new_n841), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n806), .A2(G322), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(G303), .C2(new_n800), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n773), .A2(new_n802), .B1(new_n781), .B2(new_n999), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT52), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n777), .A2(G116), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1053), .A2(new_n337), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n1045), .A2(new_n1050), .B1(new_n1057), .B2(new_n790), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n768), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n769), .B1(new_n206), .B2(new_n224), .C1(new_n245), .C2(new_n1006), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n754), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT110), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1042), .A2(new_n1059), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(KEYINPUT111), .B1(new_n979), .B2(new_n970), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n977), .B2(new_n980), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n979), .A2(new_n970), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n704), .B1(new_n1067), .B2(KEYINPUT111), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1041), .B(new_n1064), .C1(new_n1066), .C2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(G390));
  INV_X1    g0870(.A(new_n919), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n889), .A2(new_n873), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n891), .A2(new_n875), .ZN(new_n1073));
  AOI21_X1  g0873(.A(KEYINPUT38), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(KEYINPUT39), .B1(new_n1075), .B2(new_n887), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n757), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n787), .B(new_n849), .C1(new_n210), .C2(new_n799), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n254), .B(new_n1078), .C1(G77), .C2(new_n777), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n810), .A2(G283), .B1(new_n806), .B2(G294), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1079), .B(new_n1080), .C1(new_n206), .C2(new_n791), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(G116), .B2(new_n782), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(KEYINPUT54), .B(G143), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n791), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n785), .A2(new_n277), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT53), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n777), .A2(G159), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n254), .B1(new_n781), .B2(new_n850), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G137), .B2(new_n800), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G50), .A2(new_n837), .B1(new_n806), .B2(G125), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1086), .A2(new_n1087), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1084), .B(new_n1091), .C1(G128), .C2(new_n810), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n768), .B1(new_n1082), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1077), .A2(new_n754), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n282), .B2(new_n832), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n899), .A2(G330), .A3(new_n822), .A4(new_n900), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n825), .A2(new_n913), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n900), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n918), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1098), .A2(new_n1099), .B1(new_n917), .B2(new_n919), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n634), .A2(new_n821), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n720), .A2(new_n683), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n869), .B1(new_n1102), .B2(new_n913), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n884), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1074), .B1(new_n1104), .B2(KEYINPUT38), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n1103), .A2(new_n1105), .A3(new_n918), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1096), .B1(new_n1100), .B2(new_n1106), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n1071), .A2(new_n1076), .B1(new_n914), .B2(new_n918), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1102), .A2(new_n913), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1099), .B(new_n893), .C1(new_n1110), .C2(new_n869), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n828), .B1(new_n897), .B2(new_n898), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1112), .A2(G330), .A3(new_n822), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1113), .A2(new_n869), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1108), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1107), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1095), .B1(new_n984), .B2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT113), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n746), .A2(new_n747), .A3(new_n823), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n900), .ZN(new_n1120));
  NOR3_X1   g0920(.A1(new_n1100), .A2(new_n1106), .A3(new_n1120), .ZN(new_n1121));
  NOR4_X1   g0921(.A1(new_n861), .A2(new_n869), .A3(new_n747), .A4(new_n823), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n861), .A2(new_n747), .A3(new_n823), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1125), .A2(new_n900), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1126), .A2(new_n1114), .A3(new_n1109), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n900), .B1(new_n829), .B2(new_n822), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1097), .B1(new_n1128), .B2(new_n1122), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(KEYINPUT112), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1096), .B1(new_n1119), .B2(new_n900), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT112), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1131), .A2(new_n1132), .A3(new_n1097), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1127), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n903), .A2(G330), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n652), .B(new_n1135), .C1(new_n909), .C2(new_n910), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1124), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1136), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1120), .B(new_n1110), .C1(new_n900), .C2(new_n1125), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1097), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1113), .A2(new_n869), .ZN(new_n1141));
  AOI211_X1 g0941(.A(KEYINPUT112), .B(new_n1140), .C1(new_n1141), .C2(new_n1096), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1132), .B1(new_n1131), .B2(new_n1097), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1139), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1138), .A2(new_n1144), .A3(new_n1116), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1137), .A2(new_n1145), .A3(new_n703), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1118), .A2(new_n1146), .ZN(G378));
  XOR2_X1   g0947(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n304), .B(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n291), .A2(new_n871), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1154), .A2(new_n757), .B1(new_n214), .B2(new_n832), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n799), .A2(new_n850), .ZN(new_n1156));
  OR3_X1    g0956(.A1(new_n785), .A2(new_n1083), .A3(KEYINPUT116), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n782), .A2(G128), .ZN(new_n1158));
  OAI21_X1  g0958(.A(KEYINPUT116), .B1(new_n785), .B2(new_n1083), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT117), .Z(new_n1161));
  AOI211_X1 g0961(.A(new_n1156), .B(new_n1161), .C1(G125), .C2(new_n810), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1162), .B1(new_n844), .B2(new_n791), .C1(new_n277), .C2(new_n778), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1163), .A2(KEYINPUT59), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n837), .A2(G159), .ZN(new_n1165));
  AOI21_X1  g0965(.A(G41), .B1(new_n806), .B2(G124), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1164), .A2(new_n252), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1163), .A2(KEYINPUT59), .ZN(new_n1168));
  AOI21_X1  g0968(.A(G41), .B1(new_n308), .B2(G33), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n1167), .A2(new_n1168), .B1(G50), .B2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n794), .A2(new_n808), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n789), .A2(new_n219), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT114), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n210), .B2(new_n781), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n992), .B(new_n1174), .C1(G97), .C2(new_n800), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n324), .B(new_n394), .C1(new_n216), .C2(new_n785), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1176), .B(KEYINPUT115), .Z(new_n1177));
  OAI211_X1 g0977(.A(new_n1175), .B(new_n1177), .C1(new_n384), .C2(new_n791), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1171), .B(new_n1178), .C1(G116), .C2(new_n810), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT58), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n768), .B1(new_n1170), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1155), .A2(new_n754), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT118), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1186));
  OAI21_X1  g0986(.A(KEYINPUT119), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1186), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT119), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1188), .A2(new_n1189), .A3(new_n1184), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1154), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n902), .B2(new_n747), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n901), .A2(KEYINPUT40), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n861), .A2(new_n823), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT40), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1195), .A2(new_n1196), .A3(new_n888), .A4(new_n900), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1194), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1198), .A2(G330), .A3(new_n1154), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1193), .A2(new_n921), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n921), .B1(new_n1193), .B2(new_n1199), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n984), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1191), .A2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1138), .B1(new_n1134), .B2(new_n1124), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(KEYINPUT120), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT120), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1138), .B(new_n1207), .C1(new_n1134), .C2(new_n1124), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1206), .A2(new_n1202), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT57), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n704), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1206), .A2(KEYINPUT57), .A3(new_n1202), .A4(new_n1208), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1204), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(G375));
  NAND2_X1  g1014(.A1(new_n832), .A2(new_n334), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n900), .A2(new_n758), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n786), .A2(G159), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n324), .B1(G128), .B2(new_n806), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n792), .A2(G150), .B1(new_n777), .B2(G50), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1173), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT121), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1083), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G137), .A2(new_n782), .B1(new_n800), .B2(new_n1222), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1221), .B(new_n1223), .C1(new_n850), .C2(new_n773), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n778), .A2(new_n384), .B1(new_n773), .B2(new_n841), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n806), .A2(G303), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n216), .A2(new_n789), .B1(new_n791), .B2(new_n210), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n337), .B1(new_n785), .B2(new_n206), .ZN(new_n1228));
  NOR4_X1   g1028(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1229), .B1(new_n706), .B2(new_n799), .C1(new_n808), .C2(new_n781), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n857), .B1(new_n1224), .B2(new_n1230), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1216), .A2(new_n755), .A3(new_n1231), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1144), .A2(new_n984), .B1(new_n1215), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n958), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1138), .A2(new_n1144), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1233), .B1(new_n1235), .B2(new_n1237), .ZN(G381));
  INV_X1    g1038(.A(G384), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1146), .A2(new_n1117), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(KEYINPUT122), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT122), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1146), .A2(new_n1242), .A3(new_n1117), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1241), .A2(new_n1243), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n985), .A2(new_n1069), .A3(new_n1009), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1213), .A2(new_n1239), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(G393), .A2(G396), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1233), .B(new_n1247), .C1(new_n1235), .C2(new_n1237), .ZN(new_n1248));
  OAI21_X1  g1048(.A(KEYINPUT123), .B1(new_n1246), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1250), .A2(new_n703), .A3(new_n1212), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1204), .ZN(new_n1252));
  AND4_X1   g1052(.A1(new_n1251), .A2(new_n1252), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT123), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1248), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1239), .A4(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1249), .A2(new_n1256), .ZN(G407));
  INV_X1    g1057(.A(G213), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1244), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(G375), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1258), .B1(new_n1260), .B2(new_n681), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G407), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT124), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(G407), .A2(KEYINPUT124), .A3(new_n1261), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(G409));
  XOR2_X1   g1066(.A(G393), .B(G396), .Z(new_n1267));
  AOI21_X1  g1067(.A(new_n1069), .B1(new_n985), .B2(new_n1009), .ZN(new_n1268));
  OAI21_X1  g1068(.A(KEYINPUT127), .B1(new_n1245), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(G387), .A2(G390), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT127), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n985), .A2(new_n1069), .A3(new_n1009), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1267), .B1(new_n1269), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1267), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1275), .B1(new_n1276), .B2(KEYINPUT127), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1274), .A2(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1258), .A2(G343), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT60), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1234), .A2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1134), .A2(KEYINPUT60), .A3(new_n1136), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1281), .A2(new_n1236), .A3(new_n703), .A4(new_n1282), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1283), .A2(G384), .A3(new_n1233), .ZN(new_n1284));
  AOI21_X1  g1084(.A(G384), .B1(new_n1283), .B2(new_n1233), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G2897), .B(new_n1279), .C1(new_n1284), .C2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1285), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1283), .A2(G384), .A3(new_n1233), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1279), .A2(G2897), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1287), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1286), .A2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1136), .B1(new_n1144), .B2(new_n1116), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1292), .A2(new_n1207), .ZN(new_n1293));
  AOI211_X1 g1093(.A(KEYINPUT120), .B(new_n1136), .C1(new_n1144), .C2(new_n1116), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT125), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1295), .A2(new_n1296), .A3(new_n958), .A4(new_n1202), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n983), .B1(new_n1202), .B2(KEYINPUT126), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT126), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1300));
  AOI22_X1  g1100(.A1(new_n1298), .A2(new_n1300), .B1(new_n1184), .B2(new_n1188), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1206), .A2(new_n958), .A3(new_n1202), .A4(new_n1208), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(KEYINPUT125), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1297), .A2(new_n1301), .A3(new_n1303), .ZN(new_n1304));
  AOI22_X1  g1104(.A1(G378), .A2(new_n1213), .B1(new_n1304), .B2(new_n1244), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1291), .B1(new_n1305), .B2(new_n1279), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1304), .A2(new_n1244), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1251), .A2(G378), .A3(new_n1252), .ZN(new_n1309));
  AOI211_X1 g1109(.A(new_n1279), .B(new_n1307), .C1(new_n1308), .C2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT62), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1306), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1279), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1307), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1313), .A2(new_n1311), .A3(new_n1314), .A4(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT61), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1278), .B1(new_n1312), .B2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1313), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1286), .A2(new_n1290), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1321), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT63), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1320), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1278), .A2(KEYINPUT61), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1310), .A2(KEYINPUT63), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1324), .A2(new_n1325), .A3(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1319), .A2(new_n1327), .ZN(G405));
  OAI21_X1  g1128(.A(new_n1309), .B1(new_n1213), .B2(new_n1259), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n1315), .ZN(new_n1330));
  OAI211_X1 g1130(.A(new_n1309), .B(new_n1307), .C1(new_n1213), .C2(new_n1259), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(new_n1332), .B(new_n1278), .ZN(G402));
endmodule


