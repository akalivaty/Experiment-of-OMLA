//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(KEYINPUT64), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT64), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n215), .A2(G1), .A3(G13), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G20), .ZN(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n212), .B1(new_n218), .B2(new_n219), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT65), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G274), .ZN(new_n248));
  AND2_X1   g0048(.A1(G1), .A2(G13), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G41), .A2(G45), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G1), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(KEYINPUT66), .B1(new_n252), .B2(G1), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT66), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n256), .B(new_n257), .C1(G41), .C2(G45), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n250), .A2(G1), .A3(G13), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n255), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n254), .B1(new_n260), .B2(new_n222), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G33), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n264), .A2(new_n266), .A3(G232), .A4(G1698), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  NAND4_X1  g0068(.A1(new_n264), .A2(new_n266), .A3(G226), .A4(new_n268), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n267), .B(new_n269), .C1(new_n263), .C2(new_n205), .ZN(new_n270));
  AND2_X1   g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n271), .B1(new_n214), .B2(new_n216), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n262), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT13), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT13), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n262), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT75), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(new_n279), .A3(G169), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT14), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT14), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n278), .A2(new_n279), .A3(new_n282), .A4(G169), .ZN(new_n283));
  INV_X1    g0083(.A(G179), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n281), .B(new_n283), .C1(new_n284), .C2(new_n278), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n257), .A2(G20), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n214), .A2(new_n216), .A3(new_n287), .A4(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT69), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n289), .A2(new_n290), .ZN(new_n292));
  OAI211_X1 g0092(.A(G68), .B(new_n286), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n287), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n221), .ZN(new_n295));
  AND2_X1   g0095(.A1(KEYINPUT71), .A2(KEYINPUT12), .ZN(new_n296));
  NOR2_X1   g0096(.A1(KEYINPUT71), .A2(KEYINPUT12), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(new_n295), .B2(new_n297), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n214), .A2(new_n216), .A3(new_n288), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT67), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n214), .A2(new_n216), .A3(KEYINPUT67), .A4(new_n288), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT11), .ZN(new_n305));
  NOR2_X1   g0105(.A1(G20), .A2(G33), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n306), .A2(G50), .B1(G20), .B2(new_n221), .ZN(new_n307));
  INV_X1    g0107(.A(G77), .ZN(new_n308));
  INV_X1    g0108(.A(G20), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G33), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n307), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n304), .A2(new_n305), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n305), .B1(new_n304), .B2(new_n311), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n293), .B(new_n299), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT72), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n304), .A2(new_n311), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT11), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n304), .A2(new_n305), .A3(new_n311), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT72), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n319), .A2(new_n320), .A3(new_n293), .A4(new_n299), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n315), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n285), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G244), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n254), .B1(new_n260), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g0126(.A(KEYINPUT3), .B(G33), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n327), .A2(G232), .A3(new_n268), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(G1698), .ZN(new_n329));
  OAI221_X1 g0129(.A(new_n328), .B1(new_n206), .B2(new_n327), .C1(new_n329), .C2(new_n222), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n326), .B1(new_n330), .B2(new_n272), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G200), .ZN(new_n333));
  OAI211_X1 g0133(.A(G77), .B(new_n286), .C1(new_n291), .C2(new_n292), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT8), .B(G58), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n336), .A2(new_n306), .B1(G20), .B2(G77), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT15), .B(G87), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n310), .B2(new_n338), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n339), .A2(new_n300), .B1(new_n308), .B2(new_n294), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n331), .A2(G190), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n333), .A2(new_n334), .A3(new_n340), .A4(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n327), .A2(G222), .A3(new_n268), .ZN(new_n343));
  INV_X1    g0143(.A(G223), .ZN(new_n344));
  OAI221_X1 g0144(.A(new_n343), .B1(new_n308), .B2(new_n327), .C1(new_n329), .C2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n272), .ZN(new_n346));
  INV_X1    g0146(.A(new_n260), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n347), .A2(G226), .B1(new_n253), .B2(new_n251), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G169), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n304), .A2(new_n294), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n286), .A2(G50), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n353), .B(KEYINPUT68), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n203), .A2(G20), .ZN(new_n356));
  INV_X1    g0156(.A(G150), .ZN(new_n357));
  INV_X1    g0157(.A(new_n306), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n356), .B1(new_n357), .B2(new_n358), .C1(new_n310), .C2(new_n335), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n359), .A2(new_n304), .B1(new_n202), .B2(new_n294), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n351), .B(new_n361), .C1(G179), .C2(new_n349), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n332), .A2(new_n350), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n340), .A2(new_n334), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n331), .A2(new_n284), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n342), .A2(new_n362), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G200), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n346), .B2(new_n348), .ZN(new_n369));
  INV_X1    g0169(.A(new_n349), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n369), .B1(new_n370), .B2(G190), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n361), .A2(KEYINPUT9), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT9), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(new_n355), .B2(new_n360), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT70), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT10), .B1(new_n369), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NOR3_X1   g0179(.A1(new_n372), .A2(new_n376), .A3(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n379), .B1(new_n372), .B2(new_n376), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n324), .B(new_n367), .C1(new_n380), .C2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT74), .ZN(new_n384));
  INV_X1    g0184(.A(new_n277), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n276), .B1(new_n262), .B2(new_n273), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n368), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G190), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n275), .A2(new_n388), .A3(new_n277), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT73), .ZN(new_n391));
  AND3_X1   g0191(.A1(new_n322), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n391), .B1(new_n322), .B2(new_n390), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n384), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n322), .A2(new_n390), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT73), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n322), .A2(new_n390), .A3(new_n391), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(KEYINPUT74), .A3(new_n397), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n335), .B1(new_n257), .B2(G20), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n352), .A2(new_n400), .B1(new_n294), .B2(new_n335), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT76), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT7), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n327), .B2(G20), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n264), .A2(new_n266), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(KEYINPUT7), .A3(new_n309), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n221), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G58), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n409), .A2(new_n221), .ZN(new_n410));
  OAI21_X1  g0210(.A(G20), .B1(new_n410), .B2(new_n201), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n306), .A2(G159), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n402), .B(new_n403), .C1(new_n408), .C2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(KEYINPUT7), .B1(new_n406), .B2(new_n309), .ZN(new_n415));
  AOI211_X1 g0215(.A(new_n404), .B(G20), .C1(new_n264), .C2(new_n266), .ZN(new_n416));
  OAI21_X1  g0216(.A(G68), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n413), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(KEYINPUT16), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n414), .A2(new_n419), .A3(new_n300), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n417), .A2(new_n418), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n402), .B1(new_n421), .B2(new_n403), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n401), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT77), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n403), .B1(new_n408), .B2(new_n413), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT76), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n426), .A2(new_n300), .A3(new_n414), .A4(new_n419), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT77), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(new_n428), .A3(new_n401), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n255), .A2(G232), .A3(new_n258), .A4(new_n259), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n254), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT78), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n430), .A2(KEYINPUT78), .A3(new_n254), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n264), .A2(new_n266), .A3(G226), .A4(G1698), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n264), .A2(new_n266), .A3(G223), .A4(new_n268), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n435), .B(new_n436), .C1(new_n263), .C2(new_n223), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n272), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n433), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G169), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n284), .B2(new_n439), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n424), .A2(new_n429), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT18), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT17), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n431), .A2(new_n432), .B1(new_n437), .B2(new_n272), .ZN(new_n445));
  AOI21_X1  g0245(.A(G200), .B1(new_n445), .B2(new_n434), .ZN(new_n446));
  AND4_X1   g0246(.A1(new_n388), .A2(new_n433), .A3(new_n434), .A4(new_n438), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n444), .B1(new_n423), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n439), .A2(new_n368), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(G190), .B2(new_n439), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n451), .A2(new_n427), .A3(KEYINPUT17), .A4(new_n401), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT18), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n424), .A2(new_n429), .A3(new_n454), .A4(new_n441), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n443), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n383), .A2(new_n399), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(G45), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(G1), .ZN(new_n460));
  NAND2_X1  g0260(.A1(KEYINPUT5), .A2(G41), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(G274), .B1(new_n271), .B2(new_n213), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT80), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n257), .A2(G45), .ZN(new_n467));
  OR2_X1    g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n467), .B1(new_n468), .B2(new_n461), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT80), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(new_n251), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT5), .B(G41), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n472), .A2(new_n460), .B1(new_n249), .B2(new_n250), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n466), .A2(new_n471), .B1(new_n473), .B2(G257), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n264), .A2(new_n266), .A3(G244), .A4(new_n268), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT4), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G283), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n263), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G250), .A2(G1698), .ZN(new_n480));
  NAND2_X1  g0280(.A1(KEYINPUT4), .A2(G244), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n480), .B1(new_n481), .B2(G1698), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n479), .B1(new_n327), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n272), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n474), .A2(new_n485), .A3(KEYINPUT81), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT81), .B1(new_n474), .B2(new_n485), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n350), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n474), .A2(new_n485), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(G179), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT6), .ZN(new_n492));
  XNOR2_X1  g0292(.A(G97), .B(G107), .ZN(new_n493));
  XNOR2_X1  g0293(.A(KEYINPUT79), .B(G97), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n492), .A2(G107), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n492), .A2(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI22_X1  g0296(.A1(new_n496), .A2(new_n309), .B1(new_n308), .B2(new_n358), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n206), .B1(new_n405), .B2(new_n407), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n300), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n257), .A2(G33), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n302), .A2(new_n287), .A3(new_n303), .A4(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G97), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n499), .B(new_n503), .C1(G97), .C2(new_n287), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n488), .A2(new_n491), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT81), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n464), .A2(G257), .A3(new_n259), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT80), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n470), .B1(new_n469), .B2(new_n251), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n272), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(new_n477), .B2(new_n483), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n506), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n474), .A2(new_n485), .A3(KEYINPUT81), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(G190), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT82), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n513), .A2(KEYINPUT82), .A3(G190), .A4(new_n514), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n504), .B1(G200), .B2(new_n489), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT83), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT83), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n519), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n505), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n327), .A2(new_n309), .A3(G68), .ZN(new_n526));
  NOR2_X1   g0326(.A1(KEYINPUT79), .A2(G97), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(KEYINPUT79), .A2(G97), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n310), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n526), .B1(new_n530), .B2(KEYINPUT19), .ZN(new_n531));
  INV_X1    g0331(.A(new_n494), .ZN(new_n532));
  NOR2_X1   g0332(.A1(G87), .A2(G107), .ZN(new_n533));
  NAND3_X1  g0333(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n532), .A2(new_n533), .B1(new_n309), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n300), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n338), .A2(new_n294), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n502), .A2(G87), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n264), .A2(new_n266), .A3(G244), .A4(G1698), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n264), .A2(new_n266), .A3(G238), .A4(new_n268), .ZN(new_n541));
  XNOR2_X1  g0341(.A(KEYINPUT84), .B(G116), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n540), .B(new_n541), .C1(new_n263), .C2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n272), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n460), .A2(new_n248), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n467), .A2(new_n224), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n259), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G200), .ZN(new_n549));
  INV_X1    g0349(.A(new_n547), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(new_n543), .B2(new_n272), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G190), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n538), .A2(new_n539), .A3(new_n549), .A4(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n548), .A2(new_n350), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n551), .A2(new_n284), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n536), .A2(new_n537), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n501), .A2(new_n338), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n554), .B(new_n555), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n525), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(G116), .B(new_n500), .C1(new_n291), .C2(new_n292), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n542), .A2(new_n294), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n542), .A2(G20), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n300), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n309), .B1(new_n263), .B2(new_n478), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n566), .B1(new_n494), .B2(new_n263), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n568), .A2(KEYINPUT20), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT20), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n565), .A2(new_n570), .A3(new_n567), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n562), .B(new_n563), .C1(new_n569), .C2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n265), .A2(G33), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n574));
  OAI21_X1  g0374(.A(G303), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n264), .A2(new_n266), .A3(G264), .A4(G1698), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n264), .A2(new_n266), .A3(G257), .A4(new_n268), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n272), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n466), .A2(new_n471), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n473), .A2(G270), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n582), .A2(G169), .ZN(new_n583));
  AOI21_X1  g0383(.A(KEYINPUT21), .B1(new_n572), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n582), .A2(G200), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n388), .B2(new_n582), .ZN(new_n587));
  OR2_X1    g0387(.A1(new_n587), .A2(new_n572), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n582), .A2(KEYINPUT21), .A3(G169), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n579), .A2(new_n580), .A3(G179), .A4(new_n581), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT85), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n591), .A2(new_n592), .A3(new_n572), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n592), .B1(new_n591), .B2(new_n572), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n585), .B(new_n588), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n473), .A2(G264), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n224), .A2(new_n268), .ZN(new_n597));
  INV_X1    g0397(.A(G257), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G1698), .ZN(new_n599));
  AND4_X1   g0399(.A1(new_n264), .A2(new_n597), .A3(new_n266), .A4(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(G294), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT86), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT86), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G294), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n263), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n272), .B1(new_n600), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n580), .A2(new_n596), .A3(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT87), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(new_n608), .A3(G169), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n580), .A2(new_n606), .A3(G179), .A4(new_n596), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n608), .B1(new_n607), .B2(G169), .ZN(new_n612));
  OAI21_X1  g0412(.A(KEYINPUT88), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n327), .A2(new_n309), .A3(G87), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT22), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT22), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n327), .A2(new_n616), .A3(new_n309), .A4(G87), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT24), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n542), .A2(new_n263), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT23), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n309), .B2(G107), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n620), .A2(new_n309), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n618), .A2(new_n619), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n619), .B1(new_n618), .B2(new_n624), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n300), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n294), .A2(new_n206), .ZN(new_n628));
  XNOR2_X1  g0428(.A(new_n628), .B(KEYINPUT25), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n502), .B2(G107), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n607), .A2(G169), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT87), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT88), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n633), .A2(new_n634), .A3(new_n610), .A4(new_n609), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n613), .A2(new_n631), .A3(new_n635), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n607), .A2(new_n388), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n607), .A2(G200), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n627), .A2(new_n630), .A3(new_n637), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NOR4_X1   g0440(.A1(new_n458), .A2(new_n561), .A3(new_n595), .A4(new_n640), .ZN(G372));
  INV_X1    g0441(.A(new_n362), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n423), .A2(new_n441), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT18), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n423), .A2(new_n454), .A3(new_n441), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n396), .A2(new_n397), .ZN(new_n648));
  INV_X1    g0448(.A(new_n366), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n648), .A2(new_n649), .B1(new_n323), .B2(new_n285), .ZN(new_n650));
  INV_X1    g0450(.A(new_n453), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n647), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n380), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n653), .A2(KEYINPUT90), .A3(new_n381), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT90), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n382), .B2(new_n380), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n642), .B1(new_n652), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n558), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n493), .A2(new_n492), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n494), .A2(new_n495), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n662), .A2(G20), .B1(G77), .B2(new_n306), .ZN(new_n663));
  OAI21_X1  g0463(.A(G107), .B1(new_n415), .B2(new_n416), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n665), .A2(new_n300), .B1(new_n205), .B2(new_n294), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n490), .B1(new_n666), .B2(new_n503), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n667), .A2(new_n558), .A3(new_n553), .A4(new_n488), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n659), .B1(new_n668), .B2(KEYINPUT26), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT89), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n559), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT26), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n553), .A2(new_n558), .A3(KEYINPUT89), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n671), .A2(new_n505), .A3(new_n672), .A4(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n631), .B1(new_n612), .B2(new_n611), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n591), .A2(new_n572), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n676), .A2(new_n585), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n671), .A2(new_n639), .A3(new_n673), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n675), .B1(new_n525), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n658), .B1(new_n458), .B2(new_n681), .ZN(G369));
  NAND2_X1  g0482(.A1(new_n585), .A2(new_n677), .ZN(new_n683));
  INV_X1    g0483(.A(new_n595), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n257), .A2(new_n309), .A3(G13), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n687));
  INV_X1    g0487(.A(G213), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G343), .ZN(new_n690));
  XOR2_X1   g0490(.A(new_n690), .B(KEYINPUT91), .Z(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n572), .ZN(new_n693));
  MUX2_X1   g0493(.A(new_n683), .B(new_n684), .S(new_n693), .Z(new_n694));
  AND2_X1   g0494(.A1(new_n694), .A2(G330), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n691), .B1(new_n627), .B2(new_n630), .ZN(new_n696));
  OAI22_X1  g0496(.A1(new_n640), .A2(new_n696), .B1(new_n636), .B2(new_n691), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n593), .A2(new_n594), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n584), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(new_n692), .ZN(new_n701));
  INV_X1    g0501(.A(new_n640), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n676), .A2(new_n692), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n698), .A2(new_n705), .ZN(G399));
  INV_X1    g0506(.A(new_n210), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(G1), .ZN(new_n710));
  INV_X1    g0510(.A(G116), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n532), .A2(new_n711), .A3(new_n533), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n710), .A2(new_n712), .B1(new_n219), .B2(new_n709), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  INV_X1    g0514(.A(G330), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n636), .A2(new_n639), .A3(new_n691), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n595), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n522), .A2(new_n524), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n667), .A2(new_n488), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n717), .A2(new_n718), .A3(new_n560), .A4(new_n719), .ZN(new_n720));
  AND4_X1   g0520(.A1(G179), .A2(new_n579), .A3(new_n580), .A4(new_n581), .ZN(new_n721));
  AND4_X1   g0521(.A1(new_n544), .A2(new_n547), .A3(new_n596), .A4(new_n606), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n513), .A2(new_n721), .A3(new_n722), .A4(new_n514), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT93), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n582), .A2(new_n548), .A3(new_n284), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT92), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n582), .A2(new_n548), .A3(KEYINPUT92), .A4(new_n284), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n729), .A2(new_n489), .A3(new_n607), .A4(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n486), .A2(new_n487), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT93), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n551), .A2(new_n596), .A3(new_n606), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(new_n590), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n732), .A2(new_n733), .A3(KEYINPUT30), .A4(new_n735), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n725), .A2(new_n726), .A3(new_n731), .A4(new_n736), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n737), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n738));
  AOI21_X1  g0538(.A(KEYINPUT31), .B1(new_n737), .B2(new_n692), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n715), .B1(new_n720), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n681), .A2(new_n692), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n742), .A2(KEYINPUT29), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n679), .B1(new_n700), .B2(new_n636), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n744), .A2(new_n525), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n671), .A2(new_n673), .ZN(new_n746));
  OAI21_X1  g0546(.A(KEYINPUT26), .B1(new_n746), .B2(new_n719), .ZN(new_n747));
  INV_X1    g0547(.A(new_n668), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n659), .B1(new_n748), .B2(new_n672), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  OAI211_X1 g0550(.A(KEYINPUT29), .B(new_n691), .C1(new_n745), .C2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n741), .B1(new_n743), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n714), .B1(new_n752), .B2(G1), .ZN(G364));
  OR2_X1    g0553(.A1(new_n694), .A2(G330), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT94), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n309), .A2(G13), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n257), .B1(new_n756), .B2(G45), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n708), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n695), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n759), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n309), .B1(KEYINPUT97), .B2(new_n350), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(KEYINPUT97), .B2(new_n350), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n764), .A2(new_n217), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT98), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(KEYINPUT98), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n388), .A2(G179), .A3(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n309), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n205), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n309), .A2(new_n284), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n388), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n309), .A2(G179), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(new_n388), .A3(G200), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n776), .A2(new_n202), .B1(new_n778), .B2(new_n206), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n777), .A2(G190), .A3(G200), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n772), .B(new_n779), .C1(G87), .C2(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n773), .A2(new_n388), .A3(G200), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n783), .A2(KEYINPUT99), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(KEYINPUT99), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G68), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G190), .A2(G200), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n777), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G159), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT32), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n773), .A2(G190), .A3(new_n368), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n327), .B1(new_n794), .B2(new_n409), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n773), .A2(new_n789), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n795), .B1(G77), .B2(new_n797), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n782), .A2(new_n788), .A3(new_n793), .A4(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G322), .ZN(new_n800));
  INV_X1    g0600(.A(G311), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n794), .A2(new_n800), .B1(new_n796), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n790), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n327), .B(new_n802), .C1(G329), .C2(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(KEYINPUT100), .B(KEYINPUT33), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(G317), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n787), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n771), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n602), .A2(new_n604), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n808), .A2(new_n809), .B1(new_n781), .B2(G303), .ZN(new_n810));
  INV_X1    g0610(.A(new_n778), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n775), .A2(G326), .B1(new_n811), .B2(G283), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n804), .A2(new_n807), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n769), .B1(new_n799), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(G13), .A2(G33), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT96), .Z(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(G20), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n768), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n707), .A2(new_n406), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT95), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n820), .A2(G355), .B1(new_n711), .B2(new_n707), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n246), .A2(G45), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n707), .A2(new_n327), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(G45), .B2(new_n219), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n821), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n762), .B(new_n814), .C1(new_n818), .C2(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n817), .B(KEYINPUT101), .Z(new_n827));
  OAI21_X1  g0627(.A(new_n826), .B1(new_n694), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n761), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(G396));
  NAND2_X1  g0630(.A1(new_n692), .A2(new_n364), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n831), .A2(new_n366), .A3(new_n342), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(KEYINPUT103), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT103), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n831), .A2(new_n834), .A3(new_n342), .A4(new_n366), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n649), .A2(new_n692), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n833), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n833), .A2(new_n835), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n691), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n742), .A2(new_n837), .B1(new_n681), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n741), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n759), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n841), .B2(new_n840), .ZN(new_n843));
  INV_X1    g0643(.A(new_n794), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n844), .A2(G143), .B1(new_n797), .B2(G159), .ZN(new_n845));
  INV_X1    g0645(.A(G137), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n845), .B1(new_n846), .B2(new_n776), .C1(new_n786), .C2(new_n357), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n848), .A2(KEYINPUT34), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(KEYINPUT34), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n778), .A2(new_n221), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n406), .B1(new_n803), .B2(G132), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n202), .B2(new_n780), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n851), .B(new_n853), .C1(G58), .C2(new_n808), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n849), .A2(new_n850), .A3(new_n854), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n223), .A2(new_n778), .B1(new_n780), .B2(new_n206), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n772), .B(new_n856), .C1(G303), .C2(new_n775), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n794), .A2(new_n601), .B1(new_n796), .B2(new_n542), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n327), .B(new_n858), .C1(G311), .C2(new_n803), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n857), .B(new_n859), .C1(new_n478), .C2(new_n786), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n769), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n769), .A2(new_n816), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT102), .Z(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n762), .B(new_n861), .C1(new_n308), .C2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n837), .B2(new_n816), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n843), .A2(new_n866), .ZN(G384));
  AOI211_X1 g0667(.A(new_n711), .B(new_n218), .C1(new_n662), .C2(KEYINPUT35), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(KEYINPUT35), .B2(new_n662), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT36), .Z(new_n870));
  OR3_X1    g0670(.A1(new_n410), .A2(new_n219), .A3(new_n308), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n202), .A2(G68), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n257), .B(G13), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n644), .A2(new_n449), .A3(new_n452), .A4(new_n645), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n424), .A2(new_n429), .A3(new_n689), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT104), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n451), .A2(new_n427), .A3(new_n401), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n643), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT37), .B1(new_n876), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n424), .A2(new_n429), .A3(new_n689), .ZN(new_n883));
  INV_X1    g0683(.A(new_n423), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT37), .B1(new_n884), .B2(new_n451), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n442), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n875), .A2(KEYINPUT104), .A3(new_n876), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n879), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n419), .A2(new_n425), .A3(new_n304), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n401), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n689), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n456), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n441), .A2(new_n893), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n880), .A2(new_n897), .A3(new_n894), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT37), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n886), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n896), .A2(KEYINPUT38), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT39), .B1(new_n891), .B2(new_n901), .ZN(new_n902));
  AOI221_X4 g0702(.A(new_n890), .B1(new_n886), .B2(new_n899), .C1(new_n456), .C2(new_n895), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT38), .B1(new_n896), .B2(new_n900), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT39), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NOR4_X1   g0706(.A1(new_n902), .A2(new_n906), .A3(new_n324), .A4(new_n692), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n366), .A2(new_n692), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n681), .B2(new_n839), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n323), .A2(new_n692), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n324), .A2(new_n648), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n285), .B1(new_n394), .B2(new_n398), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n912), .B1(new_n913), .B2(new_n911), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n910), .B(new_n914), .C1(new_n903), .C2(new_n904), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n647), .B2(new_n689), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n907), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n751), .B(new_n457), .C1(KEYINPUT29), .C2(new_n742), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n658), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n917), .B(new_n919), .Z(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT105), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n878), .A2(new_n877), .B1(new_n882), .B2(new_n886), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT38), .B1(new_n923), .B2(new_n888), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n922), .B1(new_n924), .B2(new_n903), .ZN(new_n925));
  INV_X1    g0725(.A(new_n837), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n720), .B2(new_n740), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n927), .A2(new_n914), .A3(KEYINPUT40), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n891), .A2(KEYINPUT105), .A3(new_n901), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n925), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n927), .B(new_n914), .C1(new_n903), .C2(new_n904), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT40), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n720), .A2(new_n740), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n457), .A2(new_n935), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n934), .A2(new_n936), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n937), .A2(new_n938), .A3(new_n715), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n921), .A2(new_n939), .B1(new_n257), .B2(new_n756), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n921), .A2(new_n939), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n874), .B1(new_n940), .B2(new_n941), .ZN(G367));
  NAND2_X1  g0742(.A1(new_n692), .A2(new_n504), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n525), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n505), .A2(new_n692), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n946), .A2(new_n702), .A3(new_n701), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n947), .A2(KEYINPUT42), .ZN(new_n948));
  INV_X1    g0748(.A(new_n636), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n718), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n692), .B1(new_n950), .B2(new_n719), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n947), .B2(KEYINPUT42), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n691), .B1(new_n538), .B2(new_n539), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT106), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n954), .A2(new_n746), .ZN(new_n955));
  AOI211_X1 g0755(.A(KEYINPUT107), .B(new_n955), .C1(new_n659), .C2(new_n954), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n954), .A2(new_n659), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n956), .B1(KEYINPUT107), .B2(new_n957), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n948), .A2(new_n952), .B1(new_n958), .B2(KEYINPUT43), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n695), .A2(new_n697), .A3(new_n946), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n961), .B(new_n962), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n708), .B(KEYINPUT41), .Z(new_n964));
  INV_X1    g0764(.A(KEYINPUT108), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n965), .A2(KEYINPUT44), .ZN(new_n966));
  NOR3_X1   g0766(.A1(new_n705), .A2(new_n946), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(KEYINPUT44), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n967), .B(new_n968), .Z(new_n969));
  NAND2_X1  g0769(.A1(new_n705), .A2(new_n946), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT45), .Z(new_n971));
  AOI21_X1  g0771(.A(new_n698), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n703), .B1(new_n697), .B2(new_n701), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n695), .B(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n752), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n969), .A2(new_n971), .A3(new_n698), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n973), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n964), .B1(new_n979), .B2(new_n752), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n963), .B1(new_n980), .B2(new_n758), .ZN(new_n981));
  INV_X1    g0781(.A(new_n338), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n817), .B(new_n768), .C1(new_n707), .C2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n823), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n235), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n762), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n787), .A2(G159), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n796), .A2(new_n202), .B1(new_n790), .B2(new_n846), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n406), .B(new_n988), .C1(G150), .C2(new_n844), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n771), .A2(new_n221), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G77), .B2(new_n811), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n775), .A2(G143), .B1(new_n781), .B2(G58), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n987), .A2(new_n989), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n808), .A2(G107), .B1(new_n811), .B2(new_n494), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n844), .A2(G303), .B1(new_n797), .B2(G283), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n327), .B1(new_n803), .B2(G317), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n775), .A2(G311), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n994), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(KEYINPUT46), .B1(new_n780), .B2(new_n711), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n542), .A2(KEYINPUT46), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n999), .B1(new_n1000), .B2(new_n780), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n809), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1001), .B1(new_n786), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n993), .B1(new_n998), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT47), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n768), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n986), .B1(new_n1006), .B2(new_n1007), .C1(new_n958), .C2(new_n827), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n981), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1009), .A2(KEYINPUT109), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT109), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(new_n981), .B2(new_n1008), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(G387));
  AND2_X1   g0814(.A1(new_n975), .A2(new_n758), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1015), .A2(KEYINPUT110), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(KEYINPUT110), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n697), .A2(new_n827), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n844), .A2(G317), .B1(new_n797), .B2(G303), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n800), .B2(new_n776), .C1(new_n786), .C2(new_n801), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT48), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n808), .A2(G283), .B1(new_n781), .B2(new_n809), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n542), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n811), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n327), .B1(new_n803), .B2(G326), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1027), .A2(new_n1028), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n794), .A2(new_n202), .B1(new_n790), .B2(new_n357), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n406), .B(new_n1033), .C1(G68), .C2(new_n797), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n787), .A2(new_n336), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n808), .A2(new_n982), .B1(new_n811), .B2(G97), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n775), .A2(G159), .B1(new_n781), .B2(G77), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n769), .B1(new_n1032), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n820), .A2(new_n712), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(G107), .B2(new_n210), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT111), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AOI211_X1 g0843(.A(G45), .B(new_n712), .C1(G68), .C2(G77), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n335), .A2(G50), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT50), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n984), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n459), .B2(new_n239), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1043), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n762), .B(new_n1039), .C1(new_n818), .C2(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1016), .A2(new_n1017), .B1(new_n1018), .B2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n977), .A2(new_n709), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n752), .B2(new_n975), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1054), .ZN(G393));
  INV_X1    g0855(.A(new_n978), .ZN(new_n1056));
  NOR3_X1   g0856(.A1(new_n1056), .A2(new_n757), .A3(new_n972), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n944), .A2(new_n817), .A3(new_n945), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n243), .A2(new_n823), .B1(new_n707), .B2(new_n494), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n818), .A2(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G317), .A2(new_n775), .B1(new_n844), .B2(G311), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT52), .Z(new_n1062));
  NAND2_X1  g0862(.A1(new_n787), .A2(G303), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n406), .B1(new_n790), .B2(new_n800), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G294), .B2(new_n797), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n206), .A2(new_n778), .B1(new_n780), .B2(new_n478), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n1029), .B2(new_n808), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1062), .A2(new_n1063), .A3(new_n1065), .A4(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n776), .A2(new_n357), .B1(new_n791), .B2(new_n794), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT51), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n778), .A2(new_n223), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n406), .B(new_n1071), .C1(G143), .C2(new_n803), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n771), .A2(new_n308), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(G68), .B2(new_n781), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1070), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n786), .A2(new_n202), .B1(new_n335), .B2(new_n796), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT113), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1068), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n762), .B(new_n1060), .C1(new_n1078), .C2(new_n768), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1057), .B1(new_n1058), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n976), .B1(new_n1056), .B2(new_n972), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1081), .A2(new_n979), .A3(new_n708), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1082), .ZN(G390));
  NOR2_X1   g0883(.A1(new_n324), .A2(new_n692), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n750), .B1(new_n525), .B2(new_n744), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n909), .B1(new_n1085), .B2(new_n839), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1084), .B1(new_n1086), .B2(new_n914), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1087), .A2(new_n925), .A3(new_n929), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1084), .B1(new_n910), .B2(new_n914), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT114), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n902), .A2(new_n906), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1088), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n741), .A2(new_n837), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n914), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1096), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1088), .B(new_n1098), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1100), .A2(new_n757), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(KEYINPUT54), .B(G143), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n844), .A2(G132), .B1(new_n797), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(G128), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1104), .B1(new_n1105), .B2(new_n776), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G159), .B2(new_n808), .ZN(new_n1107));
  INV_X1    g0907(.A(G125), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n327), .B1(new_n790), .B2(new_n1108), .C1(new_n202), .C2(new_n778), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT115), .Z(new_n1110));
  NAND2_X1  g0910(.A1(new_n787), .A2(G137), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n780), .A2(new_n357), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT53), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1107), .A2(new_n1110), .A3(new_n1111), .A4(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n406), .B1(new_n780), .B2(new_n223), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n787), .A2(G107), .B1(KEYINPUT116), .B2(new_n1115), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n794), .A2(new_n711), .B1(new_n790), .B2(new_n601), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n494), .B2(new_n797), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n851), .B(new_n1073), .C1(G283), .C2(new_n775), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n1115), .A2(KEYINPUT116), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1116), .A2(new_n1118), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1114), .A2(KEYINPUT117), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n768), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT117), .B1(new_n1114), .B2(new_n1121), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n759), .B1(new_n336), .B2(new_n863), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  OR2_X1    g0925(.A1(new_n902), .A2(new_n906), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n816), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1101), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1086), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n914), .B1(new_n741), .B2(new_n837), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1098), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n910), .B1(new_n1096), .B2(new_n1131), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n457), .A2(new_n741), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n918), .A2(new_n658), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1100), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1137), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1097), .A2(new_n1099), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1140), .A2(new_n708), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1129), .A2(new_n1143), .ZN(G378));
  INV_X1    g0944(.A(new_n917), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n715), .B1(new_n931), .B2(new_n932), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n930), .A2(new_n1146), .A3(KEYINPUT122), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n361), .A2(new_n689), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n657), .A2(new_n362), .A3(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n654), .A2(new_n656), .A3(new_n362), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1150), .A2(new_n361), .A3(new_n689), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n1149), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1152), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1147), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(KEYINPUT122), .B1(new_n930), .B2(new_n1146), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AOI211_X1 g0958(.A(KEYINPUT122), .B(new_n1155), .C1(new_n930), .C2(new_n1146), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1145), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n930), .A2(new_n1146), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT122), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1164), .A2(new_n1147), .A3(new_n1155), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1161), .A2(new_n1165), .A3(new_n917), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1160), .A2(new_n758), .A3(new_n1166), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n776), .A2(new_n711), .B1(new_n778), .B2(new_n409), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n990), .B(new_n1168), .C1(G77), .C2(new_n781), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n327), .A2(G41), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n796), .A2(new_n338), .B1(new_n790), .B2(new_n478), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(G107), .C2(new_n844), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1169), .B(new_n1172), .C1(new_n205), .C2(new_n786), .ZN(new_n1173));
  XOR2_X1   g0973(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n1174));
  OR2_X1    g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1170), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n771), .A2(new_n357), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n776), .A2(new_n1108), .B1(new_n796), .B2(new_n846), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(G132), .C2(new_n787), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n794), .A2(new_n1105), .B1(new_n780), .B2(new_n1102), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT119), .Z(new_n1183));
  NAND2_X1  g0983(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1184), .A2(KEYINPUT59), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(KEYINPUT59), .ZN(new_n1186));
  AOI211_X1 g0986(.A(G33), .B(G41), .C1(new_n803), .C2(G124), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n791), .B2(new_n778), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT120), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1185), .A2(new_n1186), .A3(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n768), .B1(new_n1178), .B2(new_n1190), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT121), .Z(new_n1192));
  AOI211_X1 g0992(.A(new_n762), .B(new_n1192), .C1(new_n202), .C2(new_n864), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1155), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1193), .B1(new_n1194), .B2(new_n816), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1167), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1142), .A2(new_n1138), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1197), .A2(new_n1160), .A3(KEYINPUT57), .A4(new_n1166), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n708), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT57), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1197), .A2(new_n1160), .A3(new_n1166), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1199), .A2(KEYINPUT123), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT123), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1198), .A2(new_n1203), .A3(new_n708), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1196), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(G375));
  INV_X1    g1006(.A(new_n964), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1133), .A2(new_n1137), .A3(new_n1134), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1139), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1095), .A2(new_n1127), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n327), .B1(new_n803), .B2(G303), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n206), .B2(new_n796), .C1(new_n478), .C2(new_n794), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n775), .A2(G294), .B1(new_n781), .B2(G97), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1214), .B1(new_n308), .B2(new_n778), .C1(new_n338), .C2(new_n771), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1213), .B(new_n1215), .C1(new_n1029), .C2(new_n787), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(G150), .A2(new_n797), .B1(new_n803), .B2(G128), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1217), .B(new_n327), .C1(new_n846), .C2(new_n794), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n775), .A2(G132), .B1(new_n811), .B2(G58), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(new_n202), .B2(new_n771), .C1(new_n791), .C2(new_n780), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1218), .B(new_n1220), .C1(new_n787), .C2(new_n1103), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n768), .B1(new_n1216), .B2(new_n1221), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n759), .B(new_n1222), .C1(new_n863), .C2(G68), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT124), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1211), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n1135), .B2(new_n758), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1209), .A2(new_n1226), .ZN(G381));
  NAND3_X1  g1027(.A1(new_n1052), .A2(new_n1054), .A3(new_n829), .ZN(new_n1228));
  NOR4_X1   g1028(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1013), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(KEYINPUT125), .ZN(new_n1231));
  INV_X1    g1031(.A(G378), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1205), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT125), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1013), .A2(new_n1235), .A3(new_n1229), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1231), .A2(new_n1234), .A3(new_n1236), .ZN(G407));
  OAI211_X1 g1037(.A(G407), .B(G213), .C1(G343), .C2(new_n1233), .ZN(G409));
  NOR2_X1   g1038(.A1(new_n688), .A2(G343), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(G378), .A2(new_n1196), .ZN(new_n1240));
  OR2_X1    g1040(.A1(new_n1201), .A2(new_n964), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1239), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT126), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(G384), .A2(new_n1243), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1133), .A2(KEYINPUT60), .A3(new_n1137), .A4(new_n1134), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n708), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1139), .A2(KEYINPUT60), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1246), .B1(new_n1247), .B2(new_n1208), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1226), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1244), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(G384), .A2(new_n1243), .ZN(new_n1251));
  OR2_X1    g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1242), .B(new_n1254), .C1(new_n1205), .C2(new_n1232), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(KEYINPUT62), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT61), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1239), .A2(G2897), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1252), .A2(new_n1253), .A3(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1258), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1203), .B1(new_n1198), .B2(new_n708), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1201), .A2(new_n1200), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1263), .A2(new_n1265), .A3(new_n1204), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1196), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1232), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1242), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1261), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1198), .A2(new_n1203), .A3(new_n708), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1271), .A2(new_n1262), .A3(new_n1264), .ZN(new_n1272));
  OAI21_X1  g1072(.A(G378), .B1(new_n1272), .B2(new_n1196), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT62), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1273), .A2(new_n1274), .A3(new_n1242), .A4(new_n1254), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1256), .A2(new_n1257), .A3(new_n1270), .A4(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(G393), .A2(G396), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1228), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1011), .ZN(new_n1279));
  MUX2_X1   g1079(.A(new_n1279), .B(new_n1278), .S(G390), .Z(new_n1280));
  XNOR2_X1  g1080(.A(new_n1280), .B(new_n1009), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1276), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1273), .A2(new_n1242), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT61), .B1(new_n1284), .B2(new_n1261), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT63), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1255), .A2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1273), .A2(KEYINPUT63), .A3(new_n1242), .A4(new_n1254), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1285), .A2(new_n1281), .A3(new_n1287), .A4(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1283), .A2(new_n1289), .ZN(G405));
  NAND3_X1  g1090(.A1(new_n1233), .A2(new_n1273), .A3(new_n1254), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1254), .B1(new_n1233), .B2(new_n1273), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1282), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1293), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1295), .A2(new_n1281), .A3(new_n1291), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1294), .A2(new_n1296), .ZN(G402));
endmodule


