//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  INV_X1    g000(.A(G107), .ZN(new_n187));
  AND2_X1   g001(.A1(KEYINPUT91), .A2(G122), .ZN(new_n188));
  NOR2_X1   g002(.A1(KEYINPUT91), .A2(G122), .ZN(new_n189));
  OAI21_X1  g003(.A(G116), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT92), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT92), .ZN(new_n192));
  OAI211_X1 g006(.A(new_n192), .B(G116), .C1(new_n188), .C2(new_n189), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G122), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT93), .B1(new_n195), .B2(G116), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT93), .ZN(new_n197));
  INV_X1    g011(.A(G116), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G122), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(new_n199), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n194), .A2(KEYINPUT94), .A3(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(KEYINPUT94), .B1(new_n194), .B2(new_n200), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n187), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G128), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  XNOR2_X1  g023(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n194), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n200), .B(KEYINPUT14), .ZN(new_n212));
  OAI21_X1  g026(.A(G107), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT97), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n213), .A2(new_n214), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n203), .B(new_n210), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n194), .A2(new_n200), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT94), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n194), .A2(KEYINPUT94), .A3(new_n200), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(G107), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT95), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n203), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n208), .A2(new_n209), .ZN(new_n225));
  XOR2_X1   g039(.A(new_n225), .B(KEYINPUT96), .Z(new_n226));
  NAND2_X1  g040(.A1(new_n207), .A2(KEYINPUT13), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n205), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n204), .A2(KEYINPUT13), .A3(G128), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n209), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n224), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n223), .B1(new_n203), .B2(new_n222), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n217), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT9), .B(G234), .ZN(new_n235));
  INV_X1    g049(.A(G217), .ZN(new_n236));
  NOR3_X1   g050(.A1(new_n235), .A2(new_n236), .A3(G953), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n217), .B(new_n237), .C1(new_n232), .C2(new_n233), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G902), .ZN(new_n242));
  INV_X1    g056(.A(G478), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n243), .A2(KEYINPUT15), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n241), .A2(new_n242), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(G475), .A2(G902), .ZN(new_n248));
  XOR2_X1   g062(.A(new_n248), .B(KEYINPUT90), .Z(new_n249));
  INV_X1    g063(.A(KEYINPUT87), .ZN(new_n250));
  INV_X1    g064(.A(G140), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G125), .ZN(new_n252));
  INV_X1    g066(.A(G125), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G140), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G146), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n255), .A2(G146), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(G237), .A2(G953), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(G143), .A3(G214), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT86), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n261), .A2(KEYINPUT86), .A3(G143), .A4(G214), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n261), .A2(G214), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n204), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT18), .ZN(new_n270));
  INV_X1    g084(.A(G131), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n260), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n264), .A2(new_n265), .B1(new_n204), .B2(new_n267), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n274), .A2(new_n270), .A3(new_n271), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n250), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n272), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n274), .A2(new_n277), .B1(new_n258), .B2(new_n259), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n269), .A2(G131), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n278), .B(KEYINPUT87), .C1(new_n279), .C2(new_n270), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n255), .A2(KEYINPUT72), .A3(KEYINPUT16), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n252), .A2(KEYINPUT72), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(new_n251), .A3(G125), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT16), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(G146), .B1(new_n283), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n287), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(new_n257), .A3(new_n282), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n269), .A2(KEYINPUT17), .A3(G131), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n274), .A2(new_n271), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n279), .A2(new_n293), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n291), .B(new_n292), .C1(new_n294), .C2(KEYINPUT17), .ZN(new_n295));
  XNOR2_X1  g109(.A(G113), .B(G122), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT89), .B(G104), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n296), .B(new_n297), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n281), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT88), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n256), .A2(new_n300), .A3(KEYINPUT19), .ZN(new_n301));
  XOR2_X1   g115(.A(KEYINPUT88), .B(KEYINPUT19), .Z(new_n302));
  OAI21_X1  g116(.A(new_n301), .B1(new_n256), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n257), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n294), .A2(new_n288), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n298), .B1(new_n281), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n249), .B1(new_n299), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT20), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n281), .A2(new_n305), .ZN(new_n309));
  INV_X1    g123(.A(new_n298), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n281), .A2(new_n295), .A3(new_n298), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT20), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(new_n249), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n308), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n298), .B1(new_n281), .B2(new_n295), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n242), .B1(new_n299), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G475), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n245), .B1(new_n241), .B2(new_n242), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n247), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(G214), .B1(G237), .B2(G902), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(G110), .B(G122), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G104), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT3), .B1(new_n327), .B2(G107), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n187), .A3(G104), .ZN(new_n330));
  INV_X1    g144(.A(G101), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(G107), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n328), .A2(new_n330), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT4), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n328), .A2(new_n330), .A3(new_n332), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT73), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n328), .A2(new_n330), .A3(KEYINPUT73), .A4(new_n332), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n334), .B1(new_n339), .B2(G101), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G119), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G116), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n198), .A2(G119), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT66), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT2), .B(G113), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n348), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(new_n345), .A3(new_n346), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n331), .B1(new_n337), .B2(new_n338), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n341), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n327), .A2(G107), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n187), .A2(G104), .ZN(new_n359));
  OAI21_X1  g173(.A(G101), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n333), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n333), .A2(new_n360), .A3(KEYINPUT75), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n345), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT5), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n343), .A2(KEYINPUT5), .ZN(new_n368));
  INV_X1    g182(.A(G113), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n367), .A2(new_n370), .B1(new_n350), .B2(new_n366), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n357), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n356), .B1(new_n341), .B2(new_n355), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n326), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n339), .A2(new_n354), .A3(G101), .ZN(new_n376));
  INV_X1    g190(.A(new_n352), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT82), .B1(new_n378), .B2(new_n340), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n379), .A2(new_n357), .A3(new_n372), .A4(new_n325), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n375), .A2(KEYINPUT6), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT6), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n382), .B(new_n326), .C1(new_n373), .C2(new_n374), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n257), .A2(G143), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n204), .A2(G146), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(KEYINPUT0), .A2(G128), .ZN(new_n387));
  NAND2_X1  g201(.A1(KEYINPUT0), .A2(G128), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n386), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(G143), .B(G146), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n388), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(G125), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n384), .A2(new_n385), .A3(G128), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT1), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT64), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT64), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT1), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT65), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT65), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n391), .A2(new_n402), .A3(new_n403), .A4(G128), .ZN(new_n404));
  INV_X1    g218(.A(new_n384), .ZN(new_n405));
  OAI21_X1  g219(.A(G128), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n401), .A2(new_n404), .B1(new_n406), .B2(new_n386), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n394), .B1(new_n407), .B2(new_n253), .ZN(new_n408));
  INV_X1    g222(.A(G953), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G224), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n408), .B(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n381), .A2(new_n383), .A3(new_n411), .ZN(new_n412));
  AND4_X1   g226(.A1(new_n379), .A2(new_n357), .A3(new_n372), .A4(new_n325), .ZN(new_n413));
  OAI211_X1 g227(.A(KEYINPUT7), .B(new_n410), .C1(new_n408), .C2(KEYINPUT84), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n401), .A2(new_n404), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n406), .A2(new_n386), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n393), .B1(new_n417), .B2(G125), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n410), .A2(KEYINPUT7), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n410), .A2(KEYINPUT84), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  XOR2_X1   g235(.A(new_n325), .B(KEYINPUT8), .Z(new_n422));
  NAND3_X1  g236(.A1(new_n333), .A2(new_n360), .A3(KEYINPUT83), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n422), .B1(new_n371), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n424), .B1(new_n371), .B2(new_n423), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n414), .A2(new_n421), .A3(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(KEYINPUT85), .B(new_n242), .C1(new_n413), .C2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n242), .B1(new_n413), .B2(new_n426), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT85), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n412), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(G210), .B1(G237), .B2(G902), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n412), .A2(new_n430), .A3(new_n432), .A4(new_n427), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n324), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G952), .ZN(new_n437));
  AOI211_X1 g251(.A(G953), .B(new_n437), .C1(G234), .C2(G237), .ZN(new_n438));
  AOI211_X1 g252(.A(new_n242), .B(new_n409), .C1(G234), .C2(G237), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(G898), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n322), .A2(new_n436), .A3(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT79), .B(G469), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT11), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(new_n209), .B2(G137), .ZN(new_n446));
  INV_X1    g260(.A(G137), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(KEYINPUT11), .A3(G134), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n209), .A2(G137), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n446), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G131), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n446), .A2(new_n448), .A3(new_n271), .A4(new_n449), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n453), .A2(KEYINPUT76), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n415), .A2(new_n416), .A3(new_n361), .ZN(new_n455));
  OAI22_X1  g269(.A1(new_n391), .A2(G128), .B1(new_n396), .B2(new_n385), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n456), .B1(new_n401), .B2(new_n404), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(new_n361), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n454), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT12), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n390), .A2(new_n392), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n376), .B(new_n461), .C1(new_n353), .C2(new_n334), .ZN(new_n462));
  INV_X1    g276(.A(new_n453), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n417), .A2(new_n364), .A3(KEYINPUT10), .A4(new_n363), .ZN(new_n464));
  XNOR2_X1  g278(.A(KEYINPUT74), .B(KEYINPUT10), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n465), .B1(new_n457), .B2(new_n361), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n462), .A2(new_n463), .A3(new_n464), .A4(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT12), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n454), .B(new_n468), .C1(new_n455), .C2(new_n458), .ZN(new_n469));
  XNOR2_X1  g283(.A(G110), .B(G140), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n409), .A2(G227), .ZN(new_n471));
  XOR2_X1   g285(.A(new_n470), .B(new_n471), .Z(new_n472));
  NAND4_X1  g286(.A1(new_n460), .A2(new_n467), .A3(new_n469), .A4(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n464), .A2(new_n466), .ZN(new_n475));
  AOI211_X1 g289(.A(KEYINPUT4), .B(new_n331), .C1(new_n337), .C2(new_n338), .ZN(new_n476));
  INV_X1    g290(.A(new_n461), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n340), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n453), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n472), .B1(new_n479), .B2(new_n467), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n242), .B(new_n444), .C1(new_n474), .C2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT80), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n472), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n457), .A2(new_n361), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT10), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n407), .A2(new_n486), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n485), .A2(new_n465), .B1(new_n487), .B2(new_n365), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n463), .B1(new_n488), .B2(new_n462), .ZN(new_n489));
  INV_X1    g303(.A(new_n467), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n484), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n473), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n492), .A2(KEYINPUT80), .A3(new_n242), .A4(new_n444), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n483), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT78), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n479), .A2(new_n467), .A3(new_n472), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n460), .A2(new_n467), .A3(new_n469), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n497), .A2(KEYINPUT77), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT77), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n460), .A2(new_n467), .A3(new_n499), .A4(new_n469), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n484), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n495), .B(new_n496), .C1(new_n498), .C2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n497), .A2(KEYINPUT77), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(new_n500), .A3(new_n484), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n495), .B1(new_n505), .B2(new_n496), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n242), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n494), .B1(new_n507), .B2(G469), .ZN(new_n508));
  INV_X1    g322(.A(G221), .ZN(new_n509));
  INV_X1    g323(.A(new_n235), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n509), .B1(new_n510), .B2(new_n242), .ZN(new_n511));
  OAI21_X1  g325(.A(KEYINPUT81), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n483), .A2(new_n493), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n496), .B1(new_n498), .B2(new_n501), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT78), .ZN(new_n515));
  AOI21_X1  g329(.A(G902), .B1(new_n515), .B2(new_n502), .ZN(new_n516));
  INV_X1    g330(.A(G469), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT81), .ZN(new_n519));
  INV_X1    g333(.A(new_n511), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n443), .B1(new_n512), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n453), .A2(new_n461), .ZN(new_n523));
  INV_X1    g337(.A(new_n449), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n209), .A2(G137), .ZN(new_n525));
  OAI21_X1  g339(.A(G131), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n452), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n523), .B(new_n352), .C1(new_n407), .C2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT67), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n527), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n417), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n532), .A2(KEYINPUT67), .A3(new_n523), .A4(new_n352), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n527), .B1(new_n415), .B2(new_n416), .ZN(new_n535));
  AOI22_X1  g349(.A1(new_n451), .A2(new_n452), .B1(new_n390), .B2(new_n392), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT30), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT30), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n523), .B(new_n538), .C1(new_n407), .C2(new_n527), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n377), .ZN(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT26), .B(G101), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n261), .A2(G210), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n534), .A2(new_n541), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT31), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n534), .A2(new_n541), .A3(KEYINPUT31), .A4(new_n546), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n377), .B1(new_n535), .B2(new_n536), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n530), .A2(new_n533), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT28), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT28), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n528), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n546), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(KEYINPUT69), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT69), .ZN(new_n560));
  INV_X1    g374(.A(new_n556), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(new_n553), .B2(KEYINPUT28), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n560), .B1(new_n562), .B2(new_n546), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n551), .A2(new_n559), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(G472), .A2(G902), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(KEYINPUT32), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT70), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n564), .A2(new_n565), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT32), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT29), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n534), .A2(new_n541), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n572), .B1(new_n573), .B2(new_n546), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n557), .A2(new_n558), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n242), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n557), .A2(new_n572), .A3(new_n558), .ZN(new_n577));
  OAI21_X1  g391(.A(G472), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n564), .A2(KEYINPUT70), .A3(KEYINPUT32), .A4(new_n565), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n568), .A2(new_n571), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT23), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n581), .B1(new_n342), .B2(G128), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n206), .A2(KEYINPUT23), .A3(G119), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n582), .B(new_n583), .C1(G119), .C2(new_n206), .ZN(new_n584));
  XNOR2_X1  g398(.A(G119), .B(G128), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT24), .B(G110), .Z(new_n586));
  OAI22_X1  g400(.A1(new_n584), .A2(G110), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n288), .A2(new_n587), .A3(new_n258), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n584), .A2(G110), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n586), .A2(new_n585), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n588), .B1(new_n291), .B2(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(KEYINPUT22), .B(G137), .Z(new_n593));
  NAND3_X1  g407(.A1(new_n409), .A2(G221), .A3(G234), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n592), .B(new_n595), .Z(new_n596));
  INV_X1    g410(.A(KEYINPUT25), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n597), .A3(new_n242), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n592), .B(new_n595), .ZN(new_n599));
  OAI21_X1  g413(.A(KEYINPUT25), .B1(new_n599), .B2(G902), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n236), .B1(G234), .B2(new_n242), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(KEYINPUT71), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n598), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(G902), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n596), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n580), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n522), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT98), .B(G101), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G3));
  NAND2_X1  g425(.A1(new_n512), .A2(new_n521), .ZN(new_n612));
  INV_X1    g426(.A(new_n569), .ZN(new_n613));
  INV_X1    g427(.A(G472), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n564), .B2(new_n242), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n607), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  AOI211_X1 g432(.A(G478), .B(G902), .C1(new_n239), .C2(new_n240), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT33), .B1(new_n237), .B2(KEYINPUT99), .ZN(new_n620));
  INV_X1    g434(.A(new_n240), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n203), .A2(new_n222), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(KEYINPUT95), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(new_n224), .A3(new_n231), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n237), .B1(new_n624), .B2(new_n217), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n620), .B1(new_n621), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n620), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n239), .A2(new_n240), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n626), .A2(new_n242), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n619), .B1(new_n629), .B2(G478), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n436), .A2(new_n630), .A3(new_n320), .A4(new_n442), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n612), .A2(new_n618), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT100), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT34), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G104), .ZN(G6));
  NOR2_X1   g450(.A1(new_n621), .A2(new_n625), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n244), .B1(new_n637), .B2(G902), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n320), .B1(new_n638), .B2(new_n246), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(new_n436), .A3(new_n442), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n612), .A2(new_n618), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  INV_X1    g458(.A(new_n443), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n595), .A2(KEYINPUT36), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n592), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n604), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n603), .A2(new_n648), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n613), .A2(new_n615), .A3(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n508), .A2(KEYINPUT81), .A3(new_n511), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n519), .B1(new_n518), .B2(new_n520), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n645), .B(new_n650), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT101), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT102), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  NAND2_X1  g471(.A1(new_n580), .A2(new_n436), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n639), .ZN(new_n660));
  INV_X1    g474(.A(G900), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n439), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n438), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n660), .A2(new_n649), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n612), .A2(new_n659), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  XNOR2_X1  g482(.A(new_n664), .B(KEYINPUT39), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n612), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  AOI22_X1  g487(.A1(new_n308), .A2(new_n315), .B1(G475), .B2(new_n318), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n638), .B2(new_n246), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n675), .A2(new_n323), .A3(new_n649), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n434), .A2(new_n435), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT38), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n553), .A2(new_n558), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n547), .A2(G472), .A3(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n614), .A2(new_n242), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n685), .B(KEYINPUT103), .Z(new_n686));
  NAND4_X1  g500(.A1(new_n568), .A2(new_n686), .A3(new_n571), .A4(new_n579), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n675), .A2(KEYINPUT104), .A3(new_n323), .A4(new_n649), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n678), .A2(new_n680), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n689), .A2(KEYINPUT105), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(KEYINPUT105), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n672), .A2(new_n673), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G143), .ZN(G45));
  NAND3_X1  g507(.A1(new_n630), .A2(new_n320), .A3(new_n664), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n694), .A2(new_n649), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n612), .A2(new_n659), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G146), .ZN(G48));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n492), .A2(new_n242), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(G469), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n513), .A2(new_n520), .A3(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n513), .A2(KEYINPUT107), .A3(new_n520), .A4(new_n700), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n580), .A3(new_n607), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n698), .B1(new_n706), .B2(new_n631), .ZN(new_n707));
  AND4_X1   g521(.A1(new_n580), .A2(new_n607), .A3(new_n703), .A4(new_n704), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(KEYINPUT108), .A3(new_n632), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT41), .B(G113), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  NAND3_X1  g526(.A1(new_n608), .A2(new_n641), .A3(new_n705), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G116), .ZN(G18));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n649), .A2(new_n441), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n580), .A2(new_n322), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n703), .A2(new_n436), .A3(new_n704), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n715), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n703), .A2(new_n436), .A3(new_n704), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n322), .A2(new_n716), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(KEYINPUT109), .A3(new_n580), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  NAND2_X1  g538(.A1(new_n557), .A2(new_n558), .ZN(new_n725));
  AOI211_X1 g539(.A(G472), .B(G902), .C1(new_n551), .C2(new_n725), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n615), .A2(new_n726), .A3(new_n606), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n703), .A3(new_n704), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n436), .A2(new_n675), .A3(new_n442), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n195), .ZN(G24));
  NOR3_X1   g545(.A1(new_n615), .A2(new_n649), .A3(new_n726), .ZN(new_n732));
  AOI211_X1 g546(.A(new_n619), .B(new_n674), .C1(new_n629), .C2(G478), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(new_n733), .A3(new_n664), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n718), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n253), .ZN(G27));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n571), .B(new_n578), .C1(new_n737), .C2(new_n566), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n566), .A2(new_n737), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n607), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n434), .A2(new_n323), .A3(new_n435), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(G469), .A2(G902), .ZN(new_n743));
  XOR2_X1   g557(.A(new_n743), .B(KEYINPUT110), .Z(new_n744));
  INV_X1    g558(.A(new_n514), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n744), .B1(new_n745), .B2(G469), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n511), .B1(new_n746), .B2(new_n513), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n733), .A2(new_n664), .A3(new_n742), .A4(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(KEYINPUT42), .B1(new_n740), .B2(new_n748), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n742), .A2(new_n747), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n694), .A2(KEYINPUT42), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n608), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n271), .ZN(G33));
  NOR2_X1   g568(.A1(new_n660), .A2(new_n665), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n608), .A2(new_n755), .A3(new_n750), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G134), .ZN(G36));
  NAND2_X1  g571(.A1(new_n630), .A2(new_n674), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT43), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n758), .A2(KEYINPUT43), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n616), .A2(new_n649), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n758), .B(new_n760), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(KEYINPUT44), .A3(new_n763), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n768), .A3(new_n742), .ZN(new_n769));
  INV_X1    g583(.A(new_n744), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT45), .B1(new_n515), .B2(new_n502), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT45), .ZN(new_n772));
  OAI21_X1  g586(.A(G469), .B1(new_n514), .B2(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(KEYINPUT46), .B(new_n770), .C1(new_n771), .C2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(KEYINPUT112), .A3(new_n513), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n771), .A2(new_n773), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n744), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n775), .B1(KEYINPUT46), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT112), .B1(new_n774), .B2(new_n513), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n520), .B(new_n669), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n769), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(new_n447), .ZN(G39));
  NOR3_X1   g596(.A1(new_n694), .A2(new_n607), .A3(new_n741), .ZN(new_n783));
  INV_X1    g597(.A(new_n580), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n520), .B1(new_n778), .B2(new_n779), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT47), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g602(.A(KEYINPUT47), .B(new_n520), .C1(new_n778), .C2(new_n779), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n785), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(new_n251), .ZN(G42));
  NAND2_X1  g605(.A1(new_n513), .A2(new_n700), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT49), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n606), .A2(new_n511), .A3(new_n324), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n759), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT113), .ZN(new_n796));
  INV_X1    g610(.A(new_n687), .ZN(new_n797));
  XOR2_X1   g611(.A(new_n679), .B(KEYINPUT38), .Z(new_n798));
  OR2_X1    g612(.A1(new_n792), .A2(KEYINPUT49), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n796), .A2(new_n797), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n324), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(new_n728), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n761), .A2(new_n438), .A3(new_n762), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT50), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n806));
  NOR4_X1   g620(.A1(new_n803), .A2(new_n801), .A3(new_n806), .A4(new_n728), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n788), .B(new_n789), .C1(new_n520), .C2(new_n792), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n804), .A2(new_n727), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n741), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n808), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n705), .A2(new_n742), .ZN(new_n813));
  NOR4_X1   g627(.A1(new_n813), .A2(new_n606), .A3(new_n663), .A4(new_n687), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n630), .A2(new_n320), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n803), .A2(new_n813), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n814), .A2(new_n815), .B1(new_n816), .B2(new_n732), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n819));
  AOI211_X1 g633(.A(new_n819), .B(new_n808), .C1(new_n809), .C2(new_n811), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n818), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n812), .A2(new_n819), .A3(KEYINPUT51), .A4(new_n817), .ZN(new_n823));
  AOI211_X1 g637(.A(new_n437), .B(G953), .C1(new_n814), .C2(new_n733), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n824), .B1(new_n718), .B2(new_n810), .ZN(new_n825));
  INV_X1    g639(.A(new_n740), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n816), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n822), .A2(new_n823), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n832));
  INV_X1    g646(.A(new_n735), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n436), .A2(new_n675), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n649), .A2(new_n664), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n834), .A2(new_n687), .A3(new_n747), .A4(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n667), .A2(new_n696), .A3(new_n833), .A4(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n658), .B1(new_n521), .B2(new_n512), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n735), .B1(new_n840), .B2(new_n666), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(KEYINPUT52), .A3(new_n696), .A4(new_n836), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n749), .A2(new_n752), .A3(new_n756), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n665), .B1(new_n603), .B2(new_n648), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n580), .A2(new_n322), .A3(new_n742), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n612), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n732), .A2(new_n733), .A3(new_n664), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n750), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n844), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n730), .B1(new_n522), .B2(new_n608), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n852), .A2(new_n723), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n653), .A2(new_n713), .ZN(new_n854));
  AOI221_X4 g668(.A(new_n617), .B1(new_n631), .B2(new_n640), .C1(new_n512), .C2(new_n521), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n851), .A2(new_n853), .A3(new_n710), .A4(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n843), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n522), .A2(new_n650), .B1(new_n708), .B2(new_n641), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n612), .B(new_n618), .C1(new_n632), .C2(new_n641), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(new_n852), .A3(new_n723), .A4(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n707), .A2(new_n709), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n846), .A2(new_n612), .B1(new_n848), .B2(new_n750), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(new_n749), .A3(new_n752), .A4(new_n756), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n839), .A2(new_n842), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT53), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n832), .B1(new_n859), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n858), .B1(new_n843), .B2(new_n857), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n866), .A2(KEYINPUT53), .A3(new_n867), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(KEYINPUT54), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n831), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(G952), .A2(G953), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n800), .B1(new_n873), .B2(new_n874), .ZN(G75));
  AOI21_X1  g689(.A(new_n242), .B1(new_n870), .B2(new_n871), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(G210), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT56), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n381), .A2(new_n383), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(new_n411), .ZN(new_n880));
  XNOR2_X1  g694(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n880), .B(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n877), .A2(new_n878), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n882), .B1(new_n877), .B2(new_n878), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n409), .A2(G952), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(G51));
  XNOR2_X1  g700(.A(new_n744), .B(KEYINPUT57), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n869), .A2(new_n872), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n492), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n876), .A2(new_n776), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n885), .B1(new_n889), .B2(new_n890), .ZN(G54));
  NAND2_X1  g705(.A1(KEYINPUT58), .A2(G475), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT117), .Z(new_n893));
  AND3_X1   g707(.A1(new_n876), .A2(new_n313), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n313), .B1(new_n876), .B2(new_n893), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n894), .A2(new_n895), .A3(new_n885), .ZN(G60));
  NAND2_X1  g710(.A1(G478), .A2(G902), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT59), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n869), .A2(new_n872), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n626), .A2(new_n628), .ZN(new_n900));
  OAI22_X1  g714(.A1(new_n899), .A2(new_n900), .B1(G952), .B2(new_n409), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n900), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n899), .A2(KEYINPUT118), .A3(new_n900), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n901), .B1(new_n904), .B2(new_n905), .ZN(G63));
  NAND2_X1  g720(.A1(G217), .A2(G902), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT60), .Z(new_n908));
  OAI21_X1  g722(.A(new_n908), .B1(new_n859), .B2(new_n868), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n885), .B1(new_n909), .B2(new_n599), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n870), .A2(new_n871), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n647), .B(KEYINPUT119), .ZN(new_n913));
  AND4_X1   g727(.A1(new_n911), .A2(new_n912), .A3(new_n908), .A4(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n908), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n870), .B2(new_n871), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n911), .B1(new_n916), .B2(new_n913), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n910), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g734(.A(KEYINPUT61), .B(new_n910), .C1(new_n914), .C2(new_n917), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(G66));
  NOR2_X1   g736(.A1(new_n862), .A2(new_n863), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(G224), .A2(G953), .ZN(new_n925));
  OAI22_X1  g739(.A1(new_n924), .A2(G953), .B1(new_n440), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n879), .B1(G898), .B2(new_n409), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n926), .B(new_n927), .Z(G69));
  OAI211_X1 g742(.A(new_n608), .B(new_n742), .C1(new_n733), .C2(new_n639), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n929), .A2(new_n670), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n790), .A2(new_n781), .A3(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n841), .A2(new_n696), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n692), .A2(KEYINPUT62), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT62), .B1(new_n692), .B2(new_n932), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n409), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n540), .B(KEYINPUT121), .Z(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(new_n303), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n409), .A2(G900), .ZN(new_n940));
  INV_X1    g754(.A(new_n780), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n941), .A2(new_n742), .A3(new_n766), .A4(new_n768), .ZN(new_n942));
  INV_X1    g756(.A(new_n844), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n942), .A2(new_n932), .A3(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n790), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n941), .A2(new_n834), .A3(new_n826), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n944), .A2(KEYINPUT123), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT123), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n942), .A2(new_n946), .A3(new_n932), .A4(new_n943), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n948), .B1(new_n949), .B2(new_n790), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n940), .B1(new_n951), .B2(new_n409), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n939), .B1(new_n952), .B2(new_n938), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n409), .B1(G227), .B2(G900), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT122), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT124), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n955), .B1(new_n939), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  OAI221_X1 g772(.A(new_n939), .B1(new_n956), .B2(new_n955), .C1(new_n952), .C2(new_n938), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(G72));
  XNOR2_X1  g774(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n684), .B(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(new_n935), .B2(new_n924), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(KEYINPUT126), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT126), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n966), .B(new_n963), .C1(new_n935), .C2(new_n924), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n573), .A2(new_n558), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n965), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n963), .B1(new_n951), .B2(new_n924), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n970), .A2(new_n558), .A3(new_n573), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n573), .A2(new_n546), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n962), .B1(new_n972), .B2(new_n547), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n885), .B1(new_n912), .B2(new_n973), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n969), .A2(new_n971), .A3(new_n974), .ZN(G57));
endmodule


