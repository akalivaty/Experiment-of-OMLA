

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(n690), .A2(n689), .ZN(n694) );
  XNOR2_X1 U549 ( .A(KEYINPUT95), .B(KEYINPUT30), .ZN(n676) );
  NAND2_X1 U550 ( .A1(n867), .A2(G137), .ZN(n518) );
  AND2_X1 U551 ( .A1(n863), .A2(G125), .ZN(n510) );
  AND2_X1 U552 ( .A1(n679), .A2(n678), .ZN(n511) );
  INV_X1 U553 ( .A(n711), .ZN(n695) );
  XNOR2_X1 U554 ( .A(n677), .B(n676), .ZN(n679) );
  NAND2_X1 U555 ( .A1(n671), .A2(n767), .ZN(n711) );
  NAND2_X1 U556 ( .A1(G8), .A2(n711), .ZN(n748) );
  INV_X1 U557 ( .A(KEYINPUT17), .ZN(n515) );
  NOR2_X1 U558 ( .A1(G543), .A2(G651), .ZN(n635) );
  NOR2_X1 U559 ( .A1(n620), .A2(G651), .ZN(n629) );
  NOR2_X1 U560 ( .A1(n803), .A2(n802), .ZN(n804) );
  AND2_X1 U561 ( .A1(n521), .A2(n520), .ZN(G160) );
  INV_X1 U562 ( .A(G2104), .ZN(n513) );
  NOR2_X2 U563 ( .A1(G2105), .A2(n513), .ZN(n868) );
  NAND2_X1 U564 ( .A1(G101), .A2(n868), .ZN(n512) );
  XNOR2_X1 U565 ( .A(KEYINPUT23), .B(n512), .ZN(n514) );
  AND2_X1 U566 ( .A1(n513), .A2(G2105), .ZN(n863) );
  NOR2_X1 U567 ( .A1(n514), .A2(n510), .ZN(n521) );
  NOR2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n516) );
  XNOR2_X2 U569 ( .A(n516), .B(n515), .ZN(n867) );
  AND2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n864) );
  NAND2_X1 U571 ( .A1(G113), .A2(n864), .ZN(n517) );
  NAND2_X1 U572 ( .A1(n518), .A2(n517), .ZN(n519) );
  XOR2_X1 U573 ( .A(KEYINPUT64), .B(n519), .Z(n520) );
  NAND2_X1 U574 ( .A1(n635), .A2(G89), .ZN(n522) );
  XNOR2_X1 U575 ( .A(n522), .B(KEYINPUT4), .ZN(n524) );
  XOR2_X1 U576 ( .A(KEYINPUT0), .B(G543), .Z(n620) );
  INV_X1 U577 ( .A(G651), .ZN(n526) );
  NOR2_X1 U578 ( .A1(n620), .A2(n526), .ZN(n626) );
  NAND2_X1 U579 ( .A1(G76), .A2(n626), .ZN(n523) );
  NAND2_X1 U580 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U581 ( .A(KEYINPUT5), .B(n525), .ZN(n534) );
  NAND2_X1 U582 ( .A1(n629), .A2(G51), .ZN(n530) );
  NOR2_X1 U583 ( .A1(G543), .A2(n526), .ZN(n527) );
  XOR2_X1 U584 ( .A(KEYINPUT66), .B(n527), .Z(n528) );
  XNOR2_X1 U585 ( .A(KEYINPUT1), .B(n528), .ZN(n630) );
  NAND2_X1 U586 ( .A1(G63), .A2(n630), .ZN(n529) );
  NAND2_X1 U587 ( .A1(n530), .A2(n529), .ZN(n532) );
  XOR2_X1 U588 ( .A(KEYINPUT6), .B(KEYINPUT74), .Z(n531) );
  XNOR2_X1 U589 ( .A(n532), .B(n531), .ZN(n533) );
  NAND2_X1 U590 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U591 ( .A(KEYINPUT7), .B(n535), .ZN(G168) );
  XOR2_X1 U592 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U593 ( .A1(n629), .A2(G53), .ZN(n537) );
  NAND2_X1 U594 ( .A1(G65), .A2(n630), .ZN(n536) );
  NAND2_X1 U595 ( .A1(n537), .A2(n536), .ZN(n541) );
  NAND2_X1 U596 ( .A1(G91), .A2(n635), .ZN(n539) );
  NAND2_X1 U597 ( .A1(G78), .A2(n626), .ZN(n538) );
  NAND2_X1 U598 ( .A1(n539), .A2(n538), .ZN(n540) );
  OR2_X1 U599 ( .A1(n541), .A2(n540), .ZN(G299) );
  NAND2_X1 U600 ( .A1(n629), .A2(G52), .ZN(n543) );
  NAND2_X1 U601 ( .A1(G64), .A2(n630), .ZN(n542) );
  NAND2_X1 U602 ( .A1(n543), .A2(n542), .ZN(n548) );
  NAND2_X1 U603 ( .A1(G90), .A2(n635), .ZN(n545) );
  NAND2_X1 U604 ( .A1(G77), .A2(n626), .ZN(n544) );
  NAND2_X1 U605 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U606 ( .A(KEYINPUT9), .B(n546), .Z(n547) );
  NOR2_X1 U607 ( .A1(n548), .A2(n547), .ZN(G171) );
  AND2_X1 U608 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U609 ( .A(G132), .ZN(G219) );
  INV_X1 U610 ( .A(G57), .ZN(G237) );
  INV_X1 U611 ( .A(G120), .ZN(G236) );
  INV_X1 U612 ( .A(G108), .ZN(G238) );
  NAND2_X1 U613 ( .A1(G7), .A2(G661), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n549), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U615 ( .A(G223), .ZN(n805) );
  NAND2_X1 U616 ( .A1(n805), .A2(G567), .ZN(n550) );
  XOR2_X1 U617 ( .A(KEYINPUT11), .B(n550), .Z(G234) );
  XOR2_X1 U618 ( .A(KEYINPUT14), .B(KEYINPUT69), .Z(n552) );
  NAND2_X1 U619 ( .A1(G56), .A2(n630), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n562) );
  NAND2_X1 U621 ( .A1(n629), .A2(G43), .ZN(n553) );
  XNOR2_X1 U622 ( .A(KEYINPUT71), .B(n553), .ZN(n560) );
  NAND2_X1 U623 ( .A1(n635), .A2(G81), .ZN(n554) );
  XNOR2_X1 U624 ( .A(n554), .B(KEYINPUT12), .ZN(n556) );
  NAND2_X1 U625 ( .A1(G68), .A2(n626), .ZN(n555) );
  NAND2_X1 U626 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U627 ( .A(KEYINPUT70), .B(n557), .Z(n558) );
  XNOR2_X1 U628 ( .A(KEYINPUT13), .B(n558), .ZN(n559) );
  NOR2_X1 U629 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U630 ( .A1(n562), .A2(n561), .ZN(n922) );
  INV_X1 U631 ( .A(n922), .ZN(n563) );
  NAND2_X1 U632 ( .A1(n563), .A2(G860), .ZN(G153) );
  XOR2_X1 U633 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  NAND2_X1 U634 ( .A1(G868), .A2(G301), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n635), .A2(G92), .ZN(n570) );
  NAND2_X1 U636 ( .A1(n629), .A2(G54), .ZN(n565) );
  NAND2_X1 U637 ( .A1(G66), .A2(n630), .ZN(n564) );
  NAND2_X1 U638 ( .A1(n565), .A2(n564), .ZN(n568) );
  NAND2_X1 U639 ( .A1(G79), .A2(n626), .ZN(n566) );
  XNOR2_X1 U640 ( .A(KEYINPUT73), .B(n566), .ZN(n567) );
  NOR2_X1 U641 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U642 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U643 ( .A(KEYINPUT15), .B(n571), .Z(n692) );
  INV_X1 U644 ( .A(G868), .ZN(n647) );
  NAND2_X1 U645 ( .A1(n692), .A2(n647), .ZN(n572) );
  NAND2_X1 U646 ( .A1(n573), .A2(n572), .ZN(G284) );
  NOR2_X1 U647 ( .A1(G286), .A2(n647), .ZN(n575) );
  NOR2_X1 U648 ( .A1(G868), .A2(G299), .ZN(n574) );
  NOR2_X1 U649 ( .A1(n575), .A2(n574), .ZN(G297) );
  INV_X1 U650 ( .A(G559), .ZN(n576) );
  NOR2_X1 U651 ( .A1(G860), .A2(n576), .ZN(n577) );
  XNOR2_X1 U652 ( .A(KEYINPUT75), .B(n577), .ZN(n578) );
  INV_X1 U653 ( .A(n692), .ZN(n901) );
  NAND2_X1 U654 ( .A1(n578), .A2(n901), .ZN(n579) );
  XNOR2_X1 U655 ( .A(n579), .B(KEYINPUT16), .ZN(n580) );
  XNOR2_X1 U656 ( .A(KEYINPUT76), .B(n580), .ZN(G148) );
  NOR2_X1 U657 ( .A1(G868), .A2(n922), .ZN(n583) );
  NAND2_X1 U658 ( .A1(G868), .A2(n901), .ZN(n581) );
  NOR2_X1 U659 ( .A1(G559), .A2(n581), .ZN(n582) );
  NOR2_X1 U660 ( .A1(n583), .A2(n582), .ZN(G282) );
  XNOR2_X1 U661 ( .A(G2100), .B(KEYINPUT79), .ZN(n594) );
  NAND2_X1 U662 ( .A1(G123), .A2(n863), .ZN(n584) );
  XOR2_X1 U663 ( .A(KEYINPUT77), .B(n584), .Z(n585) );
  XNOR2_X1 U664 ( .A(n585), .B(KEYINPUT18), .ZN(n587) );
  NAND2_X1 U665 ( .A1(G111), .A2(n864), .ZN(n586) );
  NAND2_X1 U666 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U667 ( .A1(G135), .A2(n867), .ZN(n589) );
  NAND2_X1 U668 ( .A1(G99), .A2(n868), .ZN(n588) );
  NAND2_X1 U669 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U670 ( .A1(n591), .A2(n590), .ZN(n930) );
  XNOR2_X1 U671 ( .A(n930), .B(G2096), .ZN(n592) );
  XNOR2_X1 U672 ( .A(n592), .B(KEYINPUT78), .ZN(n593) );
  NAND2_X1 U673 ( .A1(n594), .A2(n593), .ZN(G156) );
  NAND2_X1 U674 ( .A1(G559), .A2(n901), .ZN(n595) );
  XNOR2_X1 U675 ( .A(n595), .B(n922), .ZN(n644) );
  NOR2_X1 U676 ( .A1(n644), .A2(G860), .ZN(n604) );
  NAND2_X1 U677 ( .A1(n629), .A2(G55), .ZN(n597) );
  NAND2_X1 U678 ( .A1(G67), .A2(n630), .ZN(n596) );
  NAND2_X1 U679 ( .A1(n597), .A2(n596), .ZN(n600) );
  NAND2_X1 U680 ( .A1(G80), .A2(n626), .ZN(n598) );
  XNOR2_X1 U681 ( .A(KEYINPUT81), .B(n598), .ZN(n599) );
  NOR2_X1 U682 ( .A1(n600), .A2(n599), .ZN(n602) );
  NAND2_X1 U683 ( .A1(n635), .A2(G93), .ZN(n601) );
  NAND2_X1 U684 ( .A1(n602), .A2(n601), .ZN(n648) );
  XOR2_X1 U685 ( .A(n648), .B(KEYINPUT80), .Z(n603) );
  XNOR2_X1 U686 ( .A(n604), .B(n603), .ZN(G145) );
  NAND2_X1 U687 ( .A1(n629), .A2(G50), .ZN(n607) );
  NAND2_X1 U688 ( .A1(n630), .A2(G62), .ZN(n605) );
  XOR2_X1 U689 ( .A(KEYINPUT83), .B(n605), .Z(n606) );
  NAND2_X1 U690 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U691 ( .A1(G88), .A2(n635), .ZN(n609) );
  NAND2_X1 U692 ( .A1(G75), .A2(n626), .ZN(n608) );
  NAND2_X1 U693 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U694 ( .A1(n611), .A2(n610), .ZN(G166) );
  NAND2_X1 U695 ( .A1(n629), .A2(G47), .ZN(n614) );
  NAND2_X1 U696 ( .A1(G60), .A2(n630), .ZN(n612) );
  XOR2_X1 U697 ( .A(KEYINPUT67), .B(n612), .Z(n613) );
  NAND2_X1 U698 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U699 ( .A1(G85), .A2(n635), .ZN(n615) );
  XNOR2_X1 U700 ( .A(KEYINPUT65), .B(n615), .ZN(n616) );
  NOR2_X1 U701 ( .A1(n617), .A2(n616), .ZN(n619) );
  NAND2_X1 U702 ( .A1(n626), .A2(G72), .ZN(n618) );
  NAND2_X1 U703 ( .A1(n619), .A2(n618), .ZN(G290) );
  NAND2_X1 U704 ( .A1(G74), .A2(G651), .ZN(n622) );
  NAND2_X1 U705 ( .A1(G87), .A2(n620), .ZN(n621) );
  NAND2_X1 U706 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U707 ( .A1(n630), .A2(n623), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n629), .A2(G49), .ZN(n624) );
  NAND2_X1 U709 ( .A1(n625), .A2(n624), .ZN(G288) );
  XOR2_X1 U710 ( .A(KEYINPUT82), .B(KEYINPUT2), .Z(n628) );
  NAND2_X1 U711 ( .A1(G73), .A2(n626), .ZN(n627) );
  XNOR2_X1 U712 ( .A(n628), .B(n627), .ZN(n634) );
  NAND2_X1 U713 ( .A1(n629), .A2(G48), .ZN(n632) );
  NAND2_X1 U714 ( .A1(G61), .A2(n630), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U716 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n635), .A2(G86), .ZN(n636) );
  NAND2_X1 U718 ( .A1(n637), .A2(n636), .ZN(G305) );
  XNOR2_X1 U719 ( .A(G166), .B(G290), .ZN(n638) );
  XNOR2_X1 U720 ( .A(n638), .B(n648), .ZN(n639) );
  XNOR2_X1 U721 ( .A(KEYINPUT19), .B(n639), .ZN(n641) );
  XNOR2_X1 U722 ( .A(G288), .B(KEYINPUT84), .ZN(n640) );
  XNOR2_X1 U723 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U724 ( .A(n642), .B(G305), .ZN(n643) );
  XNOR2_X1 U725 ( .A(n643), .B(G299), .ZN(n878) );
  XNOR2_X1 U726 ( .A(n878), .B(n644), .ZN(n645) );
  NAND2_X1 U727 ( .A1(n645), .A2(G868), .ZN(n646) );
  XOR2_X1 U728 ( .A(KEYINPUT85), .B(n646), .Z(n650) );
  NAND2_X1 U729 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U730 ( .A1(n650), .A2(n649), .ZN(G295) );
  XOR2_X1 U731 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n652) );
  NAND2_X1 U732 ( .A1(G2078), .A2(G2084), .ZN(n651) );
  XNOR2_X1 U733 ( .A(n652), .B(n651), .ZN(n653) );
  NAND2_X1 U734 ( .A1(G2090), .A2(n653), .ZN(n654) );
  XNOR2_X1 U735 ( .A(KEYINPUT21), .B(n654), .ZN(n655) );
  NAND2_X1 U736 ( .A1(n655), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U737 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U738 ( .A(KEYINPUT68), .B(G82), .Z(G220) );
  NOR2_X1 U739 ( .A1(G238), .A2(G236), .ZN(n656) );
  NAND2_X1 U740 ( .A1(G69), .A2(n656), .ZN(n657) );
  NOR2_X1 U741 ( .A1(n657), .A2(G237), .ZN(n658) );
  XNOR2_X1 U742 ( .A(n658), .B(KEYINPUT87), .ZN(n811) );
  NAND2_X1 U743 ( .A1(n811), .A2(G567), .ZN(n663) );
  NOR2_X1 U744 ( .A1(G220), .A2(G219), .ZN(n659) );
  XOR2_X1 U745 ( .A(KEYINPUT22), .B(n659), .Z(n660) );
  NOR2_X1 U746 ( .A1(G218), .A2(n660), .ZN(n661) );
  NAND2_X1 U747 ( .A1(G96), .A2(n661), .ZN(n810) );
  NAND2_X1 U748 ( .A1(n810), .A2(G2106), .ZN(n662) );
  NAND2_X1 U749 ( .A1(n663), .A2(n662), .ZN(n813) );
  NAND2_X1 U750 ( .A1(G483), .A2(G661), .ZN(n664) );
  NOR2_X1 U751 ( .A1(n813), .A2(n664), .ZN(n809) );
  NAND2_X1 U752 ( .A1(n809), .A2(G36), .ZN(G176) );
  NAND2_X1 U753 ( .A1(G138), .A2(n867), .ZN(n666) );
  NAND2_X1 U754 ( .A1(G102), .A2(n868), .ZN(n665) );
  NAND2_X1 U755 ( .A1(n666), .A2(n665), .ZN(n670) );
  NAND2_X1 U756 ( .A1(G126), .A2(n863), .ZN(n668) );
  NAND2_X1 U757 ( .A1(G114), .A2(n864), .ZN(n667) );
  NAND2_X1 U758 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U759 ( .A1(n670), .A2(n669), .ZN(G164) );
  INV_X1 U760 ( .A(G166), .ZN(G303) );
  XOR2_X1 U761 ( .A(G2078), .B(KEYINPUT25), .Z(n989) );
  NAND2_X1 U762 ( .A1(G160), .A2(G40), .ZN(n766) );
  INV_X1 U763 ( .A(n766), .ZN(n671) );
  NOR2_X1 U764 ( .A1(G164), .A2(G1384), .ZN(n767) );
  NOR2_X1 U765 ( .A1(n989), .A2(n711), .ZN(n673) );
  XNOR2_X1 U766 ( .A(G1961), .B(KEYINPUT92), .ZN(n972) );
  NOR2_X1 U767 ( .A1(n695), .A2(n972), .ZN(n672) );
  NOR2_X1 U768 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U769 ( .A(KEYINPUT93), .B(n674), .ZN(n706) );
  NOR2_X1 U770 ( .A1(G171), .A2(n706), .ZN(n680) );
  NOR2_X1 U771 ( .A1(G1966), .A2(n748), .ZN(n724) );
  NOR2_X1 U772 ( .A1(G2084), .A2(n711), .ZN(n720) );
  NOR2_X1 U773 ( .A1(n724), .A2(n720), .ZN(n675) );
  NAND2_X1 U774 ( .A1(G8), .A2(n675), .ZN(n677) );
  INV_X1 U775 ( .A(G168), .ZN(n678) );
  NOR2_X1 U776 ( .A1(n680), .A2(n511), .ZN(n682) );
  XOR2_X1 U777 ( .A(KEYINPUT31), .B(KEYINPUT96), .Z(n681) );
  XNOR2_X1 U778 ( .A(n682), .B(n681), .ZN(n710) );
  XNOR2_X1 U779 ( .A(G1996), .B(KEYINPUT94), .ZN(n988) );
  NAND2_X1 U780 ( .A1(n988), .A2(n695), .ZN(n683) );
  XNOR2_X1 U781 ( .A(n683), .B(KEYINPUT26), .ZN(n686) );
  AND2_X1 U782 ( .A1(n711), .A2(G1341), .ZN(n684) );
  NOR2_X1 U783 ( .A1(n684), .A2(n922), .ZN(n685) );
  AND2_X1 U784 ( .A1(n686), .A2(n685), .ZN(n690) );
  NAND2_X1 U785 ( .A1(G1348), .A2(n711), .ZN(n688) );
  NAND2_X1 U786 ( .A1(G2067), .A2(n695), .ZN(n687) );
  NAND2_X1 U787 ( .A1(n688), .A2(n687), .ZN(n691) );
  NOR2_X1 U788 ( .A1(n692), .A2(n691), .ZN(n689) );
  AND2_X1 U789 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U790 ( .A1(n694), .A2(n693), .ZN(n700) );
  NAND2_X1 U791 ( .A1(n695), .A2(G2072), .ZN(n696) );
  XOR2_X1 U792 ( .A(n696), .B(KEYINPUT27), .Z(n698) );
  NAND2_X1 U793 ( .A1(G1956), .A2(n711), .ZN(n697) );
  NAND2_X1 U794 ( .A1(n698), .A2(n697), .ZN(n701) );
  NOR2_X1 U795 ( .A1(G299), .A2(n701), .ZN(n699) );
  OR2_X1 U796 ( .A1(n700), .A2(n699), .ZN(n704) );
  NAND2_X1 U797 ( .A1(G299), .A2(n701), .ZN(n702) );
  XNOR2_X1 U798 ( .A(KEYINPUT28), .B(n702), .ZN(n703) );
  AND2_X1 U799 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U800 ( .A(n705), .B(KEYINPUT29), .ZN(n708) );
  NAND2_X1 U801 ( .A1(G171), .A2(n706), .ZN(n707) );
  NAND2_X1 U802 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n722) );
  NAND2_X1 U804 ( .A1(n722), .A2(G286), .ZN(n716) );
  NOR2_X1 U805 ( .A1(G1971), .A2(n748), .ZN(n713) );
  NOR2_X1 U806 ( .A1(G2090), .A2(n711), .ZN(n712) );
  NOR2_X1 U807 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U808 ( .A1(n714), .A2(G303), .ZN(n715) );
  NAND2_X1 U809 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U810 ( .A(n717), .B(KEYINPUT98), .ZN(n718) );
  NAND2_X1 U811 ( .A1(n718), .A2(G8), .ZN(n719) );
  XNOR2_X1 U812 ( .A(KEYINPUT32), .B(n719), .ZN(n727) );
  NAND2_X1 U813 ( .A1(G8), .A2(n720), .ZN(n721) );
  NAND2_X1 U814 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U815 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U816 ( .A(KEYINPUT97), .B(n725), .ZN(n726) );
  NAND2_X1 U817 ( .A1(n727), .A2(n726), .ZN(n741) );
  NOR2_X1 U818 ( .A1(G1976), .A2(G288), .ZN(n734) );
  NOR2_X1 U819 ( .A1(G1971), .A2(G303), .ZN(n728) );
  NOR2_X1 U820 ( .A1(n734), .A2(n728), .ZN(n908) );
  NAND2_X1 U821 ( .A1(n741), .A2(n908), .ZN(n729) );
  XNOR2_X1 U822 ( .A(KEYINPUT99), .B(n729), .ZN(n732) );
  NAND2_X1 U823 ( .A1(G1976), .A2(G288), .ZN(n906) );
  INV_X1 U824 ( .A(n906), .ZN(n730) );
  OR2_X1 U825 ( .A1(n748), .A2(n730), .ZN(n731) );
  NOR2_X1 U826 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U827 ( .A1(n733), .A2(KEYINPUT33), .ZN(n737) );
  NAND2_X1 U828 ( .A1(n734), .A2(KEYINPUT33), .ZN(n735) );
  NOR2_X1 U829 ( .A1(n735), .A2(n748), .ZN(n736) );
  NOR2_X1 U830 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U831 ( .A(G1981), .B(G305), .Z(n916) );
  NAND2_X1 U832 ( .A1(n738), .A2(n916), .ZN(n745) );
  NOR2_X1 U833 ( .A1(G2090), .A2(G303), .ZN(n739) );
  NAND2_X1 U834 ( .A1(G8), .A2(n739), .ZN(n740) );
  NAND2_X1 U835 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U836 ( .A1(n748), .A2(n742), .ZN(n743) );
  XNOR2_X1 U837 ( .A(n743), .B(KEYINPUT100), .ZN(n744) );
  NAND2_X1 U838 ( .A1(n745), .A2(n744), .ZN(n793) );
  NOR2_X1 U839 ( .A1(G1981), .A2(G305), .ZN(n746) );
  XNOR2_X1 U840 ( .A(n746), .B(KEYINPUT91), .ZN(n747) );
  XNOR2_X1 U841 ( .A(n747), .B(KEYINPUT24), .ZN(n749) );
  NOR2_X1 U842 ( .A1(n749), .A2(n748), .ZN(n791) );
  NAND2_X1 U843 ( .A1(G105), .A2(n868), .ZN(n750) );
  XNOR2_X1 U844 ( .A(n750), .B(KEYINPUT38), .ZN(n757) );
  NAND2_X1 U845 ( .A1(G141), .A2(n867), .ZN(n752) );
  NAND2_X1 U846 ( .A1(G129), .A2(n863), .ZN(n751) );
  NAND2_X1 U847 ( .A1(n752), .A2(n751), .ZN(n755) );
  NAND2_X1 U848 ( .A1(n864), .A2(G117), .ZN(n753) );
  XOR2_X1 U849 ( .A(KEYINPUT90), .B(n753), .Z(n754) );
  NOR2_X1 U850 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U851 ( .A1(n757), .A2(n756), .ZN(n842) );
  NOR2_X1 U852 ( .A1(G1996), .A2(n842), .ZN(n942) );
  NAND2_X1 U853 ( .A1(G131), .A2(n867), .ZN(n759) );
  NAND2_X1 U854 ( .A1(G119), .A2(n863), .ZN(n758) );
  NAND2_X1 U855 ( .A1(n759), .A2(n758), .ZN(n763) );
  NAND2_X1 U856 ( .A1(G95), .A2(n868), .ZN(n761) );
  NAND2_X1 U857 ( .A1(G107), .A2(n864), .ZN(n760) );
  NAND2_X1 U858 ( .A1(n761), .A2(n760), .ZN(n762) );
  OR2_X1 U859 ( .A1(n763), .A2(n762), .ZN(n841) );
  AND2_X1 U860 ( .A1(n841), .A2(G1991), .ZN(n765) );
  AND2_X1 U861 ( .A1(n842), .A2(G1996), .ZN(n764) );
  NOR2_X1 U862 ( .A1(n765), .A2(n764), .ZN(n928) );
  NOR2_X1 U863 ( .A1(n767), .A2(n766), .ZN(n794) );
  INV_X1 U864 ( .A(n794), .ZN(n768) );
  NOR2_X1 U865 ( .A1(n928), .A2(n768), .ZN(n795) );
  NOR2_X1 U866 ( .A1(G1991), .A2(n841), .ZN(n931) );
  NOR2_X1 U867 ( .A1(G1986), .A2(G290), .ZN(n769) );
  NOR2_X1 U868 ( .A1(n931), .A2(n769), .ZN(n770) );
  NOR2_X1 U869 ( .A1(n795), .A2(n770), .ZN(n771) );
  NOR2_X1 U870 ( .A1(n942), .A2(n771), .ZN(n772) );
  XOR2_X1 U871 ( .A(n772), .B(KEYINPUT39), .Z(n773) );
  XNOR2_X1 U872 ( .A(KEYINPUT101), .B(n773), .ZN(n785) );
  XNOR2_X1 U873 ( .A(KEYINPUT37), .B(G2067), .ZN(n787) );
  NAND2_X1 U874 ( .A1(G128), .A2(n863), .ZN(n775) );
  NAND2_X1 U875 ( .A1(G116), .A2(n864), .ZN(n774) );
  NAND2_X1 U876 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U877 ( .A(KEYINPUT35), .B(n776), .ZN(n782) );
  NAND2_X1 U878 ( .A1(n868), .A2(G104), .ZN(n777) );
  XNOR2_X1 U879 ( .A(n777), .B(KEYINPUT88), .ZN(n779) );
  NAND2_X1 U880 ( .A1(G140), .A2(n867), .ZN(n778) );
  NAND2_X1 U881 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U882 ( .A(KEYINPUT34), .B(n780), .Z(n781) );
  NAND2_X1 U883 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U884 ( .A(KEYINPUT36), .B(n783), .Z(n852) );
  OR2_X1 U885 ( .A1(n787), .A2(n852), .ZN(n784) );
  XNOR2_X1 U886 ( .A(KEYINPUT89), .B(n784), .ZN(n949) );
  NAND2_X1 U887 ( .A1(n794), .A2(n949), .ZN(n796) );
  NAND2_X1 U888 ( .A1(n785), .A2(n796), .ZN(n786) );
  XNOR2_X1 U889 ( .A(n786), .B(KEYINPUT102), .ZN(n788) );
  NAND2_X1 U890 ( .A1(n787), .A2(n852), .ZN(n927) );
  NAND2_X1 U891 ( .A1(n788), .A2(n927), .ZN(n789) );
  NAND2_X1 U892 ( .A1(n789), .A2(n794), .ZN(n801) );
  INV_X1 U893 ( .A(n801), .ZN(n790) );
  OR2_X1 U894 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U895 ( .A1(n793), .A2(n792), .ZN(n803) );
  XNOR2_X1 U896 ( .A(G1986), .B(G290), .ZN(n914) );
  AND2_X1 U897 ( .A1(n914), .A2(n794), .ZN(n799) );
  INV_X1 U898 ( .A(n795), .ZN(n797) );
  NAND2_X1 U899 ( .A1(n797), .A2(n796), .ZN(n798) );
  OR2_X1 U900 ( .A1(n799), .A2(n798), .ZN(n800) );
  AND2_X1 U901 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U902 ( .A(n804), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U903 ( .A1(n805), .A2(G2106), .ZN(n806) );
  XOR2_X1 U904 ( .A(KEYINPUT105), .B(n806), .Z(G217) );
  AND2_X1 U905 ( .A1(G15), .A2(G2), .ZN(n807) );
  NAND2_X1 U906 ( .A1(G661), .A2(n807), .ZN(G259) );
  NAND2_X1 U907 ( .A1(G3), .A2(G1), .ZN(n808) );
  NAND2_X1 U908 ( .A1(n809), .A2(n808), .ZN(G188) );
  XOR2_X1 U909 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  XNOR2_X1 U910 ( .A(G69), .B(KEYINPUT107), .ZN(G235) );
  NOR2_X1 U912 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U913 ( .A(n812), .B(KEYINPUT108), .ZN(G325) );
  INV_X1 U914 ( .A(G325), .ZN(G261) );
  INV_X1 U915 ( .A(n813), .ZN(G319) );
  XNOR2_X1 U916 ( .A(G1981), .B(G2474), .ZN(n823) );
  XOR2_X1 U917 ( .A(G1956), .B(G1961), .Z(n815) );
  XNOR2_X1 U918 ( .A(G1986), .B(G1966), .ZN(n814) );
  XNOR2_X1 U919 ( .A(n815), .B(n814), .ZN(n819) );
  XOR2_X1 U920 ( .A(G1971), .B(G1976), .Z(n817) );
  XNOR2_X1 U921 ( .A(G1996), .B(G1991), .ZN(n816) );
  XNOR2_X1 U922 ( .A(n817), .B(n816), .ZN(n818) );
  XOR2_X1 U923 ( .A(n819), .B(n818), .Z(n821) );
  XNOR2_X1 U924 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n820) );
  XNOR2_X1 U925 ( .A(n821), .B(n820), .ZN(n822) );
  XNOR2_X1 U926 ( .A(n823), .B(n822), .ZN(G229) );
  XOR2_X1 U927 ( .A(G2678), .B(G2090), .Z(n825) );
  XNOR2_X1 U928 ( .A(G2084), .B(G2078), .ZN(n824) );
  XNOR2_X1 U929 ( .A(n825), .B(n824), .ZN(n826) );
  XOR2_X1 U930 ( .A(n826), .B(G2096), .Z(n828) );
  XNOR2_X1 U931 ( .A(G2067), .B(G2072), .ZN(n827) );
  XNOR2_X1 U932 ( .A(n828), .B(n827), .ZN(n832) );
  XOR2_X1 U933 ( .A(G2100), .B(KEYINPUT109), .Z(n830) );
  XNOR2_X1 U934 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n829) );
  XNOR2_X1 U935 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U936 ( .A(n832), .B(n831), .Z(G227) );
  NAND2_X1 U937 ( .A1(G100), .A2(n868), .ZN(n834) );
  NAND2_X1 U938 ( .A1(G112), .A2(n864), .ZN(n833) );
  NAND2_X1 U939 ( .A1(n834), .A2(n833), .ZN(n840) );
  NAND2_X1 U940 ( .A1(n863), .A2(G124), .ZN(n835) );
  XNOR2_X1 U941 ( .A(n835), .B(KEYINPUT44), .ZN(n837) );
  NAND2_X1 U942 ( .A1(G136), .A2(n867), .ZN(n836) );
  NAND2_X1 U943 ( .A1(n837), .A2(n836), .ZN(n838) );
  XOR2_X1 U944 ( .A(KEYINPUT111), .B(n838), .Z(n839) );
  NOR2_X1 U945 ( .A1(n840), .A2(n839), .ZN(G162) );
  XNOR2_X1 U946 ( .A(G162), .B(n841), .ZN(n844) );
  XOR2_X1 U947 ( .A(G164), .B(n842), .Z(n843) );
  XNOR2_X1 U948 ( .A(n844), .B(n843), .ZN(n851) );
  XOR2_X1 U949 ( .A(KEYINPUT114), .B(KEYINPUT112), .Z(n846) );
  XNOR2_X1 U950 ( .A(KEYINPUT46), .B(KEYINPUT115), .ZN(n845) );
  XNOR2_X1 U951 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U952 ( .A(n847), .B(KEYINPUT116), .Z(n849) );
  XNOR2_X1 U953 ( .A(n930), .B(KEYINPUT48), .ZN(n848) );
  XNOR2_X1 U954 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U955 ( .A(n851), .B(n850), .Z(n854) );
  XOR2_X1 U956 ( .A(G160), .B(n852), .Z(n853) );
  XNOR2_X1 U957 ( .A(n854), .B(n853), .ZN(n876) );
  NAND2_X1 U958 ( .A1(G139), .A2(n867), .ZN(n856) );
  NAND2_X1 U959 ( .A1(G103), .A2(n868), .ZN(n855) );
  NAND2_X1 U960 ( .A1(n856), .A2(n855), .ZN(n862) );
  NAND2_X1 U961 ( .A1(n863), .A2(G127), .ZN(n857) );
  XOR2_X1 U962 ( .A(KEYINPUT113), .B(n857), .Z(n859) );
  NAND2_X1 U963 ( .A1(n864), .A2(G115), .ZN(n858) );
  NAND2_X1 U964 ( .A1(n859), .A2(n858), .ZN(n860) );
  XOR2_X1 U965 ( .A(KEYINPUT47), .B(n860), .Z(n861) );
  NOR2_X1 U966 ( .A1(n862), .A2(n861), .ZN(n937) );
  NAND2_X1 U967 ( .A1(G130), .A2(n863), .ZN(n866) );
  NAND2_X1 U968 ( .A1(G118), .A2(n864), .ZN(n865) );
  NAND2_X1 U969 ( .A1(n866), .A2(n865), .ZN(n873) );
  NAND2_X1 U970 ( .A1(G142), .A2(n867), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G106), .A2(n868), .ZN(n869) );
  NAND2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U973 ( .A(KEYINPUT45), .B(n871), .Z(n872) );
  NOR2_X1 U974 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n937), .B(n874), .ZN(n875) );
  XNOR2_X1 U976 ( .A(n876), .B(n875), .ZN(n877) );
  NOR2_X1 U977 ( .A1(G37), .A2(n877), .ZN(G395) );
  XNOR2_X1 U978 ( .A(n901), .B(G286), .ZN(n881) );
  XOR2_X1 U979 ( .A(G171), .B(n878), .Z(n879) );
  XNOR2_X1 U980 ( .A(n922), .B(n879), .ZN(n880) );
  XNOR2_X1 U981 ( .A(n881), .B(n880), .ZN(n882) );
  NOR2_X1 U982 ( .A1(G37), .A2(n882), .ZN(G397) );
  XNOR2_X1 U983 ( .A(G2454), .B(G2446), .ZN(n892) );
  XOR2_X1 U984 ( .A(KEYINPUT104), .B(G2430), .Z(n884) );
  XNOR2_X1 U985 ( .A(G2451), .B(G2443), .ZN(n883) );
  XNOR2_X1 U986 ( .A(n884), .B(n883), .ZN(n888) );
  XOR2_X1 U987 ( .A(G2427), .B(KEYINPUT103), .Z(n886) );
  XNOR2_X1 U988 ( .A(G1341), .B(G1348), .ZN(n885) );
  XNOR2_X1 U989 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U990 ( .A(n888), .B(n887), .Z(n890) );
  XNOR2_X1 U991 ( .A(G2435), .B(G2438), .ZN(n889) );
  XNOR2_X1 U992 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U993 ( .A(n892), .B(n891), .ZN(n893) );
  NAND2_X1 U994 ( .A1(n893), .A2(G14), .ZN(n900) );
  NAND2_X1 U995 ( .A1(G319), .A2(n900), .ZN(n897) );
  NOR2_X1 U996 ( .A1(G229), .A2(G227), .ZN(n894) );
  XOR2_X1 U997 ( .A(KEYINPUT117), .B(n894), .Z(n895) );
  XNOR2_X1 U998 ( .A(n895), .B(KEYINPUT49), .ZN(n896) );
  NOR2_X1 U999 ( .A1(n897), .A2(n896), .ZN(n899) );
  NOR2_X1 U1000 ( .A1(G395), .A2(G397), .ZN(n898) );
  NAND2_X1 U1001 ( .A1(n899), .A2(n898), .ZN(G225) );
  INV_X1 U1002 ( .A(G225), .ZN(G308) );
  INV_X1 U1003 ( .A(n900), .ZN(G401) );
  XNOR2_X1 U1004 ( .A(n901), .B(G1348), .ZN(n903) );
  XNOR2_X1 U1005 ( .A(G171), .B(G1961), .ZN(n902) );
  NAND2_X1 U1006 ( .A1(n903), .A2(n902), .ZN(n904) );
  XNOR2_X1 U1007 ( .A(KEYINPUT123), .B(n904), .ZN(n912) );
  NAND2_X1 U1008 ( .A1(G1971), .A2(G303), .ZN(n905) );
  NAND2_X1 U1009 ( .A1(n906), .A2(n905), .ZN(n910) );
  XOR2_X1 U1010 ( .A(G1956), .B(G299), .Z(n907) );
  NAND2_X1 U1011 ( .A1(n908), .A2(n907), .ZN(n909) );
  NOR2_X1 U1012 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1013 ( .A1(n912), .A2(n911), .ZN(n913) );
  NOR2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n915) );
  XNOR2_X1 U1015 ( .A(KEYINPUT124), .B(n915), .ZN(n921) );
  XNOR2_X1 U1016 ( .A(G1966), .B(G168), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(n918), .B(KEYINPUT57), .ZN(n919) );
  XNOR2_X1 U1019 ( .A(KEYINPUT122), .B(n919), .ZN(n920) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n924) );
  XNOR2_X1 U1021 ( .A(G1341), .B(n922), .ZN(n923) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n926) );
  XOR2_X1 U1023 ( .A(KEYINPUT56), .B(G16), .Z(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n956) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n936) );
  XNOR2_X1 U1026 ( .A(G2084), .B(G160), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(n929), .B(KEYINPUT118), .ZN(n933) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1030 ( .A(KEYINPUT119), .B(n934), .Z(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n947) );
  XOR2_X1 U1032 ( .A(G2072), .B(n937), .Z(n939) );
  XOR2_X1 U1033 ( .A(G164), .B(G2078), .Z(n938) );
  NOR2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1035 ( .A(KEYINPUT50), .B(n940), .Z(n945) );
  XOR2_X1 U1036 ( .A(G2090), .B(G162), .Z(n941) );
  NOR2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(KEYINPUT51), .B(n943), .ZN(n944) );
  NOR2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(n950), .B(KEYINPUT52), .ZN(n952) );
  INV_X1 U1043 ( .A(KEYINPUT55), .ZN(n951) );
  NAND2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1045 ( .A1(G29), .A2(n953), .ZN(n954) );
  XOR2_X1 U1046 ( .A(KEYINPUT120), .B(n954), .Z(n955) );
  NOR2_X1 U1047 ( .A1(n956), .A2(n955), .ZN(n1005) );
  XNOR2_X1 U1048 ( .A(G16), .B(KEYINPUT125), .ZN(n980) );
  XOR2_X1 U1049 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n978) );
  XOR2_X1 U1050 ( .A(G1348), .B(KEYINPUT59), .Z(n957) );
  XNOR2_X1 U1051 ( .A(G4), .B(n957), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(G19), .B(G1341), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(G1981), .B(G6), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(G1956), .B(G20), .ZN(n960) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(n964), .B(KEYINPUT60), .ZN(n971) );
  XNOR2_X1 U1059 ( .A(G1976), .B(G23), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(G1971), .B(G22), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n968) );
  XOR2_X1 U1062 ( .A(G1986), .B(G24), .Z(n967) );
  NAND2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(KEYINPUT58), .B(n969), .ZN(n970) );
  NOR2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(n972), .B(G5), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(G21), .B(G1966), .ZN(n973) );
  NOR2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(n978), .B(n977), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1072 ( .A1(n981), .A2(G11), .ZN(n1003) );
  XNOR2_X1 U1073 ( .A(G2067), .B(G26), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(G33), .B(G2072), .ZN(n982) );
  NOR2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1076 ( .A1(G28), .A2(n984), .ZN(n987) );
  XOR2_X1 U1077 ( .A(G25), .B(G1991), .Z(n985) );
  XNOR2_X1 U1078 ( .A(KEYINPUT121), .B(n985), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(n988), .B(G32), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(G27), .B(n989), .ZN(n990) );
  NOR2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(n994), .B(KEYINPUT53), .ZN(n997) );
  XOR2_X1 U1085 ( .A(G2084), .B(G34), .Z(n995) );
  XNOR2_X1 U1086 ( .A(KEYINPUT54), .B(n995), .ZN(n996) );
  NAND2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(G35), .B(G2090), .ZN(n998) );
  NOR2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1090 ( .A(KEYINPUT55), .B(n1000), .Z(n1001) );
  NOR2_X1 U1091 ( .A1(G29), .A2(n1001), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(KEYINPUT62), .B(n1006), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(KEYINPUT127), .B(n1007), .ZN(G311) );
  INV_X1 U1096 ( .A(G311), .ZN(G150) );
endmodule

