//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n543,
    new_n544, new_n546, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n458), .B1(KEYINPUT67), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n461), .B1(KEYINPUT67), .B2(new_n460), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT68), .Z(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n466), .A2(new_n468), .A3(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(G101), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n466), .A2(new_n468), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n464), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n476), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(new_n464), .B2(G112), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n478), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND4_X1  g059(.A1(new_n466), .A2(new_n468), .A3(G138), .A4(new_n464), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g062(.A(KEYINPUT3), .B(G2104), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n488), .A2(KEYINPUT4), .A3(G138), .A4(new_n464), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n488), .A2(G126), .A3(G2105), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n492));
  OAI21_X1  g067(.A(G2105), .B1(new_n492), .B2(G114), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(KEYINPUT69), .ZN(new_n495));
  OAI211_X1 g070(.A(G2104), .B(new_n491), .C1(new_n493), .C2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n487), .A2(new_n489), .A3(new_n490), .A4(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  NAND2_X1  g073(.A1(G75), .A2(G543), .ZN(new_n499));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G62), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n499), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G651), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(G50), .A3(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n511));
  XOR2_X1   g086(.A(KEYINPUT6), .B(G651), .Z(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(new_n504), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n501), .A2(new_n503), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(new_n508), .A3(KEYINPUT70), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n510), .B1(new_n516), .B2(G88), .ZN(G166));
  NAND2_X1  g092(.A1(new_n512), .A2(KEYINPUT71), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n508), .A2(new_n519), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n518), .A2(G543), .A3(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n514), .A2(G63), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n521), .A2(G51), .B1(G651), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n516), .A2(G89), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(G286));
  INV_X1    g102(.A(G286), .ZN(G168));
  XNOR2_X1  g103(.A(KEYINPUT72), .B(G52), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n521), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G651), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n513), .A2(new_n515), .A3(G90), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n530), .A2(new_n533), .A3(new_n534), .ZN(G171));
  NAND3_X1  g110(.A1(new_n518), .A2(G543), .A3(new_n520), .ZN(new_n536));
  INV_X1    g111(.A(G43), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n536), .A2(new_n537), .B1(new_n532), .B2(new_n538), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n513), .A2(new_n515), .A3(G81), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  NAND3_X1  g117(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G36), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT73), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n544), .A2(new_n548), .ZN(G188));
  INV_X1    g124(.A(KEYINPUT9), .ZN(new_n550));
  INV_X1    g125(.A(G53), .ZN(new_n551));
  OAI211_X1 g126(.A(KEYINPUT74), .B(new_n550), .C1(new_n536), .C2(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n513), .A2(new_n515), .A3(G91), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n514), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n554), .A2(new_n532), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  OR3_X1    g131(.A1(new_n536), .A2(KEYINPUT74), .A3(new_n551), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT74), .B1(new_n536), .B2(new_n551), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n557), .A2(KEYINPUT9), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G299));
  NAND3_X1  g135(.A1(new_n530), .A2(new_n533), .A3(new_n534), .ZN(G301));
  INV_X1    g136(.A(G166), .ZN(G303));
  NAND2_X1  g137(.A1(new_n516), .A2(G87), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n521), .A2(G49), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(G288));
  NAND2_X1  g141(.A1(new_n516), .A2(G86), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n508), .A2(G48), .A3(G543), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT77), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n568), .B(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n514), .A2(KEYINPUT75), .A3(G61), .ZN(new_n571));
  NAND2_X1  g146(.A1(G73), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n504), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n571), .A2(new_n572), .A3(new_n575), .ZN(new_n576));
  AND3_X1   g151(.A1(new_n576), .A2(KEYINPUT76), .A3(G651), .ZN(new_n577));
  AOI21_X1  g152(.A(KEYINPUT76), .B1(new_n576), .B2(G651), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n567), .B(new_n570), .C1(new_n577), .C2(new_n578), .ZN(G305));
  NAND2_X1  g154(.A1(new_n516), .A2(G85), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n581), .A2(new_n532), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n521), .A2(G47), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  XOR2_X1   g160(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n586));
  NAND3_X1  g161(.A1(new_n516), .A2(G92), .A3(new_n586), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n514), .A2(G66), .ZN(new_n588));
  NAND2_X1  g163(.A1(G79), .A2(G543), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT79), .Z(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n586), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n513), .A2(new_n515), .ZN(new_n593));
  INV_X1    g168(.A(G92), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n521), .A2(G54), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n587), .A2(new_n591), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n585), .B1(new_n598), .B2(G868), .ZN(G321));
  XNOR2_X1  g174(.A(G321), .B(KEYINPUT80), .ZN(G284));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(G299), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(new_n601), .B2(G168), .ZN(G297));
  OAI21_X1  g178(.A(new_n602), .B1(new_n601), .B2(G168), .ZN(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n598), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND2_X1  g181(.A1(new_n598), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G868), .B2(new_n541), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g185(.A1(new_n464), .A2(G111), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n465), .B1(new_n611), .B2(KEYINPUT82), .ZN(new_n612));
  OAI221_X1 g187(.A(new_n612), .B1(KEYINPUT82), .B2(new_n611), .C1(G99), .C2(G2105), .ZN(new_n613));
  AOI22_X1  g188(.A1(G123), .A2(new_n477), .B1(new_n479), .B2(G135), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT83), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(G2096), .Z(new_n618));
  NAND2_X1  g193(.A1(new_n479), .A2(G2104), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT13), .B(G2100), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n618), .A2(new_n623), .ZN(G156));
  XNOR2_X1  g199(.A(G2427), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2430), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT15), .B(G2435), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(KEYINPUT14), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT84), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n629), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n635), .B(new_n636), .Z(new_n637));
  AND2_X1   g212(.A1(new_n637), .A2(G14), .ZN(G401));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2067), .B(G2678), .Z(new_n641));
  NOR2_X1   g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n640), .A2(new_n641), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(new_n644), .A3(KEYINPUT17), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT18), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2072), .B(G2078), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n647), .B(new_n648), .C1(new_n646), .C2(new_n642), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(new_n648), .B2(new_n647), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2096), .B(G2100), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(G227));
  XOR2_X1   g227(.A(G1971), .B(G1976), .Z(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  XOR2_X1   g231(.A(G1961), .B(G1966), .Z(new_n657));
  AND2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g233(.A(KEYINPUT20), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n655), .A2(KEYINPUT20), .A3(new_n658), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n660), .B1(new_n655), .B2(new_n662), .ZN(new_n663));
  AOI211_X1 g238(.A(new_n659), .B(new_n663), .C1(new_n661), .C2(new_n655), .ZN(new_n664));
  XOR2_X1   g239(.A(G1986), .B(G1996), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G1981), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G1991), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n666), .B(new_n669), .ZN(G229));
  AOI22_X1  g245(.A1(new_n488), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT93), .ZN(new_n672));
  AOI22_X1  g247(.A1(new_n672), .A2(G2105), .B1(G139), .B2(new_n479), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT25), .Z(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  MUX2_X1   g251(.A(G33), .B(new_n676), .S(G29), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2072), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n679));
  INV_X1    g254(.A(G29), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G26), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n477), .A2(G128), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n479), .A2(G140), .ZN(new_n684));
  NOR2_X1   g259(.A1(G104), .A2(G2105), .ZN(new_n685));
  OAI21_X1  g260(.A(G2104), .B1(new_n464), .B2(G116), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n683), .B(new_n684), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  AND3_X1   g262(.A1(new_n687), .A2(KEYINPUT91), .A3(G29), .ZN(new_n688));
  AOI21_X1  g263(.A(KEYINPUT91), .B1(new_n687), .B2(G29), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n682), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G2067), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n680), .A2(G27), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G164), .B2(new_n680), .ZN(new_n693));
  MUX2_X1   g268(.A(new_n692), .B(new_n693), .S(KEYINPUT95), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G2078), .ZN(new_n695));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G4), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(new_n598), .B2(new_n696), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT90), .Z(new_n699));
  AOI211_X1 g274(.A(new_n691), .B(new_n695), .C1(new_n699), .C2(G1348), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n699), .A2(G1348), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n696), .A2(G20), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT97), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT23), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G299), .B2(G16), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1956), .ZN(new_n707));
  INV_X1    g282(.A(G2090), .ZN(new_n708));
  INV_X1    g283(.A(G35), .ZN(new_n709));
  OAI21_X1  g284(.A(KEYINPUT96), .B1(new_n709), .B2(G29), .ZN(new_n710));
  OR3_X1    g285(.A1(new_n709), .A2(KEYINPUT96), .A3(G29), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n710), .B(new_n711), .C1(G162), .C2(new_n680), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT29), .Z(new_n713));
  OAI21_X1  g288(.A(new_n707), .B1(new_n708), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT98), .ZN(new_n715));
  OR2_X1    g290(.A1(KEYINPUT24), .A2(G34), .ZN(new_n716));
  NAND2_X1  g291(.A1(KEYINPUT24), .A2(G34), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n716), .A2(new_n680), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G160), .B2(new_n680), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(G2084), .ZN(new_n720));
  OR2_X1    g295(.A1(G29), .A2(G32), .ZN(new_n721));
  AOI22_X1  g296(.A1(G129), .A2(new_n477), .B1(new_n479), .B2(G141), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n723));
  NAND3_X1  g298(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT26), .Z(new_n725));
  NAND3_X1  g300(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n721), .B1(new_n726), .B2(new_n680), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT27), .B(G1996), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n617), .A2(new_n680), .ZN(new_n730));
  AOI211_X1 g305(.A(new_n729), .B(new_n730), .C1(G2084), .C2(new_n719), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n713), .A2(new_n708), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n696), .A2(G19), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n541), .B2(new_n696), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G1341), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n727), .A2(new_n728), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT31), .B(G11), .ZN(new_n737));
  INV_X1    g312(.A(G28), .ZN(new_n738));
  AOI21_X1  g313(.A(G29), .B1(new_n738), .B2(KEYINPUT30), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(KEYINPUT30), .B2(new_n738), .ZN(new_n740));
  AND3_X1   g315(.A1(new_n736), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n731), .A2(new_n732), .A3(new_n735), .A4(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(G16), .A2(G21), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G286), .B2(new_n696), .ZN(new_n744));
  INV_X1    g319(.A(G1966), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT94), .ZN(new_n747));
  NAND2_X1  g322(.A1(G171), .A2(G16), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G5), .B2(G16), .ZN(new_n749));
  INV_X1    g324(.A(G1961), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n744), .A2(new_n745), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n752), .B(new_n753), .C1(G1341), .C2(new_n734), .ZN(new_n754));
  NOR4_X1   g329(.A1(new_n742), .A2(new_n747), .A3(new_n751), .A4(new_n754), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n702), .A2(new_n715), .A3(new_n720), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n696), .A2(G6), .ZN(new_n757));
  INV_X1    g332(.A(G305), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(new_n696), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT89), .Z(new_n760));
  XOR2_X1   g335(.A(KEYINPUT32), .B(G1981), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G1976), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n696), .A2(G23), .ZN(new_n764));
  AND3_X1   g339(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(new_n696), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(KEYINPUT33), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n766), .A2(KEYINPUT33), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n763), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n769), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n771), .A2(G1976), .A3(new_n767), .ZN(new_n772));
  NOR2_X1   g347(.A1(G166), .A2(new_n696), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n696), .B2(G22), .ZN(new_n774));
  INV_X1    g349(.A(G1971), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AND3_X1   g351(.A1(new_n770), .A2(new_n772), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n774), .A2(new_n775), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n759), .B(KEYINPUT89), .ZN(new_n779));
  INV_X1    g354(.A(new_n761), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n762), .A2(new_n777), .A3(new_n778), .A4(new_n781), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT88), .B(KEYINPUT34), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT36), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n477), .A2(G119), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n479), .A2(G131), .ZN(new_n787));
  OR2_X1    g362(.A1(G95), .A2(G2105), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n788), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  MUX2_X1   g365(.A(G25), .B(new_n790), .S(G29), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT86), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT35), .B(G1991), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n696), .A2(G24), .ZN(new_n795));
  INV_X1    g370(.A(G290), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(new_n796), .B2(new_n696), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT87), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1986), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n784), .A2(new_n785), .A3(new_n794), .A4(new_n799), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n762), .A2(new_n777), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n801), .A2(new_n783), .A3(new_n778), .A4(new_n781), .ZN(new_n802));
  INV_X1    g377(.A(new_n783), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n782), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n802), .A2(new_n794), .A3(new_n804), .A4(new_n799), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(KEYINPUT36), .ZN(new_n806));
  AOI211_X1 g381(.A(new_n678), .B(new_n756), .C1(new_n800), .C2(new_n806), .ZN(G311));
  AOI21_X1  g382(.A(new_n756), .B1(new_n800), .B2(new_n806), .ZN(new_n808));
  INV_X1    g383(.A(new_n678), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(G150));
  NAND2_X1  g385(.A1(G80), .A2(G543), .ZN(new_n811));
  INV_X1    g386(.A(G67), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n504), .B2(new_n812), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n521), .A2(G55), .B1(G651), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n516), .A2(G93), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G860), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT37), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n598), .A2(G559), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT38), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n816), .A2(new_n541), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n814), .B(new_n815), .C1(new_n540), .C2(new_n539), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT39), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n820), .B(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n818), .B1(new_n825), .B2(G860), .ZN(G145));
  INV_X1    g401(.A(G37), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n726), .B(new_n687), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G164), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n673), .A2(KEYINPUT100), .A3(new_n675), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT100), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n676), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n828), .B(new_n497), .ZN(new_n834));
  INV_X1    g409(.A(new_n830), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n477), .A2(G130), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n479), .A2(G142), .ZN(new_n839));
  NOR2_X1   g414(.A1(G106), .A2(G2105), .ZN(new_n840));
  OAI21_X1  g415(.A(G2104), .B1(new_n464), .B2(G118), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n838), .B(new_n839), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n790), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n621), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT101), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n837), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(G160), .B(KEYINPUT99), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G162), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n617), .ZN(new_n849));
  INV_X1    g424(.A(new_n844), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n846), .B(new_n849), .C1(new_n837), .C2(new_n850), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n837), .A2(new_n845), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n852), .A2(KEYINPUT102), .A3(new_n846), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT102), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n837), .A2(new_n854), .A3(new_n845), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n827), .B(new_n851), .C1(new_n856), .C2(new_n849), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g433(.A1(new_n816), .A2(new_n601), .ZN(new_n859));
  NAND2_X1  g434(.A1(G299), .A2(new_n598), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n556), .A2(new_n597), .A3(new_n559), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(KEYINPUT103), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n863));
  NAND3_X1  g438(.A1(G299), .A2(new_n598), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT41), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n860), .A2(new_n861), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT104), .B1(new_n867), .B2(KEYINPUT41), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n860), .A2(new_n861), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT104), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT41), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n866), .A2(new_n868), .A3(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n607), .B(new_n823), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n865), .ZN(new_n876));
  OAI21_X1  g451(.A(KEYINPUT105), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(KEYINPUT105), .B2(new_n875), .ZN(new_n878));
  NAND2_X1  g453(.A1(G288), .A2(G166), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(G288), .A2(G166), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n880), .A2(new_n796), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n765), .A2(G303), .ZN(new_n883));
  AOI21_X1  g458(.A(G290), .B1(new_n883), .B2(new_n879), .ZN(new_n884));
  OAI21_X1  g459(.A(G305), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n796), .B1(new_n880), .B2(new_n881), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(new_n879), .A3(G290), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n886), .A2(new_n758), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT42), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n878), .B(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n859), .B1(new_n891), .B2(new_n601), .ZN(G295));
  OAI21_X1  g467(.A(new_n859), .B1(new_n891), .B2(new_n601), .ZN(G331));
  NAND2_X1  g468(.A1(G286), .A2(G171), .ZN(new_n894));
  NAND4_X1  g469(.A1(G301), .A2(new_n525), .A3(new_n526), .A4(new_n523), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n823), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT106), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT106), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n896), .B2(new_n823), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n896), .A2(new_n823), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n865), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n871), .B1(new_n862), .B2(new_n864), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n870), .B1(new_n869), .B2(new_n871), .ZN(new_n907));
  AOI211_X1 g482(.A(KEYINPUT104), .B(KEYINPUT41), .C1(new_n860), .C2(new_n861), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n897), .A2(new_n898), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n902), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n905), .B(new_n889), .C1(new_n909), .C2(new_n912), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n873), .A2(new_n911), .B1(new_n904), .B2(new_n903), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n889), .B(new_n915), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n913), .B(new_n827), .C1(new_n914), .C2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(G37), .B1(new_n914), .B2(new_n889), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n889), .B(KEYINPUT107), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n911), .A2(new_n865), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n867), .A2(new_n871), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT41), .B1(new_n862), .B2(new_n864), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n903), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n921), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n920), .A2(KEYINPUT43), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT44), .B1(new_n919), .B2(new_n927), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n917), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT108), .B1(new_n917), .B2(KEYINPUT43), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n920), .A2(new_n918), .A3(new_n926), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n928), .B1(new_n932), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g508(.A1(new_n469), .A2(new_n470), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(G2105), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n472), .A2(new_n473), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n464), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n937), .A3(G40), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT110), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT110), .ZN(new_n940));
  NAND3_X1  g515(.A1(G160), .A2(new_n940), .A3(G40), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G1384), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n487), .A2(new_n489), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n490), .A2(new_n496), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  XOR2_X1   g521(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n942), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G1996), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n726), .B(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G2067), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n687), .B(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n790), .A2(new_n793), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n790), .A2(new_n793), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G1986), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n960), .B1(new_n961), .B2(new_n796), .ZN(new_n962));
  NOR2_X1   g537(.A1(G290), .A2(G1986), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n950), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n943), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n949), .A2(new_n939), .A3(new_n941), .A4(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G2078), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT53), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n946), .A2(KEYINPUT50), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n497), .A2(new_n972), .A3(new_n943), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n971), .A2(new_n939), .A3(new_n941), .A4(new_n973), .ZN(new_n974));
  AOI22_X1  g549(.A1(new_n969), .A2(new_n970), .B1(new_n750), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT116), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT45), .B1(new_n497), .B2(new_n943), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n976), .B1(new_n942), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n946), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n947), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n946), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n982), .A2(KEYINPUT116), .A3(new_n939), .A4(new_n941), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n978), .A2(new_n968), .A3(new_n980), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT121), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT53), .B1(new_n984), .B2(KEYINPUT121), .ZN(new_n987));
  OAI211_X1 g562(.A(G301), .B(new_n975), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT123), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT54), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n943), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n947), .B1(new_n497), .B2(new_n943), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n991), .A2(new_n992), .A3(new_n938), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n993), .A2(KEYINPUT53), .A3(new_n968), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT122), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n994), .B(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n975), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n990), .B1(new_n997), .B2(G171), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n940), .B1(G160), .B2(G40), .ZN(new_n999));
  INV_X1    g574(.A(G40), .ZN(new_n1000));
  NOR4_X1   g575(.A1(new_n471), .A2(new_n474), .A3(KEYINPUT110), .A4(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT116), .B1(new_n1002), .B2(new_n982), .ZN(new_n1003));
  AND4_X1   g578(.A1(KEYINPUT116), .A2(new_n982), .A3(new_n939), .A4(new_n941), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT121), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1005), .A2(new_n1006), .A3(new_n968), .A4(new_n980), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1007), .A2(KEYINPUT53), .A3(new_n985), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT123), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1008), .A2(new_n1009), .A3(G301), .A4(new_n975), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n989), .A2(new_n998), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(G301), .B1(new_n1008), .B2(new_n975), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n997), .A2(G171), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n990), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n942), .A2(new_n946), .ZN(new_n1015));
  INV_X1    g590(.A(G8), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(G288), .A2(new_n763), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT52), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g595(.A(KEYINPUT113), .B(G86), .Z(new_n1021));
  OAI21_X1  g596(.A(new_n570), .B1(new_n593), .B2(new_n1021), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n576), .A2(G651), .ZN(new_n1023));
  OAI21_X1  g598(.A(G1981), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(G305), .B2(G1981), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT49), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g602(.A(KEYINPUT49), .B(new_n1024), .C1(G305), .C2(G1981), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n1017), .A3(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(KEYINPUT112), .B(G1976), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT52), .B1(G288), .B2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1017), .B(new_n1031), .C1(new_n763), .C2(G288), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1020), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G303), .A2(G8), .ZN(new_n1034));
  XOR2_X1   g609(.A(new_n1034), .B(KEYINPUT55), .Z(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n974), .A2(G2090), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n991), .A2(new_n992), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1971), .B1(new_n1038), .B2(new_n1002), .ZN(new_n1039));
  OAI21_X1  g614(.A(G8), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n966), .A2(new_n775), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1042), .B(KEYINPUT111), .C1(G2090), .C2(new_n974), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1035), .A2(G8), .A3(new_n1043), .A4(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1033), .A2(new_n1041), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n978), .A2(new_n980), .A3(new_n983), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n745), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n971), .A2(new_n973), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n1052));
  INV_X1    g627(.A(G2084), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1002), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT117), .B1(new_n974), .B2(G2084), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1050), .A2(G168), .A3(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1016), .A2(KEYINPUT120), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT51), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1049), .A2(new_n745), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1061), .A2(new_n1016), .A3(G168), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1057), .A2(new_n1064), .A3(new_n1058), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1060), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1011), .A2(new_n1014), .A3(new_n1048), .A4(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT124), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  XOR2_X1   g644(.A(G299), .B(KEYINPUT57), .Z(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT56), .B(G2072), .ZN(new_n1071));
  INV_X1    g646(.A(G1956), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n967), .A2(new_n1071), .B1(new_n1072), .B2(new_n974), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1348), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1015), .A2(new_n953), .B1(new_n974), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1076), .A2(new_n597), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1074), .B(KEYINPUT61), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT58), .B(G1341), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1015), .A2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n966), .A2(G1996), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n541), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n1083), .B(KEYINPUT59), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1076), .A2(new_n597), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT60), .B1(new_n1085), .B2(new_n1077), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT60), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1076), .A2(new_n1087), .A3(new_n598), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1084), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  OAI221_X1 g664(.A(new_n1078), .B1(new_n1070), .B2(new_n1073), .C1(new_n1079), .C2(new_n1089), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1057), .A2(new_n1064), .A3(new_n1058), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1064), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1047), .B1(new_n1093), .B2(new_n1063), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1094), .A2(KEYINPUT124), .A3(new_n1014), .A4(new_n1011), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1069), .A2(new_n1090), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1045), .A2(new_n1043), .A3(G8), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT118), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1045), .A2(new_n1043), .A3(new_n1099), .A4(G8), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1098), .A2(new_n1036), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n1033), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1061), .A2(new_n1016), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(G168), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1046), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1101), .A2(KEYINPUT119), .A3(new_n1033), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1104), .A2(KEYINPUT63), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT63), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1047), .B2(new_n1106), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(G305), .A2(G1981), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n765), .A2(new_n763), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(KEYINPUT114), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1114), .B1(new_n1029), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT115), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n1119), .A2(new_n1120), .A3(new_n1018), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1091), .A2(new_n1092), .A3(new_n1062), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1047), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1012), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1125), .B1(new_n1066), .B2(KEYINPUT62), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1121), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1107), .A2(new_n1033), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1113), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n964), .B1(new_n1096), .B2(new_n1129), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n942), .A2(G1996), .A3(new_n949), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(KEYINPUT46), .ZN(new_n1132));
  XOR2_X1   g707(.A(new_n1132), .B(KEYINPUT125), .Z(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(KEYINPUT46), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT126), .ZN(new_n1135));
  INV_X1    g710(.A(new_n954), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n950), .B1(new_n1136), .B2(new_n726), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1133), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(KEYINPUT47), .ZN(new_n1139));
  OAI22_X1  g714(.A1(new_n955), .A2(new_n958), .B1(G2067), .B2(new_n687), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n950), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n959), .A2(new_n950), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n963), .A2(new_n950), .ZN(new_n1143));
  XOR2_X1   g718(.A(new_n1143), .B(KEYINPUT48), .Z(new_n1144));
  OAI211_X1 g719(.A(new_n1139), .B(new_n1141), .C1(new_n1142), .C2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT127), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1130), .A2(new_n1146), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g722(.A1(new_n917), .A2(KEYINPUT43), .ZN(new_n1149));
  INV_X1    g723(.A(KEYINPUT108), .ZN(new_n1150));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g725(.A1(new_n920), .A2(new_n918), .A3(new_n926), .ZN(new_n1152));
  NAND3_X1  g726(.A1(new_n917), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n1153));
  NAND3_X1  g727(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NOR2_X1   g728(.A1(G401), .A2(G227), .ZN(new_n1155));
  AND2_X1   g729(.A1(new_n857), .A2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g730(.A1(G229), .A2(new_n462), .ZN(new_n1157));
  AND3_X1   g731(.A1(new_n1154), .A2(new_n1156), .A3(new_n1157), .ZN(G308));
  NAND3_X1  g732(.A1(new_n1154), .A2(new_n1156), .A3(new_n1157), .ZN(G225));
endmodule


