

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744;

  INV_X1 U368 ( .A(G125), .ZN(n389) );
  INV_X2 U369 ( .A(G953), .ZN(n733) );
  NAND2_X1 U370 ( .A1(n742), .A2(n740), .ZN(n559) );
  NAND2_X2 U371 ( .A1(n532), .A2(n385), .ZN(n384) );
  XNOR2_X2 U372 ( .A(n472), .B(n364), .ZN(n731) );
  XNOR2_X2 U373 ( .A(n441), .B(G134), .ZN(n472) );
  AND2_X1 U374 ( .A1(n373), .A2(n381), .ZN(n380) );
  AND2_X1 U375 ( .A1(n365), .A2(n347), .ZN(n582) );
  NAND2_X1 U376 ( .A1(n549), .A2(n660), .ZN(n665) );
  OR2_X1 U377 ( .A1(n601), .A2(G902), .ZN(n451) );
  NOR2_X2 U378 ( .A1(n665), .A2(n547), .ZN(n542) );
  NAND2_X1 U379 ( .A1(n744), .A2(n634), .ZN(n505) );
  AND2_X1 U380 ( .A1(n526), .A2(n741), .ZN(n527) );
  XNOR2_X1 U381 ( .A(n349), .B(KEYINPUT104), .ZN(n677) );
  NAND2_X1 U382 ( .A1(n351), .A2(n350), .ZN(n349) );
  INV_X1 U383 ( .A(n387), .ZN(n351) );
  INV_X1 U384 ( .A(KEYINPUT79), .ZN(n369) );
  NAND2_X1 U385 ( .A1(n514), .A2(n513), .ZN(n528) );
  AND2_X1 U386 ( .A1(n509), .A2(n508), .ZN(n514) );
  OR2_X1 U387 ( .A1(n527), .A2(KEYINPUT83), .ZN(n385) );
  NOR2_X1 U388 ( .A1(n528), .A2(KEYINPUT83), .ZN(n386) );
  XNOR2_X1 U389 ( .A(n443), .B(n442), .ZN(n364) );
  INV_X1 U390 ( .A(KEYINPUT4), .ZN(n442) );
  XNOR2_X1 U391 ( .A(n396), .B(n359), .ZN(n397) );
  NAND2_X1 U392 ( .A1(n540), .A2(n674), .ZN(n363) );
  INV_X1 U393 ( .A(KEYINPUT30), .ZN(n362) );
  XNOR2_X1 U394 ( .A(n488), .B(n487), .ZN(n616) );
  XNOR2_X1 U395 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U396 ( .A(n730), .B(n481), .ZN(n488) );
  XNOR2_X1 U397 ( .A(n502), .B(n358), .ZN(n578) );
  INV_X1 U398 ( .A(KEYINPUT87), .ZN(n358) );
  XNOR2_X1 U399 ( .A(n498), .B(n497), .ZN(n501) );
  XNOR2_X1 U400 ( .A(KEYINPUT22), .B(KEYINPUT68), .ZN(n497) );
  XNOR2_X1 U401 ( .A(n436), .B(n390), .ZN(n437) );
  BUF_X1 U402 ( .A(n499), .Z(n589) );
  XNOR2_X1 U403 ( .A(n367), .B(n366), .ZN(n365) );
  INV_X1 U404 ( .A(KEYINPUT78), .ZN(n366) );
  AND2_X1 U405 ( .A1(G224), .A2(n733), .ZN(n396) );
  XOR2_X1 U406 ( .A(KEYINPUT4), .B(KEYINPUT18), .Z(n395) );
  XOR2_X1 U407 ( .A(G119), .B(G110), .Z(n427) );
  XNOR2_X1 U408 ( .A(G113), .B(G143), .ZN(n483) );
  XNOR2_X1 U409 ( .A(n419), .B(n418), .ZN(n496) );
  INV_X1 U410 ( .A(KEYINPUT0), .ZN(n418) );
  XNOR2_X1 U411 ( .A(n460), .B(n448), .ZN(n601) );
  NAND2_X1 U412 ( .A1(n378), .A2(n377), .ZN(n376) );
  INV_X1 U413 ( .A(n386), .ZN(n377) );
  XNOR2_X1 U414 ( .A(KEYINPUT10), .B(G140), .ZN(n388) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n469) );
  XNOR2_X1 U416 ( .A(G107), .B(KEYINPUT9), .ZN(n352) );
  XNOR2_X1 U417 ( .A(n354), .B(KEYINPUT102), .ZN(n353) );
  XNOR2_X1 U418 ( .A(KEYINPUT101), .B(KEYINPUT7), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n731), .B(G146), .ZN(n460) );
  XOR2_X1 U420 ( .A(G104), .B(G101), .Z(n454) );
  XNOR2_X1 U421 ( .A(n456), .B(n399), .ZN(n400) );
  BUF_X1 U422 ( .A(n682), .Z(n692) );
  INV_X1 U423 ( .A(n548), .ZN(n360) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U426 ( .A(n489), .B(n490), .ZN(n387) );
  BUF_X1 U427 ( .A(n496), .Z(n420) );
  OR2_X2 U428 ( .A1(n501), .A2(n356), .ZN(n355) );
  NOR2_X1 U429 ( .A1(n589), .A2(n524), .ZN(n525) );
  XOR2_X1 U430 ( .A(n653), .B(KEYINPUT82), .Z(n347) );
  XNOR2_X1 U431 ( .A(n476), .B(G478), .ZN(n520) );
  INV_X1 U432 ( .A(n520), .ZN(n350) );
  XOR2_X1 U433 ( .A(n406), .B(KEYINPUT89), .Z(n348) );
  NOR2_X1 U434 ( .A1(n677), .A2(n494), .ZN(n495) );
  XNOR2_X2 U435 ( .A(n355), .B(KEYINPUT32), .ZN(n744) );
  NAND2_X1 U436 ( .A1(n357), .A2(n500), .ZN(n356) );
  INV_X1 U437 ( .A(n578), .ZN(n357) );
  XNOR2_X1 U438 ( .A(n398), .B(n397), .ZN(n401) );
  OR2_X2 U439 ( .A1(n531), .A2(KEYINPUT44), .ZN(n532) );
  XNOR2_X1 U440 ( .A(n359), .B(n388), .ZN(n730) );
  XNOR2_X2 U441 ( .A(n389), .B(G146), .ZN(n359) );
  AND2_X1 U442 ( .A1(n361), .A2(n360), .ZN(n541) );
  XNOR2_X2 U443 ( .A(n451), .B(n450), .ZN(n540) );
  NAND2_X1 U444 ( .A1(n368), .A2(n570), .ZN(n367) );
  XNOR2_X1 U445 ( .A(n743), .B(n369), .ZN(n368) );
  XNOR2_X2 U446 ( .A(n371), .B(n370), .ZN(n447) );
  XNOR2_X2 U447 ( .A(G113), .B(KEYINPUT3), .ZN(n370) );
  XNOR2_X2 U448 ( .A(G101), .B(G116), .ZN(n371) );
  XNOR2_X1 U449 ( .A(n447), .B(n482), .ZN(n372) );
  XNOR2_X1 U450 ( .A(n372), .B(n393), .ZN(n715) );
  NAND2_X1 U451 ( .A1(n374), .A2(n533), .ZN(n373) );
  NAND2_X1 U452 ( .A1(n375), .A2(n382), .ZN(n374) );
  NAND2_X1 U453 ( .A1(n383), .A2(n528), .ZN(n382) );
  INV_X1 U454 ( .A(n384), .ZN(n375) );
  NAND2_X1 U455 ( .A1(n380), .A2(n376), .ZN(n719) );
  AND2_X1 U456 ( .A1(n379), .A2(n382), .ZN(n378) );
  NOR2_X1 U457 ( .A1(n384), .A2(n533), .ZN(n379) );
  NAND2_X1 U458 ( .A1(n386), .A2(n533), .ZN(n381) );
  AND2_X1 U459 ( .A1(n527), .A2(KEYINPUT83), .ZN(n383) );
  NAND2_X1 U460 ( .A1(n350), .A2(n387), .ZN(n648) );
  NAND2_X1 U461 ( .A1(n520), .A2(n387), .ZN(n564) );
  NOR2_X1 U462 ( .A1(n350), .A2(n387), .ZN(n641) );
  AND2_X1 U463 ( .A1(n562), .A2(n561), .ZN(n645) );
  XNOR2_X2 U464 ( .A(n547), .B(n462), .ZN(n590) );
  XNOR2_X2 U465 ( .A(n461), .B(n701), .ZN(n547) );
  BUF_X1 U466 ( .A(n534), .Z(n594) );
  NAND2_X1 U467 ( .A1(n719), .A2(n732), .ZN(n598) );
  XNOR2_X2 U468 ( .A(n505), .B(KEYINPUT85), .ZN(n530) );
  XOR2_X1 U469 ( .A(n435), .B(KEYINPUT96), .Z(n390) );
  AND2_X1 U470 ( .A1(n479), .A2(G214), .ZN(n391) );
  INV_X1 U471 ( .A(n441), .ZN(n399) );
  XNOR2_X1 U472 ( .A(n480), .B(n391), .ZN(n481) );
  XNOR2_X1 U473 ( .A(n401), .B(n400), .ZN(n402) );
  INV_X1 U474 ( .A(KEYINPUT28), .ZN(n551) );
  XNOR2_X1 U475 ( .A(n551), .B(KEYINPUT108), .ZN(n552) );
  INV_X1 U476 ( .A(n590), .ZN(n502) );
  XNOR2_X1 U477 ( .A(n407), .B(n348), .ZN(n534) );
  XNOR2_X1 U478 ( .A(n493), .B(n492), .ZN(n506) );
  NOR2_X1 U479 ( .A1(n522), .A2(n549), .ZN(n504) );
  AND2_X1 U480 ( .A1(n604), .A2(G953), .ZN(n714) );
  XOR2_X1 U481 ( .A(G122), .B(G104), .Z(n482) );
  XOR2_X1 U482 ( .A(KEYINPUT69), .B(KEYINPUT16), .Z(n392) );
  XNOR2_X1 U483 ( .A(n427), .B(n392), .ZN(n393) );
  INV_X1 U484 ( .A(n715), .ZN(n403) );
  XNOR2_X1 U485 ( .A(KEYINPUT17), .B(KEYINPUT75), .ZN(n394) );
  XNOR2_X1 U486 ( .A(n395), .B(n394), .ZN(n398) );
  XOR2_X1 U487 ( .A(KEYINPUT65), .B(G107), .Z(n456) );
  XNOR2_X2 U488 ( .A(G143), .B(G128), .ZN(n441) );
  XNOR2_X1 U489 ( .A(n403), .B(n402), .ZN(n623) );
  INV_X1 U490 ( .A(KEYINPUT15), .ZN(n404) );
  XNOR2_X1 U491 ( .A(n404), .B(G902), .ZN(n599) );
  NOR2_X2 U492 ( .A1(n623), .A2(n599), .ZN(n407) );
  NOR2_X1 U493 ( .A1(G902), .A2(G237), .ZN(n405) );
  XOR2_X1 U494 ( .A(KEYINPUT72), .B(n405), .Z(n408) );
  NAND2_X1 U495 ( .A1(n408), .A2(G210), .ZN(n406) );
  NAND2_X1 U496 ( .A1(n408), .A2(G214), .ZN(n674) );
  NAND2_X1 U497 ( .A1(n534), .A2(n674), .ZN(n571) );
  XNOR2_X1 U498 ( .A(n571), .B(KEYINPUT19), .ZN(n562) );
  XOR2_X1 U499 ( .A(KEYINPUT71), .B(KEYINPUT14), .Z(n410) );
  NAND2_X1 U500 ( .A1(G237), .A2(G234), .ZN(n409) );
  XNOR2_X1 U501 ( .A(n410), .B(n409), .ZN(n413) );
  NAND2_X1 U502 ( .A1(n413), .A2(G902), .ZN(n411) );
  XNOR2_X1 U503 ( .A(n411), .B(KEYINPUT91), .ZN(n535) );
  NOR2_X1 U504 ( .A1(G898), .A2(n733), .ZN(n718) );
  NAND2_X1 U505 ( .A1(n535), .A2(n718), .ZN(n412) );
  XNOR2_X1 U506 ( .A(KEYINPUT92), .B(n412), .ZN(n416) );
  NAND2_X1 U507 ( .A1(G952), .A2(n413), .ZN(n690) );
  NOR2_X1 U508 ( .A1(G953), .A2(n690), .ZN(n414) );
  XNOR2_X1 U509 ( .A(KEYINPUT90), .B(n414), .ZN(n537) );
  INV_X1 U510 ( .A(n537), .ZN(n415) );
  NAND2_X1 U511 ( .A1(n416), .A2(n415), .ZN(n417) );
  NAND2_X1 U512 ( .A1(n562), .A2(n417), .ZN(n419) );
  XOR2_X1 U513 ( .A(KEYINPUT74), .B(KEYINPUT93), .Z(n422) );
  XNOR2_X1 U514 ( .A(G128), .B(G137), .ZN(n421) );
  XNOR2_X1 U515 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U516 ( .A(n423), .B(n730), .ZN(n431) );
  NAND2_X1 U517 ( .A1(G234), .A2(n733), .ZN(n424) );
  XOR2_X1 U518 ( .A(KEYINPUT8), .B(n424), .Z(n470) );
  NAND2_X1 U519 ( .A1(G221), .A2(n470), .ZN(n426) );
  XOR2_X1 U520 ( .A(KEYINPUT23), .B(KEYINPUT94), .Z(n425) );
  XNOR2_X1 U521 ( .A(n426), .B(n425), .ZN(n429) );
  XOR2_X1 U522 ( .A(n427), .B(KEYINPUT24), .Z(n428) );
  XNOR2_X1 U523 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U524 ( .A(n431), .B(n430), .ZN(n609) );
  NOR2_X1 U525 ( .A1(G902), .A2(n609), .ZN(n438) );
  XOR2_X1 U526 ( .A(KEYINPUT95), .B(KEYINPUT20), .Z(n434) );
  INV_X1 U527 ( .A(n599), .ZN(n432) );
  NAND2_X1 U528 ( .A1(G234), .A2(n432), .ZN(n433) );
  XNOR2_X1 U529 ( .A(n434), .B(n433), .ZN(n439) );
  NAND2_X1 U530 ( .A1(n439), .A2(G217), .ZN(n436) );
  XNOR2_X1 U531 ( .A(KEYINPUT25), .B(KEYINPUT73), .ZN(n435) );
  XNOR2_X2 U532 ( .A(n438), .B(n437), .ZN(n549) );
  NAND2_X1 U533 ( .A1(n439), .A2(G221), .ZN(n440) );
  XOR2_X1 U534 ( .A(n440), .B(KEYINPUT21), .Z(n660) );
  XNOR2_X1 U535 ( .A(G137), .B(G131), .ZN(n443) );
  NOR2_X1 U536 ( .A1(G953), .A2(G237), .ZN(n479) );
  AND2_X1 U537 ( .A1(n479), .A2(G210), .ZN(n445) );
  XNOR2_X1 U538 ( .A(KEYINPUT5), .B(G119), .ZN(n444) );
  XNOR2_X1 U539 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U540 ( .A(n447), .B(n446), .ZN(n448) );
  INV_X1 U541 ( .A(KEYINPUT67), .ZN(n449) );
  XNOR2_X1 U542 ( .A(n449), .B(G472), .ZN(n450) );
  XNOR2_X1 U543 ( .A(KEYINPUT103), .B(KEYINPUT6), .ZN(n452) );
  XNOR2_X1 U544 ( .A(n540), .B(n452), .ZN(n499) );
  INV_X1 U545 ( .A(n499), .ZN(n574) );
  NOR2_X1 U546 ( .A1(n665), .A2(n574), .ZN(n463) );
  XNOR2_X1 U547 ( .A(G110), .B(G140), .ZN(n453) );
  XNOR2_X1 U548 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U549 ( .A(n456), .B(n455), .Z(n458) );
  NAND2_X1 U550 ( .A1(G227), .A2(n733), .ZN(n457) );
  XNOR2_X1 U551 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U552 ( .A(n460), .B(n459), .ZN(n705) );
  OR2_X1 U553 ( .A1(n705), .A2(G902), .ZN(n461) );
  INV_X1 U554 ( .A(G469), .ZN(n701) );
  INV_X1 U555 ( .A(KEYINPUT1), .ZN(n462) );
  NAND2_X1 U556 ( .A1(n463), .A2(n590), .ZN(n466) );
  XNOR2_X1 U557 ( .A(KEYINPUT86), .B(KEYINPUT33), .ZN(n464) );
  XNOR2_X1 U558 ( .A(n464), .B(KEYINPUT66), .ZN(n465) );
  XNOR2_X2 U559 ( .A(n466), .B(n465), .ZN(n682) );
  NAND2_X1 U560 ( .A1(n420), .A2(n682), .ZN(n467) );
  XNOR2_X1 U561 ( .A(n467), .B(KEYINPUT34), .ZN(n491) );
  XNOR2_X1 U562 ( .A(G116), .B(G122), .ZN(n468) );
  XNOR2_X1 U563 ( .A(n469), .B(n468), .ZN(n474) );
  NAND2_X1 U564 ( .A1(G217), .A2(n470), .ZN(n471) );
  XNOR2_X1 U565 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U566 ( .A(n474), .B(n473), .ZN(n712) );
  INV_X1 U567 ( .A(G902), .ZN(n475) );
  NAND2_X1 U568 ( .A1(n712), .A2(n475), .ZN(n476) );
  XNOR2_X1 U569 ( .A(KEYINPUT13), .B(G475), .ZN(n490) );
  XOR2_X1 U570 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n478) );
  XNOR2_X1 U571 ( .A(G131), .B(KEYINPUT11), .ZN(n477) );
  XNOR2_X1 U572 ( .A(n478), .B(n477), .ZN(n480) );
  XNOR2_X1 U573 ( .A(n482), .B(KEYINPUT98), .ZN(n486) );
  XOR2_X1 U574 ( .A(KEYINPUT97), .B(KEYINPUT100), .Z(n484) );
  XNOR2_X1 U575 ( .A(n484), .B(n483), .ZN(n485) );
  NOR2_X1 U576 ( .A1(G902), .A2(n616), .ZN(n489) );
  NOR2_X2 U577 ( .A1(n491), .A2(n564), .ZN(n493) );
  XNOR2_X1 U578 ( .A(KEYINPUT80), .B(KEYINPUT35), .ZN(n492) );
  BUF_X2 U579 ( .A(n506), .Z(n529) );
  XNOR2_X1 U580 ( .A(n529), .B(G122), .ZN(G24) );
  INV_X1 U581 ( .A(n660), .ZN(n494) );
  NAND2_X1 U582 ( .A1(n496), .A2(n495), .ZN(n498) );
  NOR2_X1 U583 ( .A1(n549), .A2(n589), .ZN(n500) );
  INV_X1 U584 ( .A(n540), .ZN(n663) );
  INV_X1 U585 ( .A(n501), .ZN(n503) );
  NAND2_X1 U586 ( .A1(n503), .A2(n502), .ZN(n522) );
  NAND2_X1 U587 ( .A1(n663), .A2(n504), .ZN(n634) );
  AND2_X1 U588 ( .A1(n506), .A2(KEYINPUT84), .ZN(n507) );
  NAND2_X1 U589 ( .A1(n530), .A2(n507), .ZN(n509) );
  OR2_X1 U590 ( .A1(n510), .A2(KEYINPUT44), .ZN(n508) );
  INV_X1 U591 ( .A(KEYINPUT84), .ZN(n510) );
  NAND2_X1 U592 ( .A1(n510), .A2(KEYINPUT44), .ZN(n511) );
  NOR2_X1 U593 ( .A1(n529), .A2(n511), .ZN(n512) );
  NAND2_X1 U594 ( .A1(n530), .A2(n512), .ZN(n513) );
  INV_X1 U595 ( .A(n420), .ZN(n516) );
  NOR2_X1 U596 ( .A1(n665), .A2(n663), .ZN(n515) );
  NAND2_X1 U597 ( .A1(n515), .A2(n590), .ZN(n669) );
  NOR2_X1 U598 ( .A1(n516), .A2(n669), .ZN(n517) );
  XNOR2_X1 U599 ( .A(n517), .B(KEYINPUT31), .ZN(n650) );
  INV_X1 U600 ( .A(n542), .ZN(n518) );
  NOR2_X1 U601 ( .A1(n518), .A2(n540), .ZN(n519) );
  NAND2_X1 U602 ( .A1(n420), .A2(n519), .ZN(n637) );
  NAND2_X1 U603 ( .A1(n650), .A2(n637), .ZN(n521) );
  INV_X1 U604 ( .A(n648), .ZN(n646) );
  NOR2_X1 U605 ( .A1(n646), .A2(n641), .ZN(n679) );
  INV_X1 U606 ( .A(n679), .ZN(n563) );
  NAND2_X1 U607 ( .A1(n521), .A2(n563), .ZN(n526) );
  INV_X1 U608 ( .A(n522), .ZN(n523) );
  NAND2_X1 U609 ( .A1(n549), .A2(n523), .ZN(n524) );
  XNOR2_X1 U610 ( .A(n525), .B(KEYINPUT105), .ZN(n741) );
  NAND2_X1 U611 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U612 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n533) );
  XOR2_X1 U613 ( .A(KEYINPUT46), .B(KEYINPUT81), .Z(n560) );
  XOR2_X1 U614 ( .A(KEYINPUT38), .B(n594), .Z(n675) );
  INV_X1 U615 ( .A(n675), .ZN(n543) );
  NAND2_X1 U616 ( .A1(G953), .A2(n535), .ZN(n536) );
  NOR2_X1 U617 ( .A1(G900), .A2(n536), .ZN(n538) );
  NOR2_X1 U618 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U619 ( .A(KEYINPUT76), .B(n539), .ZN(n548) );
  NAND2_X1 U620 ( .A1(n542), .A2(n541), .ZN(n566) );
  NOR2_X1 U621 ( .A1(n543), .A2(n566), .ZN(n544) );
  XOR2_X1 U622 ( .A(n544), .B(KEYINPUT39), .Z(n586) );
  AND2_X1 U623 ( .A1(n646), .A2(n586), .ZN(n546) );
  XNOR2_X1 U624 ( .A(KEYINPUT109), .B(KEYINPUT40), .ZN(n545) );
  XNOR2_X1 U625 ( .A(n546), .B(n545), .ZN(n742) );
  XNOR2_X1 U626 ( .A(KEYINPUT110), .B(KEYINPUT42), .ZN(n558) );
  XOR2_X1 U627 ( .A(n547), .B(KEYINPUT107), .Z(n555) );
  NOR2_X1 U628 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U629 ( .A1(n550), .A2(n660), .ZN(n572) );
  NOR2_X1 U630 ( .A1(n572), .A2(n663), .ZN(n553) );
  NOR2_X1 U631 ( .A1(n555), .A2(n554), .ZN(n561) );
  NAND2_X1 U632 ( .A1(n675), .A2(n674), .ZN(n678) );
  NOR2_X1 U633 ( .A1(n677), .A2(n678), .ZN(n556) );
  XNOR2_X1 U634 ( .A(KEYINPUT41), .B(n556), .ZN(n673) );
  INV_X1 U635 ( .A(n673), .ZN(n693) );
  NAND2_X1 U636 ( .A1(n561), .A2(n693), .ZN(n557) );
  XNOR2_X1 U637 ( .A(n558), .B(n557), .ZN(n740) );
  XNOR2_X1 U638 ( .A(n560), .B(n559), .ZN(n584) );
  NAND2_X1 U639 ( .A1(n645), .A2(n563), .ZN(n579) );
  NAND2_X1 U640 ( .A1(n579), .A2(KEYINPUT47), .ZN(n570) );
  INV_X1 U641 ( .A(n564), .ZN(n568) );
  INV_X1 U642 ( .A(n594), .ZN(n565) );
  NOR2_X1 U643 ( .A1(n565), .A2(n566), .ZN(n567) );
  NAND2_X1 U644 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X2 U645 ( .A(KEYINPUT106), .B(n569), .ZN(n743) );
  INV_X1 U646 ( .A(n571), .ZN(n573) );
  NOR2_X1 U647 ( .A1(n648), .A2(n572), .ZN(n587) );
  NAND2_X1 U648 ( .A1(n573), .A2(n587), .ZN(n575) );
  NOR2_X1 U649 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U650 ( .A(KEYINPUT36), .B(n576), .Z(n577) );
  NOR2_X1 U651 ( .A1(n578), .A2(n577), .ZN(n653) );
  NOR2_X1 U652 ( .A1(n579), .A2(KEYINPUT47), .ZN(n580) );
  XOR2_X1 U653 ( .A(KEYINPUT70), .B(n580), .Z(n581) );
  NAND2_X1 U654 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U655 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U656 ( .A(KEYINPUT48), .B(n585), .Z(n597) );
  NAND2_X1 U657 ( .A1(n586), .A2(n641), .ZN(n656) );
  AND2_X1 U658 ( .A1(n674), .A2(n587), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n589), .A2(n588), .ZN(n591) );
  NOR2_X1 U660 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U661 ( .A(n592), .B(KEYINPUT43), .ZN(n593) );
  NOR2_X1 U662 ( .A1(n594), .A2(n593), .ZN(n657) );
  INV_X1 U663 ( .A(n657), .ZN(n595) );
  NAND2_X1 U664 ( .A1(n656), .A2(n595), .ZN(n596) );
  NOR2_X1 U665 ( .A1(n597), .A2(n596), .ZN(n732) );
  XNOR2_X2 U666 ( .A(n598), .B(KEYINPUT2), .ZN(n658) );
  NAND2_X2 U667 ( .A1(n658), .A2(n599), .ZN(n709) );
  INV_X1 U668 ( .A(G472), .ZN(n600) );
  NOR2_X1 U669 ( .A1(n709), .A2(n600), .ZN(n603) );
  XNOR2_X1 U670 ( .A(n601), .B(KEYINPUT62), .ZN(n602) );
  XNOR2_X1 U671 ( .A(n603), .B(n602), .ZN(n605) );
  INV_X1 U672 ( .A(G952), .ZN(n604) );
  INV_X1 U673 ( .A(n714), .ZN(n629) );
  NAND2_X1 U674 ( .A1(n605), .A2(n629), .ZN(n607) );
  XOR2_X1 U675 ( .A(KEYINPUT111), .B(KEYINPUT63), .Z(n606) );
  XNOR2_X1 U676 ( .A(n607), .B(n606), .ZN(G57) );
  INV_X1 U677 ( .A(G217), .ZN(n608) );
  NOR2_X1 U678 ( .A1(n709), .A2(n608), .ZN(n610) );
  XNOR2_X1 U679 ( .A(n610), .B(n609), .ZN(n611) );
  NAND2_X1 U680 ( .A1(n611), .A2(n629), .ZN(n612) );
  XNOR2_X1 U681 ( .A(n612), .B(KEYINPUT123), .ZN(G66) );
  INV_X1 U682 ( .A(G475), .ZN(n613) );
  NOR2_X1 U683 ( .A1(n709), .A2(n613), .ZN(n618) );
  XNOR2_X1 U684 ( .A(KEYINPUT88), .B(KEYINPUT122), .ZN(n614) );
  XOR2_X1 U685 ( .A(n614), .B(KEYINPUT59), .Z(n615) );
  XNOR2_X1 U686 ( .A(n616), .B(n615), .ZN(n617) );
  XNOR2_X1 U687 ( .A(n618), .B(n617), .ZN(n619) );
  NAND2_X1 U688 ( .A1(n619), .A2(n629), .ZN(n621) );
  INV_X1 U689 ( .A(KEYINPUT60), .ZN(n620) );
  XNOR2_X1 U690 ( .A(n621), .B(n620), .ZN(G60) );
  INV_X1 U691 ( .A(G210), .ZN(n622) );
  NOR2_X1 U692 ( .A1(n709), .A2(n622), .ZN(n628) );
  BUF_X1 U693 ( .A(n623), .Z(n626) );
  XNOR2_X1 U694 ( .A(KEYINPUT77), .B(KEYINPUT54), .ZN(n624) );
  XNOR2_X1 U695 ( .A(n624), .B(KEYINPUT55), .ZN(n625) );
  XNOR2_X1 U696 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U697 ( .A(n628), .B(n627), .ZN(n630) );
  NAND2_X1 U698 ( .A1(n630), .A2(n629), .ZN(n632) );
  XOR2_X1 U699 ( .A(KEYINPUT120), .B(KEYINPUT56), .Z(n631) );
  XNOR2_X1 U700 ( .A(n632), .B(n631), .ZN(G51) );
  XOR2_X1 U701 ( .A(G110), .B(KEYINPUT113), .Z(n633) );
  XNOR2_X1 U702 ( .A(n634), .B(n633), .ZN(G12) );
  NOR2_X1 U703 ( .A1(n648), .A2(n637), .ZN(n635) );
  XOR2_X1 U704 ( .A(KEYINPUT112), .B(n635), .Z(n636) );
  XNOR2_X1 U705 ( .A(G104), .B(n636), .ZN(G6) );
  INV_X1 U706 ( .A(n641), .ZN(n651) );
  NOR2_X1 U707 ( .A1(n651), .A2(n637), .ZN(n639) );
  XNOR2_X1 U708 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n638) );
  XNOR2_X1 U709 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U710 ( .A(G107), .B(n640), .ZN(G9) );
  XOR2_X1 U711 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n643) );
  NAND2_X1 U712 ( .A1(n645), .A2(n641), .ZN(n642) );
  XNOR2_X1 U713 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U714 ( .A(G128), .B(n644), .ZN(G30) );
  NAND2_X1 U715 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U716 ( .A(G146), .B(n647), .ZN(G48) );
  NOR2_X1 U717 ( .A1(n648), .A2(n650), .ZN(n649) );
  XOR2_X1 U718 ( .A(G113), .B(n649), .Z(G15) );
  NOR2_X1 U719 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U720 ( .A(G116), .B(n652), .Z(G18) );
  XOR2_X1 U721 ( .A(KEYINPUT37), .B(KEYINPUT115), .Z(n655) );
  XNOR2_X1 U722 ( .A(G125), .B(n653), .ZN(n654) );
  XNOR2_X1 U723 ( .A(n655), .B(n654), .ZN(G27) );
  XNOR2_X1 U724 ( .A(G134), .B(n656), .ZN(G36) );
  XOR2_X1 U725 ( .A(G140), .B(n657), .Z(G42) );
  BUF_X1 U726 ( .A(n658), .Z(n659) );
  INV_X1 U727 ( .A(n659), .ZN(n698) );
  XOR2_X1 U728 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n689) );
  NOR2_X1 U729 ( .A1(n660), .A2(n549), .ZN(n661) );
  XNOR2_X1 U730 ( .A(n661), .B(KEYINPUT49), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n662), .B(KEYINPUT116), .ZN(n664) );
  NAND2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n668) );
  AND2_X1 U733 ( .A1(n665), .A2(n502), .ZN(n666) );
  XNOR2_X1 U734 ( .A(n666), .B(KEYINPUT50), .ZN(n667) );
  OR2_X1 U735 ( .A1(n668), .A2(n667), .ZN(n670) );
  NAND2_X1 U736 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U737 ( .A(KEYINPUT51), .B(n671), .ZN(n672) );
  NOR2_X1 U738 ( .A1(n673), .A2(n672), .ZN(n686) );
  NOR2_X1 U739 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U740 ( .A1(n677), .A2(n676), .ZN(n681) );
  NOR2_X1 U741 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U742 ( .A1(n681), .A2(n680), .ZN(n684) );
  INV_X1 U743 ( .A(n692), .ZN(n683) );
  NOR2_X1 U744 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U745 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U746 ( .A(n687), .B(KEYINPUT52), .ZN(n688) );
  XNOR2_X1 U747 ( .A(n689), .B(n688), .ZN(n691) );
  NOR2_X1 U748 ( .A1(n691), .A2(n690), .ZN(n696) );
  NAND2_X1 U749 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U750 ( .A1(n694), .A2(n733), .ZN(n695) );
  NOR2_X1 U751 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U752 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U753 ( .A(n699), .B(KEYINPUT53), .ZN(n700) );
  XNOR2_X1 U754 ( .A(KEYINPUT119), .B(n700), .ZN(G75) );
  BUF_X1 U755 ( .A(n709), .Z(n702) );
  NOR2_X1 U756 ( .A1(n702), .A2(n701), .ZN(n707) );
  XOR2_X1 U757 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n703) );
  XNOR2_X1 U758 ( .A(n703), .B(KEYINPUT121), .ZN(n704) );
  XNOR2_X1 U759 ( .A(n705), .B(n704), .ZN(n706) );
  XNOR2_X1 U760 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U761 ( .A1(n714), .A2(n708), .ZN(G54) );
  INV_X1 U762 ( .A(n709), .ZN(n710) );
  NAND2_X1 U763 ( .A1(n710), .A2(G478), .ZN(n711) );
  XOR2_X1 U764 ( .A(n712), .B(n711), .Z(n713) );
  NOR2_X1 U765 ( .A1(n714), .A2(n713), .ZN(G63) );
  BUF_X1 U766 ( .A(n715), .Z(n716) );
  XNOR2_X1 U767 ( .A(n716), .B(G107), .ZN(n717) );
  NOR2_X1 U768 ( .A1(n718), .A2(n717), .ZN(n729) );
  AND2_X1 U769 ( .A1(n719), .A2(n733), .ZN(n726) );
  XOR2_X1 U770 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n721) );
  NAND2_X1 U771 ( .A1(G224), .A2(G953), .ZN(n720) );
  XNOR2_X1 U772 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U773 ( .A(KEYINPUT124), .B(n722), .ZN(n723) );
  NAND2_X1 U774 ( .A1(n723), .A2(G898), .ZN(n724) );
  XOR2_X1 U775 ( .A(KEYINPUT126), .B(n724), .Z(n725) );
  NOR2_X1 U776 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U777 ( .A(n727), .B(KEYINPUT127), .ZN(n728) );
  XNOR2_X1 U778 ( .A(n729), .B(n728), .ZN(G69) );
  XNOR2_X1 U779 ( .A(n731), .B(n730), .ZN(n735) );
  XNOR2_X1 U780 ( .A(n732), .B(n735), .ZN(n734) );
  NAND2_X1 U781 ( .A1(n734), .A2(n733), .ZN(n739) );
  XOR2_X1 U782 ( .A(G227), .B(n735), .Z(n736) );
  NAND2_X1 U783 ( .A1(n736), .A2(G900), .ZN(n737) );
  NAND2_X1 U784 ( .A1(n737), .A2(G953), .ZN(n738) );
  NAND2_X1 U785 ( .A1(n739), .A2(n738), .ZN(G72) );
  XNOR2_X1 U786 ( .A(G137), .B(n740), .ZN(G39) );
  XNOR2_X1 U787 ( .A(G101), .B(n741), .ZN(G3) );
  XNOR2_X1 U788 ( .A(G131), .B(n742), .ZN(G33) );
  XNOR2_X1 U789 ( .A(G143), .B(n743), .ZN(G45) );
  XNOR2_X1 U790 ( .A(n744), .B(G119), .ZN(G21) );
endmodule

