//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:34:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1285, new_n1286, new_n1287, new_n1289, new_n1290, new_n1291,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  OAI21_X1  g0003(.A(KEYINPUT64), .B1(new_n203), .B2(G50), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  NOR2_X1   g0005(.A1(G58), .A2(G68), .ZN(new_n206));
  INV_X1    g0006(.A(KEYINPUT64), .ZN(new_n207));
  INV_X1    g0007(.A(G50), .ZN(new_n208));
  NAND3_X1  g0008(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  AND3_X1   g0009(.A1(new_n204), .A2(new_n205), .A3(new_n209), .ZN(G353));
  OAI21_X1  g0010(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n216));
  AND3_X1   g0016(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n217));
  AOI21_X1  g0017(.A(KEYINPUT65), .B1(G1), .B2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n203), .A2(G50), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n216), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT66), .Z(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  INV_X1    g0028(.A(G238), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n228), .B1(new_n202), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT67), .B(G77), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n230), .B1(G244), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(KEYINPUT68), .ZN(new_n233));
  AOI22_X1  g0033(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n234));
  AOI22_X1  g0034(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n232), .A2(KEYINPUT68), .ZN(new_n237));
  OAI21_X1  g0037(.A(new_n212), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g0038(.A(new_n227), .B1(KEYINPUT1), .B2(new_n238), .ZN(new_n239));
  AOI21_X1  g0039(.A(new_n239), .B1(KEYINPUT1), .B2(new_n238), .ZN(G361));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  INV_X1    g0041(.A(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(KEYINPUT2), .B(G226), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G264), .B(G270), .Z(new_n246));
  XNOR2_X1  g0046(.A(G250), .B(G257), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G358));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n208), .A2(G68), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n202), .A2(G50), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(G58), .B(G77), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n252), .B(new_n257), .ZN(G351));
  INV_X1    g0058(.A(KEYINPUT81), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT8), .B(G58), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n260), .B1(new_n261), .B2(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G1), .A2(G13), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT65), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n266));
  NAND3_X1  g0066(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  AND4_X1   g0068(.A1(new_n265), .A2(new_n266), .A3(new_n267), .A4(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n266), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n262), .A2(new_n269), .B1(new_n270), .B2(new_n260), .ZN(new_n271));
  OR2_X1    g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n272), .A2(KEYINPUT7), .A3(new_n220), .A4(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT75), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n279), .A2(KEYINPUT75), .A3(KEYINPUT7), .A4(new_n220), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n272), .A2(new_n220), .A3(new_n273), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT7), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n276), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G68), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT76), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G58), .A2(G68), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n286), .B(G20), .C1(new_n288), .C2(new_n206), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G159), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n203), .A2(new_n287), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n286), .B1(new_n293), .B2(G20), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT16), .ZN(new_n295));
  NOR3_X1   g0095(.A1(new_n292), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n285), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n283), .A2(KEYINPUT77), .A3(new_n274), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT77), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n279), .A2(new_n301), .A3(KEYINPUT7), .A4(new_n220), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n300), .A2(G68), .A3(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n292), .A2(new_n294), .ZN(new_n304));
  AOI21_X1  g0104(.A(KEYINPUT16), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n271), .B1(new_n299), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT78), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT78), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n308), .B(new_n271), .C1(new_n299), .C2(new_n305), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G41), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(new_n217), .B2(new_n218), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G87), .ZN(new_n312));
  OR2_X1    g0112(.A1(G223), .A2(G1698), .ZN(new_n313));
  INV_X1    g0113(.A(G226), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G1698), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n313), .B(new_n315), .C1(new_n277), .C2(new_n278), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n311), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G274), .ZN(new_n318));
  AND2_X1   g0118(.A1(G1), .A2(G13), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n318), .B1(new_n319), .B2(new_n310), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n319), .A2(new_n310), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(G232), .A3(new_n321), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n317), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G169), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(G179), .B2(new_n327), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n307), .A2(new_n309), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT18), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT18), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n307), .A2(new_n309), .A3(new_n334), .A4(new_n331), .ZN(new_n335));
  INV_X1    g0135(.A(new_n271), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n303), .A2(new_n304), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n295), .ZN(new_n338));
  INV_X1    g0138(.A(new_n298), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n339), .B1(new_n285), .B2(new_n296), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n336), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G200), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n317), .B2(new_n326), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n316), .A2(new_n312), .ZN(new_n344));
  INV_X1    g0144(.A(new_n311), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G190), .ZN(new_n347));
  INV_X1    g0147(.A(G41), .ZN(new_n348));
  INV_X1    g0148(.A(G45), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n261), .A2(new_n350), .B1(new_n319), .B2(new_n310), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n351), .A2(G232), .B1(new_n320), .B2(new_n322), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n346), .A2(new_n347), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n343), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT79), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n343), .A2(new_n353), .A3(KEYINPUT79), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AND3_X1   g0158(.A1(new_n341), .A2(KEYINPUT17), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT17), .B1(new_n341), .B2(new_n358), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n333), .A2(new_n335), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT80), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT80), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n333), .A2(new_n361), .A3(new_n364), .A4(new_n335), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n220), .A2(G33), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT71), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n220), .A2(KEYINPUT71), .A3(G33), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(G77), .A3(new_n369), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n290), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT74), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(new_n373), .A3(new_n298), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n373), .B1(new_n372), .B2(new_n298), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT11), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n372), .A2(new_n298), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT74), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT11), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(new_n380), .A3(new_n374), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n270), .A2(new_n202), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n382), .B(KEYINPUT12), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n261), .A2(G20), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n269), .A2(G68), .A3(new_n384), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n377), .A2(new_n381), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n242), .A2(G1698), .ZN(new_n388));
  OAI221_X1 g0188(.A(new_n388), .B1(G226), .B2(G1698), .C1(new_n277), .C2(new_n278), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G97), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n311), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT13), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n351), .A2(G238), .B1(new_n320), .B2(new_n322), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n324), .A2(new_n321), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n323), .B1(new_n229), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT13), .B1(new_n391), .B2(new_n397), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n395), .A2(new_n398), .A3(G190), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n342), .B1(new_n395), .B2(new_n398), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n387), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n395), .A2(new_n398), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G169), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT14), .ZN(new_n404));
  INV_X1    g0204(.A(new_n402), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G179), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT14), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n402), .A2(new_n407), .A3(G169), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n404), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n401), .B1(new_n409), .B2(new_n387), .ZN(new_n410));
  AOI21_X1  g0210(.A(G1698), .B1(new_n272), .B2(new_n273), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G222), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n272), .A2(new_n273), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(G223), .A3(G1698), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n279), .A2(new_n231), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n345), .ZN(new_n417));
  OR2_X1    g0217(.A1(new_n314), .A2(KEYINPUT69), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n314), .A2(KEYINPUT69), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n324), .A2(new_n418), .A3(new_n321), .A4(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n323), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT70), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT70), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n420), .A2(new_n323), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n417), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n328), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n368), .A2(new_n369), .ZN(new_n427));
  INV_X1    g0227(.A(G150), .ZN(new_n428));
  INV_X1    g0228(.A(new_n290), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n427), .A2(new_n260), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n220), .B1(new_n204), .B2(new_n209), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n298), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n208), .B1(new_n261), .B2(G20), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n269), .A2(new_n433), .B1(new_n208), .B2(new_n270), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n426), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n425), .A2(G179), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n425), .A2(G200), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT9), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n417), .A2(G190), .A3(new_n422), .A4(new_n424), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n432), .A2(KEYINPUT9), .A3(new_n434), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT10), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n443), .A2(new_n444), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT10), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(new_n439), .A4(new_n441), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n438), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n231), .A2(G20), .ZN(new_n451));
  XNOR2_X1  g0251(.A(KEYINPUT15), .B(G87), .ZN(new_n452));
  OAI221_X1 g0252(.A(new_n451), .B1(new_n429), .B2(new_n260), .C1(new_n366), .C2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n298), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n269), .A2(G77), .A3(new_n384), .ZN(new_n455));
  INV_X1    g0255(.A(new_n231), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n270), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT73), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n454), .A2(KEYINPUT73), .A3(new_n455), .A4(new_n457), .ZN(new_n461));
  INV_X1    g0261(.A(G1698), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n413), .A2(G232), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n413), .A2(G238), .A3(G1698), .ZN(new_n464));
  INV_X1    g0264(.A(G107), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n463), .B(new_n464), .C1(new_n465), .C2(new_n413), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n345), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n351), .A2(G244), .B1(new_n320), .B2(new_n322), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G200), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n460), .A2(new_n461), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n469), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(KEYINPUT72), .A3(G190), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT72), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n469), .B2(new_n347), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n460), .A2(new_n461), .ZN(new_n477));
  AOI21_X1  g0277(.A(G169), .B1(new_n467), .B2(new_n468), .ZN(new_n478));
  INV_X1    g0278(.A(G179), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n478), .B1(new_n472), .B2(new_n479), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n471), .A2(new_n476), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n410), .A2(new_n450), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  AND4_X1   g0283(.A1(new_n259), .A2(new_n363), .A3(new_n365), .A4(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n482), .B1(new_n362), .B2(KEYINPUT80), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n259), .B1(new_n485), .B2(new_n365), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n300), .A2(G107), .A3(new_n302), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT6), .ZN(new_n489));
  INV_X1    g0289(.A(G97), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(new_n465), .ZN(new_n491));
  NOR2_X1   g0291(.A1(G97), .A2(G107), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n465), .A2(KEYINPUT82), .A3(KEYINPUT6), .A4(G97), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT82), .ZN(new_n495));
  NAND2_X1  g0295(.A1(KEYINPUT6), .A2(G97), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(G107), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n493), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n498), .A2(G20), .B1(G77), .B2(new_n290), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n339), .B1(new_n488), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n266), .A2(G97), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT83), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n261), .B2(G33), .ZN(new_n504));
  INV_X1    g0304(.A(G33), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n505), .A2(KEYINPUT83), .A3(G1), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n269), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n502), .B1(new_n508), .B2(new_n490), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n500), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n349), .A2(G1), .ZN(new_n511));
  AND2_X1   g0311(.A1(KEYINPUT5), .A2(G41), .ZN(new_n512));
  NOR2_X1   g0312(.A1(KEYINPUT5), .A2(G41), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n514), .A2(G257), .A3(new_n324), .ZN(new_n515));
  OAI211_X1 g0315(.A(G244), .B(new_n462), .C1(new_n277), .C2(new_n278), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT4), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n413), .A2(KEYINPUT4), .A3(G244), .A4(new_n462), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G283), .ZN(new_n520));
  OAI211_X1 g0320(.A(G250), .B(G1698), .C1(new_n277), .C2(new_n278), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n518), .A2(new_n519), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n515), .B1(new_n522), .B2(new_n345), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT84), .ZN(new_n524));
  XNOR2_X1  g0324(.A(KEYINPUT5), .B(G41), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n320), .A2(new_n511), .A3(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n523), .A2(new_n524), .A3(G190), .A4(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n520), .B(new_n521), .C1(new_n516), .C2(new_n517), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT4), .B1(new_n411), .B2(G244), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n345), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n515), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n526), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT84), .B1(new_n532), .B2(G200), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n532), .A2(new_n347), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n510), .B(new_n527), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n532), .A2(new_n328), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n523), .A2(new_n479), .A3(new_n526), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n536), .B(new_n537), .C1(new_n500), .C2(new_n509), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n525), .A2(new_n511), .B1(new_n319), .B2(new_n310), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n261), .A2(G45), .ZN(new_n541));
  INV_X1    g0341(.A(new_n513), .ZN(new_n542));
  NAND2_X1  g0342(.A1(KEYINPUT5), .A2(G41), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n540), .A2(G264), .B1(new_n320), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(G257), .B(G1698), .C1(new_n277), .C2(new_n278), .ZN(new_n546));
  OAI211_X1 g0346(.A(G250), .B(new_n462), .C1(new_n277), .C2(new_n278), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G294), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n345), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n545), .A2(new_n347), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(G200), .B1(new_n545), .B2(new_n550), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n508), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT25), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n266), .B2(G107), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n270), .A2(KEYINPUT25), .A3(new_n465), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n555), .A2(G107), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT89), .ZN(new_n560));
  OAI21_X1  g0360(.A(KEYINPUT23), .B1(new_n220), .B2(G107), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT23), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n562), .A2(new_n465), .A3(G20), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n220), .A2(G33), .A3(G116), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT88), .ZN(new_n566));
  OR2_X1    g0366(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n567));
  NAND2_X1  g0367(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT22), .ZN(new_n571));
  AOI21_X1  g0371(.A(G20), .B1(new_n272), .B2(new_n273), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n571), .B1(new_n572), .B2(G87), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n220), .B(G87), .C1(new_n277), .C2(new_n278), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n574), .A2(KEYINPUT22), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n570), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n567), .A2(new_n566), .A3(new_n568), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n574), .A2(KEYINPUT22), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n413), .A2(new_n571), .A3(new_n220), .A4(G87), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n577), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n582), .A3(new_n570), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n560), .B1(new_n584), .B2(new_n298), .ZN(new_n585));
  AOI211_X1 g0385(.A(KEYINPUT89), .B(new_n339), .C1(new_n578), .C2(new_n583), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n554), .B(new_n559), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n559), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n581), .A2(new_n582), .A3(new_n570), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n582), .B1(new_n581), .B2(new_n570), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n298), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT89), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n584), .A2(new_n560), .A3(new_n298), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n588), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n545), .A2(new_n550), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n328), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(G179), .B2(new_n595), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n587), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n269), .A2(G116), .A3(new_n507), .ZN(new_n599));
  INV_X1    g0399(.A(G116), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n270), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(G20), .B1(G33), .B2(G283), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n505), .A2(G97), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n602), .A2(new_n603), .B1(G20), .B2(new_n600), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n604), .A2(new_n298), .A3(KEYINPUT20), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT20), .B1(new_n604), .B2(new_n298), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n599), .B(new_n601), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n540), .A2(G270), .B1(new_n320), .B2(new_n544), .ZN(new_n608));
  OAI211_X1 g0408(.A(G264), .B(G1698), .C1(new_n277), .C2(new_n278), .ZN(new_n609));
  OAI211_X1 g0409(.A(G257), .B(new_n462), .C1(new_n277), .C2(new_n278), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n272), .A2(G303), .A3(new_n273), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n345), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n607), .A2(new_n614), .A3(KEYINPUT21), .A4(G169), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n514), .A2(G270), .A3(new_n324), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n526), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n345), .B2(new_n612), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n618), .A2(new_n607), .A3(G179), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n328), .B1(new_n608), .B2(new_n613), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT21), .B1(new_n621), .B2(new_n607), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n614), .A2(G200), .ZN(new_n624));
  INV_X1    g0424(.A(new_n607), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n624), .B(new_n625), .C1(new_n347), .C2(new_n614), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT85), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(new_n508), .B2(new_n452), .ZN(new_n628));
  INV_X1    g0428(.A(new_n452), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n269), .A2(KEYINPUT85), .A3(new_n629), .A4(new_n507), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT19), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n220), .B1(new_n390), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(G87), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n492), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n220), .B(G68), .C1(new_n277), .C2(new_n278), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n631), .B1(new_n366), .B2(new_n490), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n638), .A2(new_n298), .B1(new_n270), .B2(new_n452), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n628), .A2(new_n630), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(G33), .A2(G116), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n229), .A2(new_n462), .ZN(new_n642));
  INV_X1    g0442(.A(G244), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(G1698), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n642), .B(new_n644), .C1(new_n277), .C2(new_n278), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n311), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n320), .A2(new_n511), .ZN(new_n647));
  INV_X1    g0447(.A(G250), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n648), .B1(new_n261), .B2(G45), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n324), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(G169), .B1(new_n646), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n645), .A2(new_n641), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n345), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n320), .A2(new_n511), .B1(new_n324), .B2(new_n649), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G179), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n640), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(G238), .A2(G1698), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(new_n643), .B2(G1698), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n660), .A2(new_n413), .B1(G33), .B2(G116), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n655), .B1(new_n661), .B2(new_n311), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G200), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n555), .A2(G87), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n654), .A2(G190), .A3(new_n655), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n663), .A2(new_n639), .A3(new_n664), .A4(new_n665), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n658), .A2(KEYINPUT86), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(KEYINPUT86), .B1(new_n658), .B2(new_n666), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n623), .B(new_n626), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  NOR4_X1   g0469(.A1(new_n487), .A2(new_n539), .A3(new_n598), .A4(new_n669), .ZN(G372));
  INV_X1    g0470(.A(new_n487), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n658), .B(KEYINPUT90), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n658), .A2(new_n666), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n587), .A2(new_n538), .A3(new_n535), .A4(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n622), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n676), .A2(new_n619), .A3(new_n615), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n559), .B1(new_n585), .B2(new_n586), .ZN(new_n678));
  INV_X1    g0478(.A(new_n597), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n672), .B1(new_n675), .B2(new_n680), .ZN(new_n681));
  OAI22_X1  g0481(.A1(new_n500), .A2(new_n509), .B1(new_n532), .B2(G179), .ZN(new_n682));
  INV_X1    g0482(.A(new_n536), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT91), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n509), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n488), .A2(new_n499), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n685), .B1(new_n686), .B2(new_n339), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT91), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n687), .A2(new_n688), .A3(new_n536), .A4(new_n537), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT26), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n684), .A2(new_n689), .A3(new_n690), .A4(new_n674), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT86), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n673), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n658), .A2(KEYINPUT86), .A3(new_n666), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n538), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n691), .B1(new_n695), .B2(new_n690), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n681), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n671), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n477), .A2(new_n480), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n401), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(new_n387), .B2(new_n409), .ZN(new_n701));
  INV_X1    g0501(.A(new_n361), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n331), .A2(new_n306), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT18), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n446), .A2(new_n449), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n438), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n698), .A2(new_n709), .ZN(G369));
  NAND3_X1  g0510(.A1(new_n261), .A2(new_n220), .A3(G13), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT27), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT27), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n713), .A2(new_n261), .A3(new_n220), .A4(G13), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n712), .A2(G213), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT92), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n712), .A2(KEYINPUT92), .A3(G213), .A4(new_n714), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(G343), .ZN(new_n720));
  OAI21_X1  g0520(.A(KEYINPUT93), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT93), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n717), .A2(new_n722), .A3(G343), .A4(new_n718), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n625), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n677), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n676), .A2(new_n626), .A3(new_n619), .A4(new_n615), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n727), .B1(new_n728), .B2(new_n726), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G330), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n592), .A2(new_n593), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n597), .B1(new_n732), .B2(new_n559), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n724), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n594), .A2(new_n725), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n734), .B1(new_n598), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT94), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n724), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n733), .A2(new_n739), .ZN(new_n740));
  AOI211_X1 g0540(.A(new_n588), .B(new_n553), .C1(new_n592), .C2(new_n593), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n733), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n677), .A2(new_n725), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n737), .A2(new_n740), .A3(new_n745), .ZN(G399));
  INV_X1    g0546(.A(KEYINPUT95), .ZN(new_n747));
  INV_X1    g0547(.A(new_n213), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n747), .B1(new_n748), .B2(G41), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n213), .A2(KEYINPUT95), .A3(new_n348), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n634), .A2(G116), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n751), .A2(G1), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(new_n222), .B2(new_n751), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT28), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT29), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n684), .A2(new_n689), .A3(KEYINPUT26), .A4(new_n674), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT96), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n757), .B(new_n758), .C1(KEYINPUT26), .C2(new_n695), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n623), .B1(new_n594), .B2(new_n597), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n673), .B1(new_n594), .B2(new_n554), .ZN(new_n761));
  AND2_X1   g0561(.A1(new_n535), .A2(new_n538), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n673), .B1(new_n538), .B2(KEYINPUT91), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n764), .A2(KEYINPUT96), .A3(KEYINPUT26), .A4(new_n689), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n759), .A2(new_n672), .A3(new_n763), .A4(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n756), .B1(new_n766), .B2(new_n725), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n756), .B(new_n739), .C1(new_n681), .C2(new_n696), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G330), .ZN(new_n770));
  INV_X1    g0570(.A(new_n669), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n742), .A2(new_n762), .A3(new_n771), .A4(new_n739), .ZN(new_n772));
  AND3_X1   g0572(.A1(new_n608), .A2(G179), .A3(new_n613), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n545), .A2(new_n550), .ZN(new_n774));
  INV_X1    g0574(.A(new_n662), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n773), .A2(new_n774), .A3(new_n523), .A4(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(KEYINPUT30), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT30), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n545), .A2(new_n550), .A3(new_n654), .A4(new_n655), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n608), .A2(new_n613), .A3(G179), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n778), .B1(new_n781), .B2(new_n523), .ZN(new_n782));
  AND3_X1   g0582(.A1(new_n530), .A2(new_n526), .A3(new_n531), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n595), .A2(new_n614), .A3(new_n479), .A4(new_n662), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n777), .A2(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(KEYINPUT31), .B1(new_n785), .B2(new_n724), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n784), .A2(new_n783), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n776), .A2(KEYINPUT30), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n781), .A2(new_n778), .A3(new_n523), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT31), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n790), .A2(new_n739), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n786), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n770), .B1(new_n772), .B2(new_n793), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n767), .A2(new_n769), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n755), .B1(new_n795), .B2(G1), .ZN(G364));
  INV_X1    g0596(.A(new_n751), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n220), .A2(G13), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n261), .B1(new_n798), .B2(G45), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n731), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(G330), .B2(new_n729), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n801), .B(KEYINPUT97), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n219), .B1(G20), .B2(new_n328), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n806), .A2(KEYINPUT99), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(KEYINPUT99), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G13), .A2(G33), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(G20), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n279), .A2(new_n213), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(new_n349), .B2(new_n223), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n257), .B2(new_n349), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n748), .A2(new_n279), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n817), .A2(G355), .B1(new_n600), .B2(new_n748), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT98), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n813), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(new_n820), .B2(new_n819), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n220), .A2(G179), .ZN(new_n823));
  NOR2_X1   g0623(.A1(G190), .A2(G200), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(G159), .ZN(new_n826));
  OAI21_X1  g0626(.A(KEYINPUT32), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(G20), .A2(G179), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(G200), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(new_n347), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n830), .A2(G190), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n827), .B1(new_n832), .B2(new_n208), .C1(new_n202), .C2(new_n834), .ZN(new_n835));
  NOR3_X1   g0635(.A1(new_n347), .A2(G179), .A3(G200), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n836), .A2(new_n220), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n823), .A2(G190), .A3(G200), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n838), .A2(G97), .B1(new_n840), .B2(G87), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n823), .A2(new_n347), .A3(G200), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(G107), .ZN(new_n844));
  INV_X1    g0644(.A(new_n825), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(G159), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n841), .B(new_n844), .C1(KEYINPUT32), .C2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n829), .A2(new_n824), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n828), .A2(new_n347), .A3(G200), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n413), .B1(new_n456), .B2(new_n848), .C1(new_n201), .C2(new_n850), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n835), .A2(new_n847), .A3(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(G317), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT33), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n853), .A2(KEYINPUT33), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n833), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n831), .A2(G326), .ZN(new_n857));
  INV_X1    g0657(.A(G294), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n856), .B(new_n857), .C1(new_n858), .C2(new_n837), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n845), .A2(G329), .B1(new_n849), .B2(G322), .ZN(new_n860));
  INV_X1    g0660(.A(G311), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n860), .B(new_n279), .C1(new_n861), .C2(new_n848), .ZN(new_n862));
  INV_X1    g0662(.A(G283), .ZN(new_n863));
  INV_X1    g0663(.A(G303), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n863), .A2(new_n842), .B1(new_n839), .B2(new_n864), .ZN(new_n865));
  NOR3_X1   g0665(.A1(new_n859), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n852), .A2(new_n866), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n805), .B(new_n822), .C1(new_n809), .C2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n812), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n868), .B1(new_n729), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n803), .A2(new_n870), .ZN(G396));
  NAND2_X1  g0671(.A1(new_n697), .A2(new_n739), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT100), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n699), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n471), .A2(new_n476), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n477), .A2(new_n724), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n477), .A2(new_n480), .A3(KEYINPUT100), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n874), .A2(new_n875), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n699), .B2(new_n725), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n872), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n879), .B(new_n739), .C1(new_n681), .C2(new_n696), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n794), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT101), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n801), .B1(new_n883), .B2(new_n884), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n809), .ZN(new_n889));
  INV_X1    g0689(.A(new_n848), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n890), .A2(G159), .B1(G143), .B2(new_n849), .ZN(new_n891));
  INV_X1    g0691(.A(G137), .ZN(new_n892));
  OAI221_X1 g0692(.A(new_n891), .B1(new_n832), .B2(new_n892), .C1(new_n428), .C2(new_n834), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT34), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n842), .A2(new_n202), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n279), .B(new_n897), .C1(G132), .C2(new_n845), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n838), .A2(G58), .B1(new_n840), .B2(G50), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n895), .A2(new_n896), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n832), .A2(new_n864), .B1(new_n839), .B2(new_n465), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(G87), .B2(new_n843), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n413), .B1(G294), .B2(new_n849), .ZN(new_n903));
  AOI22_X1  g0703(.A1(G311), .A2(new_n845), .B1(new_n890), .B2(G116), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n838), .A2(G97), .B1(new_n833), .B2(G283), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n902), .A2(new_n903), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n889), .B1(new_n900), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n809), .A2(new_n810), .ZN(new_n908));
  AOI211_X1 g0708(.A(new_n805), .B(new_n907), .C1(new_n205), .C2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n879), .B2(new_n811), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n888), .A2(new_n910), .ZN(G384));
  OR2_X1    g0711(.A1(new_n498), .A2(KEYINPUT35), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n498), .A2(KEYINPUT35), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n912), .A2(G116), .A3(new_n221), .A4(new_n913), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT36), .Z(new_n915));
  NAND3_X1  g0715(.A1(new_n223), .A2(new_n231), .A3(new_n287), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n261), .B(G13), .C1(new_n916), .C2(new_n253), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n874), .A2(new_n877), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n725), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n882), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n387), .A2(new_n724), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n410), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n409), .A2(new_n387), .A3(new_n724), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n921), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n285), .A2(new_n304), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n295), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n336), .B1(new_n929), .B2(new_n340), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n930), .A2(new_n719), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n362), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n719), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n307), .A2(new_n309), .A3(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT37), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n341), .A2(new_n358), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n332), .A2(new_n934), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n936), .B1(new_n330), .B2(new_n930), .ZN(new_n938));
  OAI21_X1  g0738(.A(KEYINPUT37), .B1(new_n938), .B2(new_n931), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT38), .B1(new_n932), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n932), .A2(KEYINPUT38), .A3(new_n940), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n927), .A2(new_n944), .B1(new_n705), .B2(new_n719), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT39), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n307), .A2(new_n309), .A3(new_n933), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n704), .A2(new_n936), .ZN(new_n948));
  OAI21_X1  g0748(.A(KEYINPUT37), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT102), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n704), .A2(new_n936), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n935), .B1(new_n952), .B2(new_n934), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(KEYINPUT102), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n951), .A2(new_n954), .A3(new_n937), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n947), .B1(new_n702), .B2(new_n705), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT38), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n943), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n946), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n409), .A2(new_n387), .A3(new_n725), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n942), .A2(KEYINPUT39), .A3(new_n943), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT103), .ZN(new_n964));
  AND3_X1   g0764(.A1(new_n945), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n964), .B1(new_n945), .B2(new_n963), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n484), .A2(new_n486), .B1(new_n767), .B2(new_n769), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n709), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n967), .B(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT105), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n957), .B2(new_n958), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n937), .B1(new_n953), .B2(KEYINPUT102), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n949), .A2(new_n950), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n956), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT38), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n977), .A2(KEYINPUT105), .A3(new_n943), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT104), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n724), .B(KEYINPUT94), .ZN(new_n980));
  NOR4_X1   g0780(.A1(new_n598), .A2(new_n669), .A3(new_n539), .A4(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n785), .A2(KEYINPUT31), .A3(new_n724), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n791), .B1(new_n790), .B2(new_n725), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n979), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n982), .A2(new_n983), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n772), .A2(new_n986), .A3(KEYINPUT104), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n923), .A2(new_n924), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n880), .A2(new_n989), .ZN(new_n990));
  AND3_X1   g0790(.A1(new_n988), .A2(KEYINPUT40), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n972), .A2(new_n978), .A3(new_n991), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n988), .B(new_n990), .C1(new_n958), .C2(new_n941), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT40), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n671), .A2(new_n988), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n997), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n998), .A2(G330), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n970), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n261), .B2(new_n798), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n970), .A2(new_n1000), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n918), .B1(new_n1002), .B2(new_n1003), .ZN(G367));
  NAND2_X1  g0804(.A1(new_n664), .A2(new_n639), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n724), .A2(new_n1005), .ZN(new_n1006));
  MUX2_X1   g0806(.A(new_n672), .B(new_n673), .S(new_n1006), .Z(new_n1007));
  INV_X1    g0807(.A(KEYINPUT43), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n538), .B(new_n535), .C1(new_n739), .C2(new_n510), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n739), .A2(new_n538), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT106), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n733), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n538), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n739), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1012), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1018), .A2(new_n745), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT42), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1009), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1017), .A2(new_n1008), .A3(new_n1007), .A4(new_n1020), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1014), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1026), .A2(new_n737), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1025), .B(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n751), .B(KEYINPUT41), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n745), .B1(new_n736), .B2(new_n744), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n731), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n730), .B(new_n745), .C1(new_n736), .C2(new_n744), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n766), .A2(new_n725), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(KEYINPUT29), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1033), .A2(new_n1035), .A3(new_n768), .A4(new_n884), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(KEYINPUT107), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT107), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n795), .A2(new_n1038), .A3(new_n1033), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(KEYINPUT108), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT108), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1037), .A2(new_n1039), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n745), .A2(new_n740), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n1018), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT44), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n745), .A2(new_n1012), .A3(new_n740), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT45), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1047), .A2(new_n737), .A3(new_n1050), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n731), .B(new_n736), .C1(new_n1046), .C2(new_n1049), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1041), .A2(new_n1043), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1029), .B1(new_n1053), .B2(new_n795), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1028), .B1(new_n1054), .B2(new_n800), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n837), .A2(new_n202), .B1(new_n456), .B2(new_n842), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n831), .A2(G143), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1057), .B(new_n413), .C1(new_n428), .C2(new_n850), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n833), .A2(G159), .B1(new_n890), .B2(G50), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1056), .B(new_n1058), .C1(KEYINPUT110), .C2(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n839), .A2(new_n201), .B1(new_n825), .B2(new_n892), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT111), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1060), .B(new_n1062), .C1(KEYINPUT110), .C2(new_n1059), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT112), .Z(new_n1064));
  OAI21_X1  g0864(.A(new_n279), .B1(new_n848), .B2(new_n863), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n850), .A2(new_n864), .B1(new_n825), .B2(new_n853), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n839), .A2(new_n600), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1065), .B(new_n1066), .C1(KEYINPUT46), .C2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(KEYINPUT46), .B2(new_n1067), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n834), .A2(new_n858), .B1(new_n842), .B2(new_n490), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n832), .A2(new_n861), .B1(new_n465), .B2(new_n837), .ZN(new_n1071));
  NOR3_X1   g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1064), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n889), .B1(new_n1073), .B2(KEYINPUT47), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(KEYINPUT47), .B2(new_n1073), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1007), .A2(new_n812), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n813), .B1(new_n213), .B2(new_n452), .C1(new_n248), .C2(new_n814), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1077), .A2(KEYINPUT109), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1077), .A2(KEYINPUT109), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n1078), .A2(new_n1079), .A3(new_n805), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1075), .A2(new_n1076), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1055), .A2(new_n1081), .ZN(G387));
  OAI211_X1 g0882(.A(new_n1040), .B(new_n797), .C1(new_n795), .C2(new_n1033), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n817), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n1084), .A2(new_n752), .B1(G107), .B2(new_n213), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n245), .A2(new_n349), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n752), .B(new_n349), .C1(new_n202), .C2(new_n205), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n1088));
  NOR3_X1   g0888(.A1(new_n1088), .A2(G50), .A3(new_n260), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1088), .B1(G50), .B2(new_n260), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n814), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1085), .B1(new_n1086), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n813), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n804), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n825), .A2(new_n428), .B1(new_n848), .B2(new_n202), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n279), .B(new_n1096), .C1(G50), .C2(new_n849), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n840), .A2(new_n231), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n837), .A2(new_n452), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n260), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1099), .B1(new_n1100), .B2(new_n833), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G159), .A2(new_n831), .B1(new_n843), .B2(G97), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1097), .A2(new_n1098), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n413), .B1(new_n845), .B2(G326), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n837), .A2(new_n863), .B1(new_n839), .B2(new_n858), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n890), .A2(G303), .B1(G317), .B2(new_n849), .ZN(new_n1106));
  INV_X1    g0906(.A(G322), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1106), .B1(new_n832), .B2(new_n1107), .C1(new_n861), .C2(new_n834), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT48), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1105), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n1109), .B2(new_n1108), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT49), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n1104), .B1(new_n600), .B2(new_n842), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1103), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1095), .B1(new_n1115), .B2(new_n809), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n736), .B2(new_n869), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT114), .Z(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n800), .B2(new_n1033), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1083), .A2(new_n1119), .ZN(G393));
  NOR2_X1   g0920(.A1(new_n252), .A2(new_n814), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(G97), .B2(new_n748), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n805), .B1(new_n813), .B2(new_n1122), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n837), .A2(new_n205), .B1(new_n848), .B2(new_n260), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n831), .A2(G150), .B1(G159), .B2(new_n849), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT51), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1124), .B(new_n1126), .C1(G50), .C2(new_n833), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n279), .B1(new_n845), .B2(G143), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1128), .B1(new_n202), .B2(new_n839), .C1(new_n633), .C2(new_n842), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT115), .Z(new_n1130));
  AOI22_X1  g0930(.A1(new_n831), .A2(G317), .B1(G311), .B2(new_n849), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT52), .Z(new_n1132));
  OAI21_X1  g0932(.A(new_n844), .B1(new_n834), .B2(new_n864), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n279), .B1(new_n848), .B2(new_n858), .C1(new_n1107), .C2(new_n825), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n837), .A2(new_n600), .B1(new_n839), .B2(new_n863), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1127), .A2(new_n1130), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1123), .B1(new_n889), .B2(new_n1137), .C1(new_n1014), .C2(new_n869), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1138), .B1(new_n1139), .B2(new_n799), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n751), .B1(new_n1139), .B2(new_n1040), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1140), .B1(new_n1053), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(G390));
  AOI21_X1  g0943(.A(new_n770), .B1(new_n985), .B2(new_n987), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n919), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n766), .A2(new_n875), .A3(new_n725), .A4(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n920), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n961), .B1(new_n1147), .B2(new_n925), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1148), .A2(new_n972), .A3(new_n978), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n959), .A2(new_n962), .B1(new_n960), .B2(new_n926), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n990), .B(new_n1144), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1151), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n772), .A2(new_n793), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1154), .A2(G330), .A3(new_n879), .A4(new_n925), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1153), .A2(new_n1149), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n981), .A2(new_n979), .A3(new_n984), .ZN(new_n1158));
  AOI21_X1  g0958(.A(KEYINPUT104), .B1(new_n772), .B2(new_n986), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n990), .B(G330), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n794), .A2(new_n879), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n989), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g0963(.A(G330), .B(new_n879), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n989), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1155), .A2(new_n1146), .A3(new_n920), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n921), .A2(new_n1163), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1144), .B1(new_n484), .B2(new_n486), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1168), .A2(new_n968), .A3(new_n709), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1157), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1152), .A2(new_n1156), .A3(new_n1170), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(new_n797), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n908), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n413), .B1(G116), .B2(new_n849), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1176), .B1(new_n490), .B2(new_n848), .C1(new_n858), .C2(new_n825), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n897), .B(new_n1177), .C1(G87), .C2(new_n840), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n832), .A2(new_n863), .B1(new_n205), .B2(new_n837), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G107), .B2(new_n833), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n839), .A2(new_n428), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT53), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n834), .A2(new_n892), .B1(new_n842), .B2(new_n208), .ZN(new_n1183));
  INV_X1    g0983(.A(G128), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n832), .A2(new_n1184), .B1(new_n826), .B2(new_n837), .ZN(new_n1185));
  INV_X1    g0985(.A(G132), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n413), .B1(new_n850), .B2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT54), .B(G143), .ZN(new_n1188));
  INV_X1    g0988(.A(G125), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n848), .A2(new_n1188), .B1(new_n825), .B2(new_n1189), .ZN(new_n1190));
  NOR4_X1   g0990(.A1(new_n1183), .A2(new_n1185), .A3(new_n1187), .A4(new_n1190), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1178), .A2(new_n1180), .B1(new_n1182), .B2(new_n1191), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n804), .B1(new_n1100), .B2(new_n1175), .C1(new_n1192), .C2(new_n889), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n959), .A2(new_n962), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1193), .B1(new_n1194), .B2(new_n810), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1157), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1195), .B1(new_n1196), .B2(new_n800), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1174), .A2(new_n1197), .ZN(G378));
  OR2_X1    g0998(.A1(new_n965), .A2(new_n966), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n770), .B1(new_n993), .B2(new_n994), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n992), .A2(new_n1200), .A3(KEYINPUT119), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n435), .A2(new_n933), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n450), .B(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT118), .ZN(new_n1204));
  XOR2_X1   g1004(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1205));
  XNOR2_X1  g1005(.A(new_n1204), .B(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1201), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT119), .B1(new_n992), .B2(new_n1200), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n992), .A2(new_n1200), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT119), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1211), .A2(new_n1212), .A3(new_n1206), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1199), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1216), .A2(new_n1201), .A3(new_n1207), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1215), .A2(new_n1217), .A3(new_n967), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1214), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1207), .A2(new_n810), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n801), .B1(new_n1175), .B2(G50), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT117), .Z(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  AOI211_X1 g1023(.A(G33), .B(G41), .C1(new_n845), .C2(G124), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n826), .B2(new_n842), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n850), .A2(new_n1184), .B1(new_n839), .B2(new_n1188), .ZN(new_n1226));
  XOR2_X1   g1026(.A(new_n1226), .B(KEYINPUT116), .Z(new_n1227));
  OAI22_X1  g1027(.A1(new_n832), .A2(new_n1189), .B1(new_n848), .B2(new_n892), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n834), .A2(new_n1186), .B1(new_n428), .B2(new_n837), .ZN(new_n1229));
  OR3_X1    g1029(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1225), .B1(new_n1230), .B2(KEYINPUT59), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(KEYINPUT59), .B2(new_n1230), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n842), .A2(new_n201), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(G116), .B2(new_n831), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n490), .B2(new_n834), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n348), .B(new_n279), .C1(new_n825), .C2(new_n863), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n850), .A2(new_n465), .B1(new_n452), .B2(new_n848), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1098), .B1(new_n202), .B2(new_n837), .ZN(new_n1238));
  OR4_X1    g1038(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT58), .ZN(new_n1240));
  OR2_X1    g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n208), .B1(G33), .B2(G41), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n279), .B2(new_n348), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1232), .A2(new_n1241), .A3(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1223), .B1(new_n1246), .B2(new_n809), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1219), .A2(new_n800), .B1(new_n1220), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT57), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1168), .A2(new_n968), .A3(new_n709), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1249), .B1(new_n1173), .B2(new_n1250), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1215), .A2(new_n1217), .A3(new_n967), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n967), .B1(new_n1217), .B2(new_n1215), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1251), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n797), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1173), .A2(new_n1250), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT57), .B1(new_n1219), .B2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1248), .B1(new_n1255), .B2(new_n1257), .ZN(G375));
  INV_X1    g1058(.A(new_n1029), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1171), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n925), .A2(new_n811), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(KEYINPUT120), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n845), .A2(G303), .B1(new_n849), .B2(G283), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1264), .B(new_n279), .C1(new_n465), .C2(new_n848), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1099), .B(new_n1265), .C1(G116), .C2(new_n833), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n832), .A2(new_n858), .B1(new_n842), .B2(new_n205), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(G97), .B2(new_n840), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n837), .A2(new_n208), .B1(new_n839), .B2(new_n826), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(G132), .B2(new_n831), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n834), .A2(new_n1188), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n850), .A2(new_n892), .B1(new_n848), .B2(new_n428), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n413), .B1(new_n825), .B2(new_n1184), .ZN(new_n1273));
  NOR4_X1   g1073(.A1(new_n1271), .A2(new_n1233), .A3(new_n1272), .A4(new_n1273), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1266), .A2(new_n1268), .B1(new_n1270), .B2(new_n1274), .ZN(new_n1275));
  OAI221_X1 g1075(.A(new_n804), .B1(G68), .B2(new_n1175), .C1(new_n1275), .C2(new_n889), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1263), .A2(new_n1276), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1144), .A2(new_n990), .B1(new_n989), .B2(new_n1161), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n882), .A2(new_n920), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n925), .B1(new_n1144), .B2(new_n879), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1155), .A2(new_n1146), .A3(new_n920), .ZN(new_n1281));
  OAI22_X1  g1081(.A1(new_n1278), .A2(new_n1279), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1277), .B1(new_n1282), .B2(new_n800), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1261), .A2(new_n1283), .ZN(G381));
  INV_X1    g1084(.A(G378), .ZN(new_n1285));
  NOR4_X1   g1085(.A1(G381), .A2(G384), .A3(G396), .A4(G393), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1285), .A2(new_n1142), .A3(new_n1286), .ZN(new_n1287));
  OR3_X1    g1087(.A1(G375), .A2(new_n1287), .A3(G387), .ZN(G407));
  NAND2_X1  g1088(.A1(new_n720), .A2(G213), .ZN(new_n1289));
  XOR2_X1   g1089(.A(new_n1289), .B(KEYINPUT121), .Z(new_n1290));
  NAND2_X1  g1090(.A1(new_n1285), .A2(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(G407), .B(G213), .C1(G375), .C2(new_n1291), .ZN(G409));
  OAI211_X1 g1092(.A(G378), .B(new_n1248), .C1(new_n1255), .C2(new_n1257), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1259), .B(new_n1256), .C1(new_n1252), .C2(new_n1253), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n800), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1220), .A2(new_n1247), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1294), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1285), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1293), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT122), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT60), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1301), .B1(new_n1282), .B2(new_n1250), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1163), .A2(new_n921), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1169), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1300), .B1(new_n1302), .B2(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(KEYINPUT60), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1307), .A2(KEYINPUT122), .A3(new_n1260), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n751), .B1(new_n1305), .B2(KEYINPUT60), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1306), .A2(new_n1308), .A3(new_n1309), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1310), .A2(G384), .A3(new_n1283), .ZN(new_n1311));
  AOI21_X1  g1111(.A(G384), .B1(new_n1310), .B2(new_n1283), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1299), .A2(new_n1289), .A3(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT63), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1289), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1317), .B1(new_n1293), .B2(new_n1298), .ZN(new_n1318));
  OAI211_X1 g1118(.A(G2897), .B(new_n1290), .C1(new_n1311), .C2(new_n1312), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT123), .ZN(new_n1320));
  INV_X1    g1120(.A(G2897), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1289), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1322), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT124), .B1(new_n1313), .B2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT124), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1323), .ZN(new_n1326));
  NOR4_X1   g1126(.A1(new_n1311), .A2(new_n1312), .A3(new_n1325), .A4(new_n1326), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1319), .B1(new_n1324), .B2(new_n1327), .ZN(new_n1328));
  OR2_X1    g1128(.A1(new_n1318), .A2(new_n1328), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1055), .A2(KEYINPUT125), .A3(G390), .A4(new_n1081), .ZN(new_n1330));
  XOR2_X1   g1130(.A(G393), .B(G396), .Z(new_n1331));
  AND2_X1   g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1025), .B1(new_n737), .B2(new_n1026), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1023), .A2(new_n1024), .A3(new_n1027), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1043), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1042), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1337));
  NOR3_X1   g1137(.A1(new_n1336), .A2(new_n1337), .A3(new_n1139), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n795), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1259), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1335), .B1(new_n1340), .B2(new_n799), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1081), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1142), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT125), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1055), .A2(new_n1081), .A3(G390), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1343), .A2(new_n1344), .A3(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1331), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1343), .A2(new_n1345), .A3(new_n1347), .ZN(new_n1348));
  AOI22_X1  g1148(.A1(new_n1332), .A2(new_n1346), .B1(new_n1348), .B2(KEYINPUT126), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT126), .ZN(new_n1350));
  NAND4_X1  g1150(.A1(new_n1343), .A2(new_n1345), .A3(new_n1350), .A4(new_n1347), .ZN(new_n1351));
  AOI21_X1  g1151(.A(KEYINPUT61), .B1(new_n1349), .B2(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1290), .B1(new_n1293), .B2(new_n1298), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1353), .A2(KEYINPUT63), .A3(new_n1313), .ZN(new_n1354));
  NAND4_X1  g1154(.A1(new_n1316), .A2(new_n1329), .A3(new_n1352), .A4(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT61), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1356), .B1(new_n1353), .B2(new_n1328), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT62), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1314), .A2(new_n1358), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1353), .A2(KEYINPUT62), .A3(new_n1313), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1357), .B1(new_n1359), .B2(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1332), .A2(new_n1346), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1348), .A2(KEYINPUT126), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1362), .A2(new_n1363), .A3(new_n1351), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1355), .B1(new_n1361), .B2(new_n1364), .ZN(G405));
  INV_X1    g1165(.A(KEYINPUT127), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1364), .A2(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(G375), .A2(new_n1285), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1368), .A2(new_n1293), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1369), .A2(new_n1313), .ZN(new_n1370));
  NAND4_X1  g1170(.A1(new_n1362), .A2(new_n1363), .A3(KEYINPUT127), .A4(new_n1351), .ZN(new_n1371));
  OAI211_X1 g1171(.A(new_n1368), .B(new_n1293), .C1(new_n1312), .C2(new_n1311), .ZN(new_n1372));
  AND4_X1   g1172(.A1(new_n1367), .A2(new_n1370), .A3(new_n1371), .A4(new_n1372), .ZN(new_n1373));
  AOI22_X1  g1173(.A1(new_n1367), .A2(new_n1371), .B1(new_n1370), .B2(new_n1372), .ZN(new_n1374));
  NOR2_X1   g1174(.A1(new_n1373), .A2(new_n1374), .ZN(G402));
endmodule


