//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  INV_X1    g0007(.A(G244), .ZN(new_n208));
  INV_X1    g0008(.A(G107), .ZN(new_n209));
  INV_X1    g0009(.A(G264), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT65), .ZN(new_n213));
  AOI211_X1 g0013(.A(new_n211), .B(new_n213), .C1(G50), .C2(G226), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G116), .A2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n214), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AND2_X1   g0018(.A1(G68), .A2(G238), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n206), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT1), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT64), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT64), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n224), .A2(G1), .A3(G13), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G20), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n206), .A2(G13), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT0), .Z(new_n232));
  NOR3_X1   g0032(.A1(new_n221), .A2(new_n229), .A3(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT66), .B(G107), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NOR2_X1   g0049(.A1(G226), .A2(G1698), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n250), .B1(new_n217), .B2(G1698), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  AOI22_X1  g0052(.A1(new_n251), .A2(new_n252), .B1(G33), .B2(G97), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n226), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(KEYINPUT70), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n255), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G97), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n217), .A2(G1698), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(G226), .B2(G1698), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n258), .B1(new_n260), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT70), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n257), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n269), .B1(G41), .B2(G45), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n254), .A2(G1), .A3(G13), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n270), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n272), .B1(new_n275), .B2(G238), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n256), .A2(new_n268), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT13), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT13), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n256), .A2(new_n268), .A3(new_n279), .A4(new_n276), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G190), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G13), .ZN(new_n284));
  INV_X1    g0084(.A(G20), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n284), .A2(new_n285), .A3(G1), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  OR3_X1    g0087(.A1(new_n287), .A2(KEYINPUT12), .A3(G68), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT12), .B1(new_n287), .B2(G68), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n223), .A2(new_n225), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n291), .B1(new_n269), .B2(G20), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n288), .A2(new_n289), .B1(new_n292), .B2(G68), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n285), .A2(G33), .ZN(new_n294));
  OAI22_X1  g0094(.A1(new_n294), .A2(new_n207), .B1(new_n285), .B2(G68), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n295), .A2(KEYINPUT71), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(KEYINPUT71), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G20), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n296), .B(new_n297), .C1(new_n202), .C2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT11), .ZN(new_n301));
  AND3_X1   g0101(.A1(new_n300), .A2(new_n301), .A3(new_n291), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(new_n300), .B2(new_n291), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n293), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G200), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(new_n278), .B2(new_n280), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n283), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n281), .A2(G169), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT72), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT14), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n278), .A2(G179), .A3(new_n280), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT73), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n313), .A2(new_n314), .B1(KEYINPUT72), .B2(KEYINPUT14), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n278), .A2(KEYINPUT73), .A3(G179), .A4(new_n280), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n281), .A2(new_n309), .A3(new_n310), .A4(G169), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n312), .A2(new_n315), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n307), .B1(new_n318), .B2(new_n304), .ZN(new_n319));
  NOR2_X1   g0119(.A1(G222), .A2(G1698), .ZN(new_n320));
  INV_X1    g0120(.A(G1698), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(G223), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n252), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n257), .B(new_n323), .C1(G77), .C2(new_n252), .ZN(new_n324));
  INV_X1    g0124(.A(new_n272), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n275), .A2(G226), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT69), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n328), .A2(G190), .B1(new_n329), .B2(KEYINPUT10), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n292), .A2(G50), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT8), .B(G58), .ZN(new_n332));
  INV_X1    g0132(.A(G150), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n332), .A2(new_n294), .B1(new_n333), .B2(new_n299), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(G20), .B2(new_n203), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n223), .A2(new_n225), .A3(new_n290), .ZN(new_n336));
  OAI221_X1 g0136(.A(new_n331), .B1(G50), .B2(new_n287), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT9), .ZN(new_n338));
  XOR2_X1   g0138(.A(KEYINPUT68), .B(G200), .Z(new_n339));
  AOI22_X1  g0139(.A1(new_n337), .A2(new_n338), .B1(new_n339), .B2(new_n327), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n330), .B(new_n340), .C1(new_n338), .C2(new_n337), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n329), .A2(KEYINPUT10), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G179), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n328), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G169), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n327), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n345), .A2(new_n337), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G20), .A2(G77), .ZN(new_n349));
  XOR2_X1   g0149(.A(KEYINPUT15), .B(G87), .Z(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n349), .B1(new_n332), .B2(new_n299), .C1(new_n294), .C2(new_n351), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(new_n291), .B1(G77), .B2(new_n292), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(G77), .B2(new_n287), .ZN(new_n354));
  NOR2_X1   g0154(.A1(G232), .A2(G1698), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n321), .A2(G238), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n252), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT67), .B(G107), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n257), .B(new_n357), .C1(new_n252), .C2(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n359), .B(new_n325), .C1(new_n208), .C2(new_n274), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n346), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n354), .B(new_n361), .C1(G179), .C2(new_n360), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n319), .A2(new_n343), .A3(new_n348), .A4(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT18), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n261), .A2(KEYINPUT74), .A3(G33), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT74), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(KEYINPUT3), .B2(new_n263), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n365), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT7), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT75), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT75), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT7), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n369), .A2(new_n285), .A3(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT74), .B1(new_n261), .B2(G33), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n262), .ZN(new_n377));
  AOI21_X1  g0177(.A(G20), .B1(new_n377), .B2(new_n365), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n375), .B(G68), .C1(new_n370), .C2(new_n378), .ZN(new_n379));
  XNOR2_X1  g0179(.A(G58), .B(G68), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n380), .A2(G20), .B1(G159), .B2(new_n298), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(KEYINPUT16), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT16), .ZN(new_n383));
  INV_X1    g0183(.A(G68), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n374), .B1(new_n252), .B2(G20), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n285), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n381), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n383), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n382), .A2(new_n389), .A3(new_n291), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n287), .A2(new_n332), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n292), .B2(new_n332), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  OR2_X1    g0193(.A1(G223), .A2(G1698), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n321), .A2(G226), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n377), .A2(new_n365), .A3(new_n394), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G33), .A2(G87), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n257), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n325), .B1(new_n274), .B2(new_n217), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(G169), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n255), .B1(new_n396), .B2(new_n397), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n403), .A2(G179), .A3(new_n400), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT76), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n399), .A2(new_n344), .A3(new_n401), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT76), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n346), .B1(new_n403), .B2(new_n400), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n364), .B1(new_n393), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n390), .A2(new_n392), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n412), .A2(KEYINPUT18), .A3(new_n405), .A4(new_n409), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n399), .A2(new_n282), .A3(new_n401), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n305), .B1(new_n403), .B2(new_n400), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(KEYINPUT77), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT77), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n399), .A2(new_n418), .A3(new_n282), .A4(new_n401), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n390), .A2(new_n417), .A3(new_n419), .A4(new_n392), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n420), .B(KEYINPUT17), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n354), .B1(new_n360), .B2(new_n339), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n282), .B2(new_n360), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n414), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n363), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(G45), .ZN(new_n426));
  NOR3_X1   g0226(.A1(new_n426), .A2(new_n271), .A3(G1), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n273), .B(G250), .C1(G1), .C2(new_n426), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G116), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n208), .A2(G1698), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(G238), .B2(G1698), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n430), .B1(new_n369), .B2(new_n432), .ZN(new_n433));
  AOI211_X1 g0233(.A(new_n427), .B(new_n429), .C1(new_n433), .C2(new_n257), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n344), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n257), .ZN(new_n436));
  INV_X1    g0236(.A(new_n427), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(new_n428), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n346), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n377), .A2(new_n285), .A3(G68), .A4(new_n365), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT19), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n285), .B1(new_n258), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G87), .ZN(new_n443));
  INV_X1    g0243(.A(G97), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n442), .B1(new_n358), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n441), .B1(new_n294), .B2(new_n444), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n440), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n448), .A2(new_n291), .B1(new_n286), .B2(new_n351), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n269), .A2(G33), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n336), .A2(new_n287), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n350), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n435), .A2(new_n439), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n339), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n427), .B1(new_n433), .B2(new_n257), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n455), .B1(new_n456), .B2(new_n428), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n448), .A2(new_n291), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n351), .A2(new_n286), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n451), .A2(G87), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT81), .B1(new_n438), .B2(new_n282), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT81), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n434), .A2(new_n464), .A3(G190), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n462), .A2(KEYINPUT80), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT80), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n457), .B2(new_n461), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n454), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n321), .A2(G244), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n365), .B(new_n471), .C1(new_n367), .C2(new_n368), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT4), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  INV_X1    g0275(.A(G250), .ZN(new_n476));
  OAI22_X1  g0276(.A1(new_n470), .A2(new_n473), .B1(new_n476), .B2(new_n321), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n252), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n474), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n257), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT5), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G41), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT78), .B1(new_n481), .B2(G41), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT78), .ZN(new_n484));
  INV_X1    g0284(.A(G41), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT5), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n427), .A2(new_n482), .A3(new_n483), .A4(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n269), .B(G45), .C1(new_n485), .C2(KEYINPUT5), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n481), .A2(G41), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n273), .B(G257), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n480), .A2(G190), .A3(new_n487), .A4(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT79), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n490), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n479), .B2(new_n257), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n495), .A2(KEYINPUT79), .A3(G190), .A4(new_n487), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT6), .ZN(new_n498));
  AND2_X1   g0298(.A1(G97), .A2(G107), .ZN(new_n499));
  NOR2_X1   g0299(.A1(G97), .A2(G107), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n209), .A2(KEYINPUT6), .A3(G97), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n503), .A2(new_n285), .B1(new_n207), .B2(new_n299), .ZN(new_n504));
  INV_X1    g0304(.A(new_n358), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n505), .B1(new_n385), .B2(new_n386), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n291), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n286), .A2(new_n444), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n336), .A2(new_n287), .A3(new_n450), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(new_n444), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n507), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n480), .A2(new_n487), .A3(new_n490), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n512), .B1(G200), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n265), .A2(new_n285), .B1(new_n371), .B2(new_n373), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n252), .A2(new_n370), .A3(G20), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n358), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n501), .A2(new_n502), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n518), .A2(G20), .B1(G77), .B2(new_n298), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n510), .B1(new_n520), .B2(new_n291), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n346), .A2(new_n513), .B1(new_n521), .B2(new_n508), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n495), .A2(new_n344), .A3(new_n487), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n497), .A2(new_n514), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(G257), .A2(G1698), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n525), .B1(new_n210), .B2(G1698), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n377), .A2(new_n526), .A3(new_n365), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n265), .A2(G303), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n255), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n273), .B(G270), .C1(new_n488), .C2(new_n489), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n487), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(G169), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n475), .B(new_n285), .C1(G33), .C2(new_n444), .ZN(new_n533));
  INV_X1    g0333(.A(G116), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G20), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n291), .A2(KEYINPUT20), .A3(new_n533), .A4(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT82), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n533), .A2(new_n535), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n539), .A2(KEYINPUT82), .A3(KEYINPUT20), .A4(new_n291), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n291), .A2(new_n533), .A3(new_n535), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT20), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n541), .A2(KEYINPUT83), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT83), .B1(new_n541), .B2(new_n542), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n538), .B(new_n540), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n287), .A2(G116), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n509), .B2(new_n534), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n532), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(KEYINPUT21), .B(G169), .C1(new_n529), .C2(new_n531), .ZN(new_n551));
  INV_X1    g0351(.A(new_n531), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n261), .A2(KEYINPUT74), .A3(G33), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(new_n262), .B2(new_n376), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n554), .A2(new_n526), .B1(G303), .B2(new_n265), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n552), .B(G179), .C1(new_n555), .C2(new_n255), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n541), .A2(new_n542), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT83), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n541), .A2(KEYINPUT83), .A3(new_n542), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n538), .A2(new_n540), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n548), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI22_X1  g0364(.A1(new_n550), .A2(KEYINPUT21), .B1(new_n557), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n529), .A2(new_n531), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G190), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n305), .B2(new_n566), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n545), .A2(new_n549), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n469), .A2(new_n524), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT86), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n443), .A2(G20), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n377), .A2(KEYINPUT22), .A3(new_n365), .A4(new_n574), .ZN(new_n575));
  NOR3_X1   g0375(.A1(new_n285), .A2(KEYINPUT23), .A3(G107), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n262), .A3(new_n264), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT22), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(KEYINPUT23), .B1(new_n358), .B2(new_n285), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n430), .A2(G20), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n575), .A2(new_n579), .A3(new_n580), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT24), .ZN(new_n584));
  AOI211_X1 g0384(.A(new_n576), .B(new_n581), .C1(new_n577), .C2(new_n578), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT24), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n585), .A2(new_n586), .A3(new_n580), .A4(new_n575), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n291), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT25), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n287), .B2(G107), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n286), .A2(KEYINPUT25), .A3(new_n209), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n451), .A2(G107), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n476), .A2(new_n321), .ZN(new_n595));
  OR2_X1    g0395(.A1(new_n321), .A2(G257), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n377), .A2(new_n365), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  XOR2_X1   g0397(.A(KEYINPUT84), .B(G294), .Z(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G33), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n257), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n273), .B(G264), .C1(new_n488), .C2(new_n489), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n601), .A2(new_n602), .A3(new_n487), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G169), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n255), .B1(new_n597), .B2(new_n599), .ZN(new_n605));
  INV_X1    g0405(.A(new_n602), .ZN(new_n606));
  INV_X1    g0406(.A(new_n487), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(G179), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT85), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n604), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n606), .B1(new_n600), .B2(new_n257), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n346), .B1(new_n612), .B2(new_n487), .ZN(new_n613));
  NOR4_X1   g0413(.A1(new_n605), .A2(new_n344), .A3(new_n606), .A4(new_n607), .ZN(new_n614));
  OAI21_X1  g0414(.A(KEYINPUT85), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n594), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n608), .A2(G190), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n603), .A2(G200), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n589), .A2(new_n593), .A3(new_n617), .A4(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n573), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n616), .A2(new_n573), .A3(new_n619), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n572), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n425), .A2(new_n622), .ZN(G372));
  INV_X1    g0423(.A(new_n348), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n307), .A2(new_n362), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n318), .A2(new_n304), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT89), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT89), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n625), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n421), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n414), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n624), .B1(new_n632), .B2(new_n343), .ZN(new_n633));
  INV_X1    g0433(.A(new_n425), .ZN(new_n634));
  XNOR2_X1  g0434(.A(new_n454), .B(KEYINPUT87), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT26), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n513), .A2(new_n346), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n637), .A2(new_n512), .A3(new_n523), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT21), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n564), .B2(new_n532), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n336), .B1(new_n584), .B2(new_n587), .ZN(new_n641));
  INV_X1    g0441(.A(new_n593), .ZN(new_n642));
  OAI22_X1  g0442(.A1(new_n641), .A2(new_n642), .B1(new_n613), .B2(new_n614), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n551), .A2(new_n556), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n569), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n640), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n638), .B1(new_n646), .B2(new_n619), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n497), .A2(new_n514), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n463), .A2(new_n465), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n346), .A2(new_n438), .B1(new_n449), .B2(new_n452), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n649), .A2(new_n462), .B1(new_n650), .B2(new_n435), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n636), .B1(new_n647), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n438), .A2(new_n339), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n654), .A2(KEYINPUT80), .A3(new_n449), .A4(new_n460), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n649), .A2(new_n655), .A3(new_n468), .ZN(new_n656));
  INV_X1    g0456(.A(new_n454), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(new_n638), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g0458(.A(KEYINPUT88), .B(KEYINPUT26), .Z(new_n659));
  OR2_X1    g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n635), .B1(new_n653), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n633), .B1(new_n634), .B2(new_n661), .ZN(G369));
  XOR2_X1   g0462(.A(KEYINPUT90), .B(KEYINPUT27), .Z(new_n663));
  NOR3_X1   g0463(.A1(new_n284), .A2(G1), .A3(G20), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G213), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n670), .B1(new_n589), .B2(new_n593), .ZN(new_n671));
  OR3_X1    g0471(.A1(new_n621), .A2(new_n620), .A3(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n616), .A2(new_n670), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n672), .A2(KEYINPUT91), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT91), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n621), .A2(new_n620), .A3(new_n671), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n676), .B1(new_n677), .B2(new_n673), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n564), .A2(new_n670), .ZN(new_n681));
  MUX2_X1   g0481(.A(new_n571), .B(new_n565), .S(new_n681), .Z(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n565), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(new_n669), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n675), .B2(new_n678), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n643), .A2(new_n669), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n685), .A2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n230), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n358), .A2(G116), .A3(new_n445), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G1), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n228), .B2(new_n695), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n658), .A2(new_n659), .ZN(new_n700));
  AOI22_X1  g0500(.A1(new_n589), .A2(new_n593), .B1(new_n604), .B2(new_n609), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n619), .B1(new_n565), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n638), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n648), .A2(new_n651), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n700), .B1(new_n706), .B2(new_n636), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n670), .B1(new_n707), .B2(new_n635), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(KEYINPUT29), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n651), .A2(KEYINPUT26), .A3(new_n638), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT94), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n658), .A2(new_n711), .A3(new_n659), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n711), .B1(new_n658), .B2(new_n659), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n710), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n686), .A2(new_n616), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n715), .A2(new_n619), .A3(new_n524), .A4(new_n651), .ZN(new_n716));
  INV_X1    g0516(.A(new_n635), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n669), .B1(new_n714), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT29), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n709), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n621), .A2(new_n620), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n469), .A2(new_n524), .A3(new_n571), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(new_n724), .A3(new_n670), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n495), .A2(G179), .A3(new_n566), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n608), .A2(new_n434), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n603), .A2(new_n438), .ZN(new_n730));
  INV_X1    g0530(.A(new_n556), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n730), .A2(KEYINPUT30), .A3(new_n495), .A4(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT92), .ZN(new_n733));
  AOI21_X1  g0533(.A(G179), .B1(new_n434), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n552), .B1(new_n555), .B2(new_n255), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n438), .A2(KEYINPUT92), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n734), .A2(new_n513), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n729), .B(new_n732), .C1(new_n737), .C2(new_n608), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n669), .ZN(new_n739));
  AOI21_X1  g0539(.A(KEYINPUT31), .B1(new_n738), .B2(new_n669), .ZN(new_n740));
  OAI21_X1  g0540(.A(KEYINPUT93), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n740), .A2(KEYINPUT93), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n725), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G330), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n722), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n699), .B1(new_n746), .B2(G1), .ZN(G364));
  OR2_X1    g0547(.A1(new_n682), .A2(G330), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n284), .A2(G20), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G45), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n695), .A2(G1), .A3(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n748), .A2(new_n683), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n226), .B1(new_n285), .B2(G169), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT95), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n285), .A2(new_n344), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n282), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(KEYINPUT97), .A3(new_n305), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(KEYINPUT97), .B1(new_n757), .B2(new_n305), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n756), .A2(new_n305), .A3(G190), .ZN(new_n763));
  XNOR2_X1  g0563(.A(KEYINPUT33), .B(G317), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n762), .A2(G322), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT100), .Z(new_n766));
  INV_X1    g0566(.A(new_n757), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n305), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G326), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n285), .A2(G179), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G190), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n774), .A2(KEYINPUT98), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(KEYINPUT98), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G329), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n339), .A2(new_n772), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n282), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G303), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n265), .B1(new_n777), .B2(new_n778), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n766), .A2(new_n771), .A3(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G283), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n779), .A2(G190), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n598), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n282), .A2(G179), .A3(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n285), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n784), .B1(new_n785), .B2(new_n787), .C1(new_n788), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n755), .A2(new_n773), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n791), .B1(G311), .B2(new_n793), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT101), .Z(new_n795));
  INV_X1    g0595(.A(G159), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n777), .A2(new_n796), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT32), .Z(new_n798));
  NAND2_X1  g0598(.A1(new_n786), .A2(G107), .ZN(new_n799));
  INV_X1    g0599(.A(new_n790), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n800), .A2(G97), .B1(new_n793), .B2(G77), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n799), .B(new_n801), .C1(new_n761), .C2(new_n216), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n780), .A2(G87), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT99), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n803), .A2(new_n804), .A3(new_n252), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n804), .B1(new_n803), .B2(new_n252), .ZN(new_n807));
  NOR4_X1   g0607(.A1(new_n798), .A2(new_n802), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n763), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n808), .B1(new_n202), .B2(new_n769), .C1(new_n384), .C2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n754), .B1(new_n795), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n754), .ZN(new_n812));
  NOR2_X1   g0612(.A1(G13), .A2(G33), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(G20), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT96), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n252), .A2(G355), .A3(new_n230), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n554), .A2(new_n693), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n248), .B2(new_n426), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n228), .A2(G45), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n818), .B1(G116), .B2(new_n230), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n811), .B1(new_n817), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n815), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n682), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n752), .B1(new_n825), .B2(new_n751), .ZN(G396));
  NOR2_X1   g0626(.A1(new_n362), .A2(new_n669), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n354), .A2(new_n669), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n423), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n827), .B1(new_n829), .B2(new_n362), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n670), .B(new_n830), .C1(new_n707), .C2(new_n635), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(KEYINPUT103), .ZN(new_n832));
  INV_X1    g0632(.A(new_n830), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n708), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n832), .B(new_n834), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n835), .A2(new_n744), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n744), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n836), .A2(new_n751), .A3(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n777), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n762), .A2(G294), .B1(G311), .B2(new_n839), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n840), .B(new_n265), .C1(new_n785), .C2(new_n809), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(G116), .B2(new_n793), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n768), .A2(G303), .B1(G97), .B2(new_n800), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n786), .A2(G87), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n780), .A2(G107), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n842), .A2(new_n843), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n768), .A2(G137), .B1(G150), .B2(new_n763), .ZN(new_n847));
  INV_X1    g0647(.A(G143), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n847), .B1(new_n796), .B2(new_n792), .C1(new_n761), .C2(new_n848), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT34), .Z(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G50), .B2(new_n780), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n839), .A2(G132), .B1(G58), .B2(new_n800), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n851), .B(new_n852), .C1(new_n384), .C2(new_n787), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n846), .B1(new_n853), .B2(new_n369), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n812), .ZN(new_n855));
  INV_X1    g0655(.A(new_n751), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n833), .A2(new_n813), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n754), .A2(new_n814), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT102), .Z(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n207), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n855), .A2(new_n856), .A3(new_n857), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n838), .A2(new_n861), .ZN(G384));
  INV_X1    g0662(.A(KEYINPUT40), .ZN(new_n863));
  INV_X1    g0663(.A(new_n392), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n382), .A2(new_n291), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n379), .A2(new_n381), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n383), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n864), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n667), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n405), .B2(new_n409), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n420), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT37), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT105), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n410), .A2(new_n667), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n412), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT37), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(new_n876), .A3(new_n420), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT105), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n871), .A2(new_n878), .A3(KEYINPUT37), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n873), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n414), .A2(new_n421), .ZN(new_n881));
  INV_X1    g0681(.A(new_n868), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(new_n869), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n880), .A2(KEYINPUT38), .A3(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT38), .B1(new_n880), .B2(new_n883), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n307), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n304), .A2(new_n669), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n626), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n318), .A2(new_n304), .A3(new_n669), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR4_X1   g0692(.A1(new_n572), .A2(new_n621), .A3(new_n620), .A4(new_n669), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n738), .A2(new_n669), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT31), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n669), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n892), .B(new_n830), .C1(new_n893), .C2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n863), .B1(new_n887), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n725), .A2(new_n896), .A3(new_n897), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT38), .ZN(new_n902));
  AOI211_X1 g0702(.A(new_n393), .B(new_n667), .C1(new_n414), .C2(new_n421), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n870), .A2(new_n393), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT106), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT37), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n875), .A2(new_n420), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n875), .A2(new_n905), .A3(KEYINPUT37), .A4(new_n420), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n902), .B1(new_n903), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n884), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n898), .B1(new_n622), .B2(new_n670), .ZN(new_n913));
  INV_X1    g0713(.A(new_n889), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n914), .B(new_n307), .C1(new_n318), .C2(new_n304), .ZN(new_n915));
  INV_X1    g0715(.A(new_n891), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n830), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n912), .A2(new_n918), .A3(KEYINPUT40), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n900), .A2(new_n425), .A3(new_n901), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n880), .A2(new_n883), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n902), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n899), .B1(new_n922), .B2(new_n884), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n919), .B(G330), .C1(new_n923), .C2(KEYINPUT40), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n901), .A2(G330), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n425), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n920), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT107), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n425), .B1(new_n709), .B2(new_n721), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n633), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n930), .B(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n922), .A2(new_n884), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT104), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n653), .A2(new_n660), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n669), .B1(new_n936), .B2(new_n717), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n935), .B(new_n827), .C1(new_n937), .C2(new_n830), .ZN(new_n938));
  INV_X1    g0738(.A(new_n827), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT104), .B1(new_n831), .B2(new_n939), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n934), .B(new_n892), .C1(new_n938), .C2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT39), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n912), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n922), .A2(KEYINPUT39), .A3(new_n884), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n626), .A2(new_n669), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n411), .A2(new_n413), .A3(new_n667), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n941), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n933), .B(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n269), .B2(new_n749), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n534), .B1(new_n518), .B2(KEYINPUT35), .ZN(new_n951));
  INV_X1    g0751(.A(new_n227), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n951), .B(new_n952), .C1(KEYINPUT35), .C2(new_n518), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT36), .ZN(new_n954));
  OAI21_X1  g0754(.A(G77), .B1(new_n216), .B2(new_n384), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n955), .A2(new_n228), .B1(G50), .B2(new_n384), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(G1), .A3(new_n284), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n950), .A2(new_n954), .A3(new_n957), .ZN(G367));
  INV_X1    g0758(.A(new_n689), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n512), .A2(new_n669), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n524), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(new_n638), .B2(new_n669), .ZN(new_n962));
  OAI21_X1  g0762(.A(KEYINPUT42), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n461), .A2(new_n669), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n651), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n717), .B2(new_n964), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n967));
  INV_X1    g0767(.A(new_n961), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n703), .B1(new_n968), .B2(new_n616), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n670), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT42), .ZN(new_n971));
  INV_X1    g0771(.A(new_n962), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n689), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n963), .A2(new_n967), .A3(new_n970), .A4(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT108), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n685), .A2(new_n962), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n963), .A2(new_n970), .A3(new_n973), .ZN(new_n978));
  INV_X1    g0778(.A(new_n967), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n976), .A2(new_n977), .A3(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n977), .B1(new_n976), .B2(new_n981), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n694), .B(KEYINPUT41), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n690), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n959), .A2(new_n988), .A3(new_n972), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(KEYINPUT109), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT109), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n691), .A2(new_n991), .A3(new_n972), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n990), .A2(KEYINPUT45), .A3(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT45), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n991), .B1(new_n691), .B2(new_n972), .ZN(new_n995));
  NOR4_X1   g0795(.A1(new_n689), .A2(KEYINPUT109), .A3(new_n690), .A4(new_n962), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n962), .B1(new_n689), .B2(new_n690), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT44), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n993), .A2(new_n997), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n684), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n680), .A2(new_n688), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n1003), .A2(new_n959), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n683), .A2(KEYINPUT110), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n683), .B(KEYINPUT110), .Z(new_n1007));
  OAI21_X1  g0807(.A(new_n1006), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1008), .A2(new_n745), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n993), .A2(new_n997), .A3(new_n1000), .A4(new_n685), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1002), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n987), .B1(new_n1011), .B2(new_n746), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n750), .A2(G1), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n985), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n819), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n816), .B1(new_n230), .B2(new_n351), .C1(new_n240), .C2(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n762), .A2(G303), .B1(new_n358), .B2(new_n800), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1017), .B(new_n369), .C1(new_n785), .C2(new_n792), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n598), .B2(new_n763), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n786), .A2(G97), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n780), .A2(G116), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT46), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n839), .A2(G317), .B1(new_n768), .B2(G311), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n768), .A2(G143), .B1(G68), .B2(new_n800), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n761), .B2(new_n333), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT111), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n780), .A2(G58), .B1(G50), .B2(new_n793), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n786), .A2(G77), .B1(G159), .B2(new_n763), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1027), .A2(new_n252), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(G137), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n777), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1024), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT47), .Z(new_n1034));
  OAI211_X1 g0834(.A(new_n856), .B(new_n1016), .C1(new_n1034), .C2(new_n754), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT112), .Z(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n824), .B2(new_n966), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1014), .A2(new_n1037), .ZN(G387));
  AOI22_X1  g0838(.A1(new_n763), .A2(G311), .B1(G303), .B2(new_n793), .ZN(new_n1039));
  INV_X1    g0839(.A(G322), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1039), .B1(new_n769), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G317), .B2(new_n762), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT48), .Z(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n785), .B2(new_n790), .C1(new_n788), .C2(new_n781), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT49), .Z(new_n1045));
  OAI221_X1 g0845(.A(new_n369), .B1(new_n777), .B2(new_n770), .C1(new_n787), .C2(new_n534), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(KEYINPUT113), .B(G150), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n839), .A2(new_n1047), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n384), .B2(new_n792), .C1(new_n207), .C2(new_n781), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n554), .B1(new_n809), .B2(new_n332), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n768), .A2(G159), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT114), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1050), .B(new_n1052), .C1(G50), .C2(new_n762), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n351), .A2(new_n790), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1053), .A2(new_n1020), .A3(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n1045), .A2(new_n1046), .B1(new_n1049), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n812), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n680), .A2(new_n815), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n332), .A2(G50), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT50), .ZN(new_n1061));
  AOI21_X1  g0861(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1061), .A2(new_n696), .A3(new_n1062), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n819), .B(new_n1063), .C1(new_n237), .C2(new_n426), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n252), .A2(new_n230), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1064), .B1(G107), .B2(new_n230), .C1(new_n696), .C2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n817), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1058), .A2(new_n856), .A3(new_n1059), .A4(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1013), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1008), .A2(new_n745), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n694), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1068), .B1(new_n1069), .B2(new_n1008), .C1(new_n1071), .C2(new_n1009), .ZN(G393));
  NAND3_X1  g0872(.A1(new_n1002), .A2(new_n1013), .A3(new_n1010), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n751), .B1(new_n962), .B2(new_n815), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n762), .A2(G311), .B1(G317), .B2(new_n768), .ZN(new_n1075));
  XOR2_X1   g0875(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n1076));
  XNOR2_X1  g0876(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(G294), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n265), .B1(new_n792), .B2(new_n1078), .C1(new_n790), .C2(new_n534), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n799), .B1(new_n1040), .B2(new_n777), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1079), .B(new_n1080), .C1(G283), .C2(new_n780), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1077), .B(new_n1081), .C1(new_n782), .C2(new_n809), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n761), .A2(new_n796), .B1(new_n769), .B2(new_n333), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT51), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n369), .B1(new_n763), .B2(G50), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n790), .A2(new_n207), .B1(new_n792), .B2(new_n332), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n780), .B2(G68), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1084), .A2(new_n844), .A3(new_n1085), .A4(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n777), .A2(new_n848), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1082), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n812), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n816), .B1(new_n444), .B2(new_n230), .C1(new_n245), .C2(new_n1015), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1074), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1073), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1002), .A2(new_n1010), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1008), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n746), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n695), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1094), .B1(new_n1098), .B2(new_n1011), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(G390));
  NAND2_X1  g0900(.A1(new_n943), .A2(new_n944), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n813), .ZN(new_n1102));
  INV_X1    g0902(.A(G132), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n761), .A2(new_n1103), .B1(new_n1031), .B2(new_n809), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(G128), .B2(new_n768), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n786), .A2(G50), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n780), .A2(new_n1047), .ZN(new_n1107));
  XOR2_X1   g0907(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1108));
  XNOR2_X1  g0908(.A(new_n1107), .B(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(G125), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n777), .A2(new_n1110), .B1(new_n796), .B2(new_n790), .ZN(new_n1111));
  XOR2_X1   g0911(.A(KEYINPUT54), .B(G143), .Z(new_n1112));
  AOI211_X1 g0912(.A(new_n265), .B(new_n1111), .C1(new_n793), .C2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1105), .A2(new_n1106), .A3(new_n1109), .A4(new_n1113), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n769), .A2(new_n785), .B1(new_n444), .B2(new_n792), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n358), .B2(new_n763), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT117), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1117), .A2(new_n252), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n839), .A2(G294), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n761), .A2(new_n534), .B1(new_n207), .B2(new_n790), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT118), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1118), .A2(new_n803), .A3(new_n1119), .A4(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n787), .A2(new_n384), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1114), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n812), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n859), .A2(new_n332), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1102), .A2(new_n856), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n945), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n829), .A2(new_n362), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n827), .B1(new_n719), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n892), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1128), .B(new_n912), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n743), .A2(G330), .A3(new_n830), .A4(new_n892), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n661), .A2(new_n669), .A3(new_n833), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n935), .B1(new_n1134), .B2(new_n827), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n831), .A2(KEYINPUT104), .A3(new_n939), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n945), .B1(new_n1137), .B2(new_n892), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1101), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1132), .B(new_n1133), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1132), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n892), .B1(new_n938), .B2(new_n940), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n1128), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1141), .B1(new_n1143), .B2(new_n1101), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n918), .A2(G330), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1140), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1127), .B1(new_n1146), .B2(new_n1069), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1131), .B1(new_n744), .B2(new_n833), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n1145), .ZN(new_n1149));
  OAI211_X1 g0949(.A(G330), .B(new_n830), .C1(new_n893), .C2(new_n898), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n1131), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1151), .A2(new_n1133), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1137), .A2(new_n1149), .B1(new_n1152), .B2(new_n1130), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n931), .A2(new_n633), .A3(new_n927), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1140), .B(new_n1155), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1156), .A2(new_n694), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1149), .A2(new_n1137), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1152), .A2(new_n1130), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1154), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1146), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1147), .B1(new_n1157), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(G378));
  NOR2_X1   g0965(.A1(G33), .A2(G41), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1166), .A2(G50), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n554), .B2(G41), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n762), .A2(G128), .B1(G132), .B2(new_n763), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n780), .A2(new_n1112), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n768), .A2(G125), .B1(G137), .B2(new_n793), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G150), .B2(new_n800), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT59), .Z(new_n1174));
  INV_X1    g0974(.A(G124), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1166), .B1(new_n777), .B2(new_n1175), .C1(new_n787), .C2(new_n796), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1168), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n777), .A2(new_n785), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n800), .A2(G68), .B1(new_n793), .B2(new_n350), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n444), .B2(new_n809), .C1(new_n787), .C2(new_n216), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1178), .B(new_n1180), .C1(G107), .C2(new_n762), .ZN(new_n1181));
  AOI211_X1 g0981(.A(G41), .B(new_n554), .C1(new_n780), .C2(G77), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(new_n534), .C2(new_n769), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1183), .B(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n812), .B1(new_n1177), .B2(new_n1185), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1186), .B(KEYINPUT120), .Z(new_n1187));
  NAND2_X1  g0987(.A1(new_n343), .A2(new_n348), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n337), .A2(new_n869), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1188), .B(new_n1189), .ZN(new_n1190));
  XOR2_X1   g0990(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1191));
  XNOR2_X1  g0991(.A(new_n1190), .B(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n813), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n856), .B1(new_n858), .B2(G50), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT121), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1187), .A2(new_n1193), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT122), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n900), .A2(new_n1192), .A3(G330), .A4(new_n919), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1192), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n924), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n948), .A2(new_n1199), .A3(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n948), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1198), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1202), .A2(KEYINPUT122), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1197), .B1(new_n1207), .B2(new_n1013), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1156), .A2(new_n1161), .ZN(new_n1209));
  AOI21_X1  g1009(.A(KEYINPUT57), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT57), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1201), .A2(new_n1199), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n941), .A2(new_n946), .A3(new_n947), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1211), .B1(new_n1214), .B2(new_n1202), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1209), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n694), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1208), .B1(new_n1210), .B2(new_n1217), .ZN(G375));
  NAND2_X1  g1018(.A1(new_n859), .A2(new_n384), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n892), .B2(new_n814), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n839), .A2(G128), .B1(new_n768), .B2(G132), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1221), .B(new_n554), .C1(new_n202), .C2(new_n790), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G159), .B2(new_n780), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n763), .A2(new_n1112), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n762), .A2(G137), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n786), .A2(G58), .B1(G150), .B2(new_n793), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n761), .A2(new_n785), .B1(new_n207), .B2(new_n787), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n252), .B(new_n1228), .C1(G116), .C2(new_n763), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1055), .B1(new_n769), .B2(new_n1078), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n358), .B2(new_n793), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1229), .B(new_n1231), .C1(new_n444), .C2(new_n781), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n777), .A2(new_n782), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1227), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n751), .B(new_n1220), .C1(new_n812), .C2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n1160), .B2(new_n1013), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1154), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n986), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1236), .B1(new_n1238), .B2(new_n1155), .ZN(G381));
  NAND3_X1  g1039(.A1(new_n1014), .A2(new_n1037), .A3(new_n1099), .ZN(new_n1240));
  OR2_X1    g1040(.A1(G381), .A2(G384), .ZN(new_n1241));
  NOR4_X1   g1041(.A1(new_n1240), .A2(G396), .A3(G393), .A4(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT122), .B1(new_n1214), .B2(new_n1202), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1206), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1013), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1196), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1156), .A2(new_n1161), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1211), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n695), .B1(new_n1209), .B2(new_n1215), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1246), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1164), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1242), .A2(new_n1253), .ZN(G407));
  OAI21_X1  g1054(.A(new_n1253), .B1(new_n1242), .B2(new_n668), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(G213), .ZN(G409));
  INV_X1    g1056(.A(G213), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1257), .A2(G343), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1207), .A2(new_n986), .A3(new_n1209), .ZN(new_n1260));
  OAI21_X1  g1060(.A(KEYINPUT123), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT123), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1214), .A2(new_n1262), .A3(new_n1202), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1261), .A2(new_n1013), .A3(new_n1263), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1164), .A2(new_n1260), .A3(new_n1196), .A4(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1259), .B(new_n1265), .C1(new_n1251), .C2(new_n1164), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT125), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT124), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT60), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1162), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1237), .A2(KEYINPUT124), .A3(new_n1270), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n694), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1236), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(G384), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1237), .A2(KEYINPUT124), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(KEYINPUT60), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1278), .A2(new_n694), .A3(new_n1162), .A4(new_n1272), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G384), .B1(new_n1279), .B2(new_n1236), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1267), .B1(new_n1276), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1279), .A2(G384), .A3(new_n1236), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1282), .A2(KEYINPUT125), .A3(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1281), .A2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(KEYINPUT62), .B1(new_n1266), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1287), .A2(G2897), .A3(new_n1258), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1258), .A2(G2897), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1281), .A2(new_n1284), .A3(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1266), .A2(new_n1288), .A3(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1258), .B1(G375), .B2(G378), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT62), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1282), .A2(KEYINPUT125), .A3(new_n1283), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT125), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1292), .A2(new_n1293), .A3(new_n1265), .A4(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT61), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1286), .A2(new_n1291), .A3(new_n1297), .A4(new_n1298), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(G393), .B(G396), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1014), .A2(new_n1037), .A3(new_n1099), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1099), .B1(new_n1014), .B2(new_n1037), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1301), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(G387), .A2(G390), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1305), .A2(new_n1240), .A3(new_n1300), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1299), .A2(new_n1307), .ZN(new_n1308));
  AND2_X1   g1108(.A1(new_n1290), .A2(new_n1288), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT61), .B1(new_n1309), .B2(new_n1266), .ZN(new_n1310));
  AND2_X1   g1110(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1311));
  XOR2_X1   g1111(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1312));
  OAI21_X1  g1112(.A(new_n1312), .B1(new_n1266), .B2(new_n1285), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1292), .A2(KEYINPUT63), .A3(new_n1265), .A4(new_n1296), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1310), .A2(new_n1311), .A3(new_n1313), .A4(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1308), .A2(new_n1315), .ZN(G405));
  NAND2_X1  g1116(.A1(G375), .A2(G378), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1252), .A2(new_n1317), .A3(new_n1296), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(KEYINPUT127), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1252), .A2(new_n1317), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1287), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT127), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1252), .A2(new_n1317), .A3(new_n1296), .A4(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1319), .A2(new_n1321), .A3(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1307), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1311), .A2(new_n1319), .A3(new_n1321), .A4(new_n1323), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(G402));
endmodule


