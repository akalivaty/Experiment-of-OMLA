//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n811, new_n812, new_n814,
    new_n815, new_n816, new_n818, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942;
  NAND2_X1  g000(.A1(KEYINPUT76), .A2(KEYINPUT36), .ZN(new_n202));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT66), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT26), .ZN(new_n207));
  NOR3_X1   g006(.A1(KEYINPUT71), .A2(G169gat), .A3(G176gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n208), .A2(new_n207), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n203), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT68), .B(G190gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT27), .B(G183gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(G183gat), .B2(G190gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT24), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n203), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n203), .A2(KEYINPUT64), .A3(new_n221), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n220), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n206), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n226), .A2(new_n227), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT25), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT69), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237));
  INV_X1    g036(.A(G183gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n212), .A2(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n239), .A2(new_n219), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n222), .B(KEYINPUT67), .ZN(new_n241));
  AOI211_X1 g040(.A(new_n237), .B(new_n232), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  NOR3_X1   g041(.A1(new_n235), .A2(new_n236), .A3(new_n242), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n231), .A2(new_n206), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(new_n227), .B2(new_n226), .ZN(new_n245));
  INV_X1    g044(.A(new_n234), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n237), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n240), .A2(new_n241), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n248), .A2(KEYINPUT25), .A3(new_n244), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT69), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n218), .B1(new_n243), .B2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G113gat), .B(G120gat), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT1), .B1(new_n252), .B2(KEYINPUT73), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n253), .B1(KEYINPUT73), .B2(new_n252), .ZN(new_n254));
  NOR2_X1   g053(.A1(G127gat), .A2(G134gat), .ZN(new_n255));
  XOR2_X1   g054(.A(KEYINPUT72), .B(G127gat), .Z(new_n256));
  AOI21_X1  g055(.A(new_n255), .B1(new_n256), .B2(G134gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n259));
  AND2_X1   g058(.A1(G127gat), .A2(G134gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n259), .B1(new_n260), .B2(new_n255), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n261), .B1(KEYINPUT74), .B2(new_n252), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n262), .B1(KEYINPUT74), .B2(new_n252), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n251), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n236), .B1(new_n235), .B2(new_n242), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n247), .A2(KEYINPUT69), .A3(new_n249), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n217), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n264), .ZN(new_n270));
  INV_X1    g069(.A(G227gat), .ZN(new_n271));
  INV_X1    g070(.A(G233gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n266), .A2(new_n270), .A3(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(G71gat), .B(G99gat), .Z(new_n275));
  XNOR2_X1  g074(.A(G15gat), .B(G43gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT33), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n274), .A2(KEYINPUT32), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT75), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT75), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n274), .A2(new_n281), .A3(KEYINPUT32), .A4(new_n278), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT34), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n266), .A2(new_n270), .ZN(new_n285));
  INV_X1    g084(.A(new_n273), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AOI211_X1 g086(.A(KEYINPUT34), .B(new_n273), .C1(new_n266), .C2(new_n270), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT32), .ZN(new_n290));
  INV_X1    g089(.A(new_n274), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n290), .B(new_n277), .C1(new_n291), .C2(KEYINPUT33), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n283), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n289), .B1(new_n283), .B2(new_n292), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n202), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n283), .A2(new_n292), .ZN(new_n296));
  INV_X1    g095(.A(new_n289), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n283), .A2(new_n289), .A3(new_n292), .ZN(new_n299));
  XOR2_X1   g098(.A(KEYINPUT76), .B(KEYINPUT36), .Z(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n298), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n295), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G8gat), .B(G36gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(G64gat), .B(G92gat), .ZN(new_n305));
  XOR2_X1   g104(.A(new_n304), .B(new_n305), .Z(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  XOR2_X1   g106(.A(G197gat), .B(G204gat), .Z(new_n308));
  AOI21_X1  g107(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G211gat), .B(G218gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n312), .B(KEYINPUT78), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT77), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n311), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n315), .B1(new_n314), .B2(new_n310), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G226gat), .A2(G233gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n269), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n218), .B1(new_n235), .B2(new_n242), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n322), .A2(new_n323), .A3(new_n319), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n318), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  OAI211_X1 g124(.A(KEYINPUT79), .B(new_n319), .C1(new_n269), .C2(KEYINPUT29), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n320), .B1(new_n251), .B2(new_n323), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n322), .A2(new_n320), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT79), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n326), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n325), .B1(new_n331), .B2(new_n318), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT80), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n319), .B1(new_n269), .B2(KEYINPUT29), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n329), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n317), .B1(new_n336), .B2(new_n326), .ZN(new_n337));
  NOR3_X1   g136(.A1(new_n337), .A2(KEYINPUT80), .A3(new_n325), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n307), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G225gat), .A2(G233gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(KEYINPUT82), .B(G148gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G141gat), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n342), .A2(KEYINPUT83), .ZN(new_n343));
  INV_X1    g142(.A(G148gat), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n342), .B(KEYINPUT83), .C1(G141gat), .C2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G155gat), .ZN(new_n346));
  INV_X1    g145(.A(G162gat), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT2), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n348), .A2(KEYINPUT84), .ZN(new_n349));
  XOR2_X1   g148(.A(G155gat), .B(G162gat), .Z(new_n350));
  AOI21_X1  g149(.A(new_n350), .B1(KEYINPUT84), .B2(new_n348), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n343), .A2(new_n345), .A3(new_n349), .A4(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G141gat), .B(G148gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT81), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n348), .B1(new_n353), .B2(new_n354), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n350), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT3), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n352), .A2(new_n360), .A3(new_n357), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n264), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n340), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n358), .A2(new_n264), .ZN(new_n365));
  XOR2_X1   g164(.A(KEYINPUT85), .B(KEYINPUT4), .Z(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n369), .B1(new_n358), .B2(new_n264), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  OR3_X1    g170(.A1(new_n364), .A2(new_n371), .A3(KEYINPUT5), .ZN(new_n372));
  INV_X1    g171(.A(new_n340), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n359), .A2(new_n265), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n373), .B1(new_n374), .B2(new_n365), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n365), .A2(KEYINPUT4), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n376), .B1(new_n365), .B2(new_n367), .ZN(new_n377));
  OAI211_X1 g176(.A(KEYINPUT5), .B(new_n375), .C1(new_n377), .C2(new_n364), .ZN(new_n378));
  XOR2_X1   g177(.A(G57gat), .B(G85gat), .Z(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT87), .ZN(new_n380));
  XOR2_X1   g179(.A(G1gat), .B(G29gat), .Z(new_n381));
  XOR2_X1   g180(.A(new_n380), .B(new_n381), .Z(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n372), .A2(new_n378), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT6), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n384), .B1(new_n372), .B2(new_n378), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n332), .A2(new_n306), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT30), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n332), .A2(KEYINPUT30), .A3(new_n306), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n339), .A2(new_n389), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT88), .ZN(new_n395));
  NAND2_X1  g194(.A1(G228gat), .A2(G233gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT78), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n312), .B(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n310), .A2(new_n311), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n323), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n360), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n358), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n362), .A2(new_n323), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n318), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n397), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT29), .B1(new_n313), .B2(new_n316), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n358), .B1(new_n407), .B2(KEYINPUT3), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n408), .A2(new_n397), .A3(new_n405), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(G22gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(G22gat), .B1(new_n406), .B2(new_n409), .ZN(new_n413));
  XNOR2_X1  g212(.A(G78gat), .B(G106gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT31), .B(G50gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  AND4_X1   g215(.A1(new_n395), .A2(new_n412), .A3(new_n413), .A4(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n413), .A2(KEYINPUT88), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n418), .A2(new_n416), .B1(new_n412), .B2(new_n413), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n394), .A2(new_n420), .ZN(new_n421));
  OR2_X1    g220(.A1(new_n374), .A2(new_n365), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT39), .B1(new_n422), .B2(new_n373), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT89), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT89), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n425), .B(KEYINPUT39), .C1(new_n422), .C2(new_n373), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n368), .B(new_n370), .C1(new_n361), .C2(new_n363), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n373), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(KEYINPUT39), .ZN(new_n430));
  INV_X1    g229(.A(new_n384), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n429), .A2(new_n432), .A3(KEYINPUT40), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT40), .B1(new_n429), .B2(new_n432), .ZN(new_n434));
  NOR3_X1   g233(.A1(new_n433), .A2(new_n434), .A3(new_n388), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n392), .A2(new_n393), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n332), .A2(new_n333), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT80), .B1(new_n337), .B2(new_n325), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n306), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n435), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  OR2_X1    g239(.A1(new_n417), .A2(new_n419), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n372), .A2(new_n378), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n431), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n387), .B(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n390), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT37), .B1(new_n334), .B2(new_n338), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT38), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT37), .ZN(new_n449));
  AOI211_X1 g248(.A(new_n448), .B(new_n306), .C1(new_n332), .C2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n331), .A2(new_n317), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n321), .A2(new_n324), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n452), .B(KEYINPUT37), .C1(new_n317), .C2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n332), .A2(new_n449), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(new_n455), .A3(new_n307), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n448), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n446), .B1(new_n451), .B2(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n303), .B(new_n421), .C1(new_n442), .C2(new_n458), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n293), .A2(new_n420), .A3(new_n294), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n436), .A2(new_n445), .A3(new_n439), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT35), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n441), .A2(new_n298), .A3(new_n299), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT35), .B1(new_n464), .B2(new_n394), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(G113gat), .B(G141gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(G169gat), .B(G197gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  XOR2_X1   g269(.A(KEYINPUT90), .B(KEYINPUT11), .Z(new_n471));
  XNOR2_X1  g270(.A(new_n470), .B(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(KEYINPUT12), .ZN(new_n473));
  XOR2_X1   g272(.A(G15gat), .B(G22gat), .Z(new_n474));
  INV_X1    g273(.A(G1gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(G15gat), .B(G22gat), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT16), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n477), .B1(new_n478), .B2(G1gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n476), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  OR2_X1    g280(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  XOR2_X1   g282(.A(G43gat), .B(G50gat), .Z(new_n484));
  INV_X1    g283(.A(KEYINPUT15), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(G29gat), .ZN(new_n487));
  INV_X1    g286(.A(G36gat), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT14), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT14), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n490), .B1(G29gat), .B2(G36gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  OAI22_X1  g291(.A1(new_n492), .A2(KEYINPUT91), .B1(new_n487), .B2(new_n488), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n492), .A2(KEYINPUT91), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n486), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n492), .B1(G29gat), .B2(G36gat), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT92), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n497), .B1(new_n484), .B2(new_n485), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n484), .A2(new_n485), .ZN(new_n499));
  XNOR2_X1  g298(.A(G43gat), .B(G50gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(KEYINPUT92), .A3(KEYINPUT15), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n496), .A2(new_n498), .A3(new_n499), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n495), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n483), .B(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(G229gat), .A2(G233gat), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n505), .B(KEYINPUT13), .Z(new_n506));
  AND2_X1   g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n495), .A2(new_n502), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n483), .B1(KEYINPUT17), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT93), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT17), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n510), .B1(new_n503), .B2(new_n511), .ZN(new_n512));
  AOI211_X1 g311(.A(KEYINPUT93), .B(KEYINPUT17), .C1(new_n495), .C2(new_n502), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n483), .A2(new_n503), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n514), .A2(new_n505), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT18), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n507), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n514), .A2(KEYINPUT18), .A3(new_n505), .A4(new_n515), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n473), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n518), .A2(new_n519), .A3(new_n473), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g322(.A1(G232gat), .A2(G233gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n524), .A2(KEYINPUT41), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT99), .ZN(new_n526));
  XNOR2_X1  g325(.A(G134gat), .B(G162gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G85gat), .A2(G92gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT7), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n532), .A2(G85gat), .A3(G92gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(G99gat), .A2(G106gat), .ZN(new_n535));
  INV_X1    g334(.A(G85gat), .ZN(new_n536));
  INV_X1    g335(.A(G92gat), .ZN(new_n537));
  AOI22_X1  g336(.A1(KEYINPUT8), .A2(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G99gat), .B(G106gat), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n534), .A2(new_n538), .A3(new_n540), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n544), .B1(new_n508), .B2(KEYINPUT17), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(new_n513), .B2(new_n512), .ZN(new_n546));
  XNOR2_X1  g345(.A(G190gat), .B(G218gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT100), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n503), .A2(new_n544), .B1(KEYINPUT41), .B2(new_n524), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n546), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n549), .B1(new_n546), .B2(new_n550), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n529), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n553), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n555), .A2(new_n528), .A3(new_n551), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G71gat), .A2(G78gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT95), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT95), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n558), .A2(new_n562), .A3(new_n559), .ZN(new_n563));
  INV_X1    g362(.A(G57gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(G64gat), .ZN(new_n565));
  INV_X1    g364(.A(G64gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(G57gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n561), .A2(new_n563), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G71gat), .B(G78gat), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT96), .B1(new_n566), .B2(G57gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT96), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n574), .A2(new_n564), .A3(G64gat), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n573), .A2(new_n575), .A3(new_n567), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n576), .A2(new_n570), .A3(new_n563), .A4(new_n561), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(KEYINPUT97), .B(KEYINPUT21), .Z(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n582), .B(G127gat), .Z(new_n583));
  INV_X1    g382(.A(new_n578), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n483), .B1(KEYINPUT21), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n583), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G183gat), .B(G211gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT98), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(new_n346), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n588), .B(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n586), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n586), .A2(new_n592), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n557), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G230gat), .A2(G233gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT102), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n542), .A2(new_n543), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n578), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n572), .A2(new_n542), .A3(new_n577), .A4(new_n543), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(KEYINPUT101), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT101), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n578), .A2(new_n603), .A3(new_n599), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT10), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT10), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n598), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n602), .A2(new_n597), .A3(new_n604), .ZN(new_n609));
  XNOR2_X1  g408(.A(G120gat), .B(G148gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n610), .B(new_n611), .Z(new_n612));
  AND2_X1   g411(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n605), .A2(new_n607), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n597), .B(KEYINPUT104), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n609), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n612), .B(KEYINPUT103), .Z(new_n619));
  AOI21_X1  g418(.A(new_n615), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n595), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n467), .A2(new_n523), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n445), .B(KEYINPUT105), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(new_n475), .ZN(G1324gat));
  NOR2_X1   g425(.A1(new_n436), .A2(new_n439), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT16), .B(G8gat), .Z(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(G8gat), .B1(new_n623), .B2(new_n627), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(KEYINPUT42), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT106), .ZN(new_n634));
  AOI21_X1  g433(.A(KEYINPUT42), .B1(new_n628), .B2(new_n629), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT42), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n638), .B1(new_n630), .B2(new_n631), .ZN(new_n639));
  OAI21_X1  g438(.A(KEYINPUT106), .B1(new_n639), .B2(new_n635), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n640), .ZN(G1325gat));
  NAND2_X1  g440(.A1(new_n298), .A2(new_n299), .ZN(new_n642));
  OR3_X1    g441(.A1(new_n623), .A2(G15gat), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(G15gat), .B1(new_n623), .B2(new_n303), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(G1326gat));
  NOR2_X1   g444(.A1(new_n623), .A2(new_n441), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT43), .B(G22gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(G1327gat));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n447), .A2(new_n450), .B1(new_n456), .B2(new_n448), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n441), .B(new_n440), .C1(new_n650), .C2(new_n446), .ZN(new_n651));
  AOI22_X1  g450(.A1(new_n295), .A2(new_n302), .B1(new_n394), .B2(new_n420), .ZN(new_n652));
  AOI22_X1  g451(.A1(new_n651), .A2(new_n652), .B1(new_n463), .B2(new_n465), .ZN(new_n653));
  INV_X1    g452(.A(new_n557), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n467), .A2(KEYINPUT44), .A3(new_n557), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n593), .A2(new_n594), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n516), .A2(new_n517), .ZN(new_n659));
  INV_X1    g458(.A(new_n507), .ZN(new_n660));
  AND4_X1   g459(.A1(new_n519), .A2(new_n659), .A3(new_n660), .A4(new_n473), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(new_n520), .ZN(new_n662));
  INV_X1    g461(.A(new_n620), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n658), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n657), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(G29gat), .B1(new_n665), .B2(new_n624), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n653), .A2(new_n654), .ZN(new_n667));
  INV_X1    g466(.A(new_n624), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n667), .A2(new_n487), .A3(new_n668), .A4(new_n664), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT45), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n666), .A2(new_n670), .ZN(G1328gat));
  NAND2_X1  g470(.A1(new_n667), .A2(new_n664), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n672), .A2(G36gat), .A3(new_n627), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT46), .ZN(new_n674));
  OAI21_X1  g473(.A(G36gat), .B1(new_n665), .B2(new_n627), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(G1329gat));
  NOR2_X1   g475(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT108), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT47), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n642), .A2(G43gat), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n467), .A2(new_n557), .A3(new_n664), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT107), .ZN(new_n683));
  INV_X1    g482(.A(new_n303), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n655), .A2(new_n656), .A3(new_n684), .A4(new_n664), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(G43gat), .ZN(new_n686));
  AOI211_X1 g485(.A(new_n677), .B(new_n680), .C1(new_n683), .C2(new_n686), .ZN(new_n687));
  AND4_X1   g486(.A1(new_n678), .A2(new_n683), .A3(new_n686), .A4(new_n679), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(G1330gat));
  INV_X1    g488(.A(G50gat), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(new_n672), .B2(new_n441), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n441), .A2(new_n690), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n665), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT48), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT48), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n696), .B(new_n691), .C1(new_n665), .C2(new_n693), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(G1331gat));
  NAND3_X1  g497(.A1(new_n595), .A2(new_n662), .A3(new_n663), .ZN(new_n699));
  OR3_X1    g498(.A1(new_n653), .A2(KEYINPUT109), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT109), .B1(new_n653), .B2(new_n699), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(new_n624), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(new_n564), .ZN(G1332gat));
  NOR2_X1   g503(.A1(new_n702), .A2(new_n627), .ZN(new_n705));
  NOR2_X1   g504(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n706));
  AND2_X1   g505(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n708), .B1(new_n705), .B2(new_n706), .ZN(G1333gat));
  INV_X1    g508(.A(G71gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n642), .B(KEYINPUT110), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n710), .B1(new_n702), .B2(new_n711), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n700), .A2(G71gat), .A3(new_n684), .A4(new_n701), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(G1334gat));
  NOR2_X1   g518(.A1(new_n702), .A2(new_n441), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(G78gat), .Z(G1335gat));
  NOR3_X1   g520(.A1(new_n658), .A2(new_n523), .A3(new_n620), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n657), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G85gat), .B1(new_n723), .B2(new_n624), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n658), .A2(new_n523), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n467), .A2(new_n557), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT51), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n728), .A2(new_n536), .A3(new_n663), .A4(new_n668), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n724), .A2(new_n729), .ZN(G1336gat));
  NOR3_X1   g529(.A1(new_n627), .A2(G92gat), .A3(new_n620), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733));
  INV_X1    g532(.A(new_n627), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n655), .A2(new_n656), .A3(new_n734), .A4(new_n722), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G92gat), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n732), .A2(new_n733), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n726), .B(new_n738), .ZN(new_n739));
  AOI22_X1  g538(.A1(new_n739), .A2(new_n731), .B1(G92gat), .B2(new_n735), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n737), .B1(new_n733), .B2(new_n740), .ZN(G1337gat));
  OAI21_X1  g540(.A(G99gat), .B1(new_n723), .B2(new_n303), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n642), .A2(G99gat), .A3(new_n620), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(G1338gat));
  NOR3_X1   g544(.A1(new_n441), .A2(G106gat), .A3(new_n620), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT53), .B1(new_n728), .B2(new_n746), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n655), .A2(new_n656), .A3(new_n420), .A4(new_n722), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT113), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G106gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n747), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n726), .A2(new_n738), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n726), .A2(new_n738), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n746), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n748), .A2(G106gat), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT53), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n753), .A2(new_n759), .ZN(G1339gat));
  NOR2_X1   g559(.A1(new_n662), .A2(G113gat), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n505), .B1(new_n514), .B2(new_n515), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n504), .A2(new_n506), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n472), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n663), .A2(new_n522), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n601), .A2(KEYINPUT101), .ZN(new_n766));
  AOI22_X1  g565(.A1(new_n572), .A2(new_n577), .B1(new_n542), .B2(new_n543), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n604), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n606), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n607), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n770), .A2(new_n771), .A3(new_n617), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT114), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n770), .A2(new_n774), .A3(new_n771), .A4(new_n617), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n773), .A2(KEYINPUT54), .A3(new_n608), .A4(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777));
  INV_X1    g576(.A(new_n617), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n777), .B(new_n778), .C1(new_n605), .C2(new_n607), .ZN(new_n779));
  INV_X1    g578(.A(new_n612), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n779), .A2(KEYINPUT55), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n615), .B1(new_n776), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n779), .A2(new_n780), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT55), .B1(new_n776), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(KEYINPUT115), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n605), .A2(new_n607), .A3(new_n778), .ZN(new_n786));
  OAI211_X1 g585(.A(KEYINPUT54), .B(new_n608), .C1(new_n786), .C2(new_n774), .ZN(new_n787));
  INV_X1    g586(.A(new_n775), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n789), .A2(KEYINPUT115), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n782), .B1(new_n785), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n765), .B1(new_n792), .B2(new_n662), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n654), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n557), .A2(new_n522), .A3(new_n764), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n795), .B(new_n782), .C1(new_n791), .C2(new_n785), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n658), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n621), .A2(new_n523), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n668), .A2(new_n627), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n799), .A2(new_n464), .A3(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(KEYINPUT116), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n801), .A2(KEYINPUT116), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n761), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n801), .ZN(new_n805));
  OAI21_X1  g604(.A(G113gat), .B1(new_n805), .B2(new_n662), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(G1340gat));
  NOR2_X1   g606(.A1(new_n620), .A2(G120gat), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n802), .B2(new_n803), .ZN(new_n809));
  OAI21_X1  g608(.A(G120gat), .B1(new_n805), .B2(new_n620), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n811), .B(new_n812), .ZN(G1341gat));
  NAND2_X1  g612(.A1(new_n801), .A2(new_n658), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n256), .A2(new_n815), .ZN(new_n816));
  XOR2_X1   g615(.A(new_n814), .B(new_n816), .Z(G1342gat));
  NAND3_X1  g616(.A1(new_n668), .A2(new_n627), .A3(new_n557), .ZN(new_n818));
  NOR4_X1   g617(.A1(new_n799), .A2(G134gat), .A3(new_n464), .A4(new_n818), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(KEYINPUT56), .ZN(new_n820));
  OAI21_X1  g619(.A(G134gat), .B1(new_n805), .B2(new_n654), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(G1343gat));
  NOR2_X1   g621(.A1(new_n799), .A2(new_n441), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n800), .A2(new_n684), .ZN(new_n826));
  INV_X1    g625(.A(new_n658), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n781), .B1(new_n787), .B2(new_n788), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n614), .ZN(new_n829));
  OAI21_X1  g628(.A(KEYINPUT119), .B1(new_n829), .B2(new_n784), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n789), .A2(new_n790), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(new_n782), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n830), .A2(new_n523), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n557), .B1(new_n834), .B2(new_n765), .ZN(new_n835));
  INV_X1    g634(.A(new_n796), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n827), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n622), .A2(new_n662), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n441), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n825), .B(new_n826), .C1(new_n824), .C2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(G141gat), .B1(new_n840), .B2(new_n662), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n823), .A2(new_n826), .ZN(new_n842));
  INV_X1    g641(.A(G141gat), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n843), .A3(new_n523), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT58), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n841), .A2(new_n847), .A3(new_n844), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(G1344gat));
  NOR2_X1   g648(.A1(new_n341), .A2(KEYINPUT59), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n850), .B1(new_n840), .B2(new_n620), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n852));
  INV_X1    g651(.A(new_n765), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n829), .A2(new_n784), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n662), .B1(new_n854), .B2(new_n832), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n853), .B1(new_n855), .B2(new_n830), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n796), .B1(new_n856), .B2(new_n557), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n798), .B1(new_n857), .B2(new_n827), .ZN(new_n858));
  OAI211_X1 g657(.A(KEYINPUT120), .B(new_n824), .C1(new_n858), .C2(new_n441), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n860), .B1(new_n839), .B2(KEYINPUT57), .ZN(new_n861));
  OAI211_X1 g660(.A(KEYINPUT57), .B(new_n420), .C1(new_n797), .C2(new_n798), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n859), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n800), .A2(new_n684), .A3(new_n620), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(G148gat), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n852), .B1(new_n866), .B2(KEYINPUT59), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n344), .B1(new_n863), .B2(new_n864), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n868), .A2(KEYINPUT121), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n851), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n823), .A2(new_n341), .A3(new_n864), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(G1345gat));
  NOR3_X1   g672(.A1(new_n840), .A2(new_n346), .A3(new_n827), .ZN(new_n874));
  AOI21_X1  g673(.A(G155gat), .B1(new_n842), .B2(new_n658), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n874), .A2(new_n875), .ZN(G1346gat));
  NOR3_X1   g675(.A1(new_n818), .A2(new_n684), .A3(G162gat), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n823), .A2(new_n877), .ZN(new_n878));
  XOR2_X1   g677(.A(new_n878), .B(KEYINPUT122), .Z(new_n879));
  OAI21_X1  g678(.A(G162gat), .B1(new_n840), .B2(new_n654), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1347gat));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n882));
  INV_X1    g681(.A(new_n711), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n624), .A2(new_n734), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT123), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n624), .A2(new_n734), .A3(KEYINPUT123), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n883), .A2(new_n886), .A3(new_n441), .A4(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n882), .B1(new_n888), .B2(new_n799), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n886), .A2(new_n887), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n711), .A2(new_n420), .ZN(new_n892));
  INV_X1    g691(.A(new_n799), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n891), .A2(new_n892), .A3(new_n893), .A4(KEYINPUT124), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G169gat), .B1(new_n895), .B2(new_n662), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT125), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n799), .A2(new_n464), .A3(new_n884), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  OR3_X1    g698(.A1(new_n899), .A2(G169gat), .A3(new_n662), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n896), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n897), .B1(new_n896), .B2(new_n900), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(new_n902), .ZN(G1348gat));
  OAI21_X1  g702(.A(G176gat), .B1(new_n895), .B2(new_n620), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n620), .A2(G176gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n899), .B2(new_n905), .ZN(G1349gat));
  OAI21_X1  g705(.A(G183gat), .B1(new_n895), .B2(new_n827), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n898), .A2(new_n213), .A3(new_n658), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT60), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n907), .A2(new_n911), .A3(new_n908), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(G1350gat));
  NAND3_X1  g712(.A1(new_n898), .A2(new_n212), .A3(new_n557), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n889), .A2(new_n894), .A3(new_n557), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT61), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n915), .A2(new_n916), .A3(G190gat), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n915), .B2(G190gat), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n914), .B1(new_n917), .B2(new_n918), .ZN(G1351gat));
  NOR2_X1   g718(.A1(new_n890), .A2(new_n684), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n863), .A2(new_n523), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G197gat), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n684), .A2(new_n884), .A3(new_n441), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n893), .A2(new_n923), .ZN(new_n924));
  OR3_X1    g723(.A1(new_n924), .A2(G197gat), .A3(new_n662), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT126), .ZN(G1352gat));
  NOR3_X1   g726(.A1(new_n924), .A2(G204gat), .A3(new_n620), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT62), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n863), .A2(new_n920), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n663), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(G204gat), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n929), .A2(new_n932), .ZN(G1353gat));
  OR3_X1    g732(.A1(new_n924), .A2(G211gat), .A3(new_n827), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n930), .A2(new_n658), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n935), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT63), .B1(new_n935), .B2(G211gat), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(G1354gat));
  NAND2_X1  g737(.A1(new_n557), .A2(G218gat), .ZN(new_n939));
  XOR2_X1   g738(.A(new_n939), .B(KEYINPUT127), .Z(new_n940));
  INV_X1    g739(.A(G218gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n893), .A2(new_n923), .A3(new_n557), .ZN(new_n942));
  AOI22_X1  g741(.A1(new_n930), .A2(new_n940), .B1(new_n941), .B2(new_n942), .ZN(G1355gat));
endmodule


