

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759;

  OR2_X1 U374 ( .A1(n669), .A2(n670), .ZN(n666) );
  NOR2_X1 U375 ( .A1(n667), .A2(n666), .ZN(n630) );
  XNOR2_X2 U376 ( .A(n550), .B(n551), .ZN(n653) );
  XNOR2_X2 U377 ( .A(n610), .B(n611), .ZN(n614) );
  AND2_X2 U378 ( .A1(n431), .A2(n361), .ZN(n434) );
  XNOR2_X2 U379 ( .A(n537), .B(n536), .ZN(n742) );
  XNOR2_X1 U380 ( .A(n624), .B(n623), .ZN(n754) );
  XNOR2_X1 U381 ( .A(n556), .B(KEYINPUT42), .ZN(n756) );
  XNOR2_X1 U382 ( .A(n485), .B(n484), .ZN(n580) );
  XNOR2_X1 U383 ( .A(n493), .B(n355), .ZN(n553) );
  NOR2_X1 U384 ( .A1(n695), .A2(G902), .ZN(n493) );
  XNOR2_X1 U385 ( .A(n513), .B(n512), .ZN(n669) );
  XNOR2_X1 U386 ( .A(n526), .B(n525), .ZN(n576) );
  XNOR2_X1 U387 ( .A(n489), .B(n456), .ZN(n379) );
  XNOR2_X1 U388 ( .A(n504), .B(n392), .ZN(n391) );
  XNOR2_X1 U389 ( .A(n368), .B(G128), .ZN(n489) );
  XNOR2_X1 U390 ( .A(n370), .B(KEYINPUT4), .ZN(n491) );
  XNOR2_X1 U391 ( .A(n482), .B(n398), .ZN(n501) );
  INV_X1 U392 ( .A(KEYINPUT65), .ZN(n370) );
  XOR2_X1 U393 ( .A(G146), .B(G125), .Z(n504) );
  NAND2_X1 U394 ( .A1(n382), .A2(n380), .ZN(n593) );
  INV_X1 U395 ( .A(G143), .ZN(n368) );
  INV_X1 U396 ( .A(n535), .ZN(n536) );
  XNOR2_X1 U397 ( .A(n568), .B(KEYINPUT46), .ZN(n437) );
  AND2_X1 U398 ( .A1(n756), .A2(n757), .ZN(n568) );
  INV_X1 U399 ( .A(n719), .ZN(n389) );
  NOR2_X1 U400 ( .A1(G953), .A2(G237), .ZN(n518) );
  INV_X1 U401 ( .A(n576), .ZN(n405) );
  OR2_X1 U402 ( .A1(G902), .A2(G237), .ZN(n544) );
  XNOR2_X1 U403 ( .A(n463), .B(n391), .ZN(n464) );
  NOR2_X1 U404 ( .A1(G902), .A2(n726), .ZN(n513) );
  INV_X1 U405 ( .A(KEYINPUT25), .ZN(n510) );
  XNOR2_X1 U406 ( .A(n491), .B(n490), .ZN(n369) );
  INV_X1 U407 ( .A(G137), .ZN(n490) );
  XOR2_X1 U408 ( .A(G122), .B(G116), .Z(n527) );
  XNOR2_X1 U409 ( .A(n478), .B(n477), .ZN(n486) );
  XNOR2_X1 U410 ( .A(G119), .B(G113), .ZN(n477) );
  XNOR2_X1 U411 ( .A(n448), .B(n447), .ZN(n531) );
  INV_X1 U412 ( .A(KEYINPUT8), .ZN(n447) );
  NAND2_X1 U413 ( .A1(n356), .A2(G234), .ZN(n448) );
  XNOR2_X1 U414 ( .A(n504), .B(n427), .ZN(n743) );
  XNOR2_X1 U415 ( .A(KEYINPUT10), .B(KEYINPUT69), .ZN(n427) );
  XNOR2_X1 U416 ( .A(n471), .B(n470), .ZN(n541) );
  XNOR2_X1 U417 ( .A(G107), .B(G104), .ZN(n470) );
  AND2_X1 U418 ( .A1(n376), .A2(n360), .ZN(n374) );
  NAND2_X1 U419 ( .A1(n631), .A2(KEYINPUT34), .ZN(n375) );
  NOR2_X1 U420 ( .A1(G902), .A2(n722), .ZN(n543) );
  AND2_X1 U421 ( .A1(n371), .A2(n424), .ZN(n422) );
  INV_X1 U422 ( .A(KEYINPUT84), .ZN(n436) );
  NAND2_X1 U423 ( .A1(n501), .A2(G234), .ZN(n502) );
  XOR2_X1 U424 ( .A(KEYINPUT95), .B(KEYINPUT97), .Z(n516) );
  INV_X1 U425 ( .A(n501), .ZN(n646) );
  NAND2_X1 U426 ( .A1(n383), .A2(n389), .ZN(n382) );
  NAND2_X1 U427 ( .A1(n385), .A2(n387), .ZN(n383) );
  NAND2_X1 U428 ( .A1(n388), .A2(n592), .ZN(n387) );
  NAND2_X1 U429 ( .A1(n384), .A2(n381), .ZN(n380) );
  AND2_X1 U430 ( .A1(n354), .A2(n437), .ZN(n384) );
  XNOR2_X1 U431 ( .A(n506), .B(n445), .ZN(n444) );
  XNOR2_X1 U432 ( .A(KEYINPUT23), .B(G119), .ZN(n506) );
  XNOR2_X1 U433 ( .A(G110), .B(G137), .ZN(n445) );
  XNOR2_X1 U434 ( .A(n428), .B(n426), .ZN(n524) );
  NAND2_X1 U435 ( .A1(G214), .A2(n544), .ZN(n656) );
  XNOR2_X1 U436 ( .A(n458), .B(n457), .ZN(n594) );
  XNOR2_X1 U437 ( .A(KEYINPUT39), .B(KEYINPUT85), .ZN(n457) );
  AND2_X1 U438 ( .A1(n569), .A2(n657), .ZN(n458) );
  XNOR2_X1 U439 ( .A(n416), .B(n415), .ZN(n588) );
  INV_X1 U440 ( .A(KEYINPUT106), .ZN(n415) );
  AND2_X1 U441 ( .A1(n534), .A2(n619), .ZN(n416) );
  XNOR2_X1 U442 ( .A(n630), .B(n372), .ZN(n620) );
  INV_X1 U443 ( .A(KEYINPUT102), .ZN(n372) );
  XNOR2_X1 U444 ( .A(n407), .B(n417), .ZN(n619) );
  XNOR2_X1 U445 ( .A(KEYINPUT99), .B(KEYINPUT6), .ZN(n417) );
  XNOR2_X1 U446 ( .A(n483), .B(KEYINPUT89), .ZN(n484) );
  XNOR2_X1 U447 ( .A(n414), .B(n412), .ZN(n488) );
  NAND2_X1 U448 ( .A1(n727), .A2(G472), .ZN(n442) );
  XNOR2_X1 U449 ( .A(n530), .B(n406), .ZN(n725) );
  XNOR2_X1 U450 ( .A(G107), .B(KEYINPUT9), .ZN(n528) );
  NAND2_X1 U451 ( .A1(n727), .A2(G478), .ZN(n455) );
  NAND2_X1 U452 ( .A1(n727), .A2(G475), .ZN(n411) );
  XOR2_X1 U453 ( .A(G146), .B(KEYINPUT76), .Z(n539) );
  XNOR2_X1 U454 ( .A(n396), .B(n365), .ZN(n397) );
  NAND2_X1 U455 ( .A1(n727), .A2(G210), .ZN(n396) );
  NOR2_X1 U456 ( .A1(n710), .A2(n595), .ZN(n660) );
  NAND2_X1 U457 ( .A1(n667), .A2(n436), .ZN(n435) );
  INV_X1 U458 ( .A(KEYINPUT17), .ZN(n392) );
  XOR2_X1 U459 ( .A(KEYINPUT77), .B(KEYINPUT18), .Z(n462) );
  INV_X1 U460 ( .A(G131), .ZN(n395) );
  INV_X1 U461 ( .A(n743), .ZN(n426) );
  XNOR2_X1 U462 ( .A(n517), .B(n519), .ZN(n428) );
  XNOR2_X1 U463 ( .A(G122), .B(G104), .ZN(n515) );
  XOR2_X1 U464 ( .A(KEYINPUT12), .B(KEYINPUT96), .Z(n521) );
  XOR2_X1 U465 ( .A(G131), .B(G140), .Z(n535) );
  XNOR2_X1 U466 ( .A(n580), .B(n548), .ZN(n657) );
  NAND2_X1 U467 ( .A1(n634), .A2(n378), .ZN(n377) );
  XNOR2_X1 U468 ( .A(n563), .B(n402), .ZN(n401) );
  INV_X1 U469 ( .A(KEYINPUT30), .ZN(n402) );
  NAND2_X1 U470 ( .A1(n407), .A2(n656), .ZN(n563) );
  INV_X1 U471 ( .A(KEYINPUT87), .ZN(n398) );
  XNOR2_X1 U472 ( .A(G902), .B(KEYINPUT15), .ZN(n482) );
  XNOR2_X1 U473 ( .A(n590), .B(KEYINPUT19), .ZN(n605) );
  XNOR2_X1 U474 ( .A(n399), .B(n394), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n400), .B(KEYINPUT92), .ZN(n399) );
  XNOR2_X1 U476 ( .A(n395), .B(G146), .ZN(n394) );
  INV_X1 U477 ( .A(KEYINPUT5), .ZN(n400) );
  XNOR2_X1 U478 ( .A(n413), .B(KEYINPUT91), .ZN(n412) );
  XNOR2_X1 U479 ( .A(G116), .B(G101), .ZN(n413) );
  INV_X1 U480 ( .A(G134), .ZN(n456) );
  AND2_X1 U481 ( .A1(n646), .A2(n645), .ZN(n424) );
  NAND2_X1 U482 ( .A1(n580), .A2(n656), .ZN(n590) );
  XNOR2_X1 U483 ( .A(n533), .B(G478), .ZN(n575) );
  XOR2_X1 U484 ( .A(KEYINPUT16), .B(KEYINPUT74), .Z(n472) );
  XNOR2_X1 U485 ( .A(n446), .B(n443), .ZN(n508) );
  XNOR2_X1 U486 ( .A(n507), .B(n444), .ZN(n443) );
  NOR2_X1 U487 ( .A1(n580), .A2(n547), .ZN(n719) );
  XNOR2_X1 U488 ( .A(n567), .B(n566), .ZN(n757) );
  NAND2_X1 U489 ( .A1(n374), .A2(n373), .ZN(n624) );
  NAND2_X1 U490 ( .A1(n614), .A2(n667), .ZN(n629) );
  NAND2_X1 U491 ( .A1(n441), .A2(n452), .ZN(n440) );
  XNOR2_X1 U492 ( .A(n442), .B(n364), .ZN(n441) );
  NAND2_X1 U493 ( .A1(n453), .A2(n452), .ZN(n451) );
  XNOR2_X1 U494 ( .A(n455), .B(n454), .ZN(n453) );
  INV_X1 U495 ( .A(KEYINPUT60), .ZN(n408) );
  NAND2_X1 U496 ( .A1(n410), .A2(n452), .ZN(n409) );
  XNOR2_X1 U497 ( .A(n411), .B(n366), .ZN(n410) );
  XNOR2_X1 U498 ( .A(n720), .B(n404), .ZN(n723) );
  XNOR2_X1 U499 ( .A(n722), .B(n721), .ZN(n404) );
  NAND2_X1 U500 ( .A1(n397), .A2(n452), .ZN(n393) );
  INV_X1 U501 ( .A(n667), .ZN(n438) );
  AND2_X1 U502 ( .A1(n433), .A2(n432), .ZN(n353) );
  AND2_X1 U503 ( .A1(n353), .A2(KEYINPUT48), .ZN(n354) );
  XOR2_X1 U504 ( .A(KEYINPUT71), .B(G472), .Z(n355) );
  XOR2_X1 U505 ( .A(G953), .B(KEYINPUT64), .Z(n356) );
  XNOR2_X1 U506 ( .A(n379), .B(n369), .ZN(n537) );
  AND2_X1 U507 ( .A1(n575), .A2(n405), .ZN(n357) );
  OR2_X1 U508 ( .A1(n562), .A2(n561), .ZN(n358) );
  AND2_X1 U509 ( .A1(n745), .A2(n423), .ZN(n652) );
  AND2_X1 U510 ( .A1(n667), .A2(n553), .ZN(n359) );
  AND2_X1 U511 ( .A1(n375), .A2(n622), .ZN(n360) );
  AND2_X1 U512 ( .A1(n587), .A2(n435), .ZN(n361) );
  AND2_X1 U513 ( .A1(n438), .A2(KEYINPUT84), .ZN(n362) );
  XOR2_X1 U514 ( .A(KEYINPUT36), .B(KEYINPUT113), .Z(n363) );
  XOR2_X1 U515 ( .A(n695), .B(KEYINPUT62), .Z(n364) );
  XOR2_X1 U516 ( .A(n650), .B(n649), .Z(n365) );
  XNOR2_X1 U517 ( .A(n724), .B(KEYINPUT59), .ZN(n366) );
  XNOR2_X1 U518 ( .A(n742), .B(n542), .ZN(n722) );
  INV_X1 U519 ( .A(KEYINPUT48), .ZN(n592) );
  XOR2_X1 U520 ( .A(n651), .B(KEYINPUT83), .Z(n367) );
  INV_X1 U521 ( .A(n730), .ZN(n452) );
  NAND2_X1 U522 ( .A1(n745), .A2(n371), .ZN(n655) );
  NAND2_X1 U523 ( .A1(n371), .A2(n736), .ZN(n737) );
  AND2_X1 U524 ( .A1(n371), .A2(n645), .ZN(n423) );
  XNOR2_X2 U525 ( .A(n642), .B(KEYINPUT45), .ZN(n371) );
  XNOR2_X2 U526 ( .A(n560), .B(KEYINPUT1), .ZN(n667) );
  XNOR2_X2 U527 ( .A(n543), .B(G469), .ZN(n560) );
  OR2_X1 U528 ( .A1(n665), .A2(n377), .ZN(n376) );
  XNOR2_X1 U529 ( .A(n621), .B(KEYINPUT33), .ZN(n665) );
  NAND2_X1 U530 ( .A1(n665), .A2(KEYINPUT34), .ZN(n373) );
  INV_X1 U531 ( .A(KEYINPUT34), .ZN(n378) );
  XNOR2_X1 U532 ( .A(n532), .B(n379), .ZN(n406) );
  AND2_X1 U533 ( .A1(n434), .A2(n389), .ZN(n381) );
  NAND2_X1 U534 ( .A1(n386), .A2(n592), .ZN(n385) );
  NAND2_X1 U535 ( .A1(n437), .A2(n353), .ZN(n386) );
  INV_X1 U536 ( .A(n434), .ZN(n388) );
  XNOR2_X1 U537 ( .A(n574), .B(KEYINPUT108), .ZN(n758) );
  NAND2_X1 U538 ( .A1(n390), .A2(n401), .ZN(n564) );
  NAND2_X1 U539 ( .A1(n429), .A2(n430), .ZN(n390) );
  XNOR2_X1 U540 ( .A(n409), .B(n408), .ZN(G60) );
  NOR2_X1 U541 ( .A1(n702), .A2(n755), .ZN(n420) );
  XNOR2_X1 U542 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U543 ( .A(n393), .B(n367), .ZN(G51) );
  INV_X1 U544 ( .A(n669), .ZN(n450) );
  NAND2_X2 U545 ( .A1(n647), .A2(n421), .ZN(n727) );
  NOR2_X1 U546 ( .A1(n358), .A2(n560), .ZN(n429) );
  NAND2_X1 U547 ( .A1(n403), .A2(n418), .ZN(n641) );
  NAND2_X1 U548 ( .A1(n625), .A2(n626), .ZN(n403) );
  NAND2_X1 U549 ( .A1(n509), .A2(G221), .ZN(n503) );
  XNOR2_X1 U550 ( .A(n502), .B(KEYINPUT20), .ZN(n509) );
  NOR2_X2 U551 ( .A1(n565), .A2(n564), .ZN(n569) );
  INV_X1 U552 ( .A(n575), .ZN(n571) );
  NAND2_X1 U553 ( .A1(n558), .A2(n450), .ZN(n449) );
  INV_X1 U554 ( .A(n553), .ZN(n407) );
  NAND2_X1 U555 ( .A1(n419), .A2(n754), .ZN(n418) );
  XNOR2_X1 U556 ( .A(n420), .B(n618), .ZN(n419) );
  NAND2_X1 U557 ( .A1(n422), .A2(n745), .ZN(n421) );
  AND2_X2 U558 ( .A1(n597), .A2(n596), .ZN(n745) );
  NAND2_X1 U559 ( .A1(n614), .A2(n359), .ZN(n425) );
  XNOR2_X1 U560 ( .A(n425), .B(KEYINPUT66), .ZN(n612) );
  NAND2_X1 U561 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U562 ( .A1(n666), .A2(n560), .ZN(n635) );
  INV_X1 U563 ( .A(n666), .ZN(n430) );
  XNOR2_X1 U564 ( .A(n584), .B(KEYINPUT79), .ZN(n431) );
  AND2_X1 U565 ( .A1(n439), .A2(n438), .ZN(n715) );
  OR2_X1 U566 ( .A1(n439), .A2(KEYINPUT84), .ZN(n432) );
  NAND2_X1 U567 ( .A1(n439), .A2(n362), .ZN(n433) );
  XNOR2_X1 U568 ( .A(n591), .B(n363), .ZN(n439) );
  XNOR2_X1 U569 ( .A(n440), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U570 ( .A1(n531), .A2(G221), .ZN(n446) );
  NOR2_X1 U571 ( .A1(n560), .A2(n449), .ZN(n559) );
  XNOR2_X1 U572 ( .A(n451), .B(KEYINPUT123), .ZN(G63) );
  INV_X1 U573 ( .A(n725), .ZN(n454) );
  NAND2_X1 U574 ( .A1(n594), .A2(n710), .ZN(n566) );
  OR2_X1 U575 ( .A1(n661), .A2(n659), .ZN(n550) );
  XNOR2_X1 U576 ( .A(n486), .B(n527), .ZN(n479) );
  XOR2_X1 U577 ( .A(n521), .B(n520), .Z(n459) );
  AND2_X1 U578 ( .A1(n518), .A2(G210), .ZN(n460) );
  INV_X1 U579 ( .A(KEYINPUT78), .ZN(n578) );
  XNOR2_X1 U580 ( .A(n579), .B(n578), .ZN(n583) );
  XNOR2_X1 U581 ( .A(n486), .B(n460), .ZN(n487) );
  INV_X1 U582 ( .A(KEYINPUT38), .ZN(n548) );
  XNOR2_X1 U583 ( .A(n488), .B(n487), .ZN(n492) );
  XNOR2_X1 U584 ( .A(n522), .B(n459), .ZN(n523) );
  INV_X1 U585 ( .A(n718), .ZN(n596) );
  XNOR2_X1 U586 ( .A(n524), .B(n523), .ZN(n724) );
  XNOR2_X1 U587 ( .A(n480), .B(n479), .ZN(n731) );
  XNOR2_X1 U588 ( .A(KEYINPUT35), .B(KEYINPUT81), .ZN(n623) );
  NOR2_X1 U589 ( .A1(n746), .A2(G952), .ZN(n730) );
  XNOR2_X1 U590 ( .A(n694), .B(n693), .ZN(G75) );
  XOR2_X2 U591 ( .A(G953), .B(KEYINPUT64), .Z(n746) );
  NAND2_X1 U592 ( .A1(G224), .A2(n746), .ZN(n461) );
  XNOR2_X1 U593 ( .A(n462), .B(n461), .ZN(n465) );
  XNOR2_X1 U594 ( .A(n489), .B(n491), .ZN(n463) );
  XNOR2_X1 U595 ( .A(n465), .B(n464), .ZN(n481) );
  INV_X1 U596 ( .A(G110), .ZN(n466) );
  NAND2_X1 U597 ( .A1(n466), .A2(G101), .ZN(n469) );
  INV_X1 U598 ( .A(G101), .ZN(n467) );
  NAND2_X1 U599 ( .A1(n467), .A2(G110), .ZN(n468) );
  NAND2_X1 U600 ( .A1(n469), .A2(n468), .ZN(n471) );
  XNOR2_X1 U601 ( .A(n541), .B(n472), .ZN(n480) );
  INV_X1 U602 ( .A(KEYINPUT3), .ZN(n473) );
  NAND2_X1 U603 ( .A1(KEYINPUT88), .A2(n473), .ZN(n476) );
  INV_X1 U604 ( .A(KEYINPUT88), .ZN(n474) );
  NAND2_X1 U605 ( .A1(n474), .A2(KEYINPUT3), .ZN(n475) );
  NAND2_X1 U606 ( .A1(n476), .A2(n475), .ZN(n478) );
  XNOR2_X1 U607 ( .A(n481), .B(n731), .ZN(n648) );
  NAND2_X1 U608 ( .A1(n648), .A2(n501), .ZN(n485) );
  NAND2_X1 U609 ( .A1(G210), .A2(n544), .ZN(n483) );
  XNOR2_X1 U610 ( .A(n492), .B(n537), .ZN(n695) );
  NAND2_X1 U611 ( .A1(G237), .A2(G234), .ZN(n494) );
  XNOR2_X1 U612 ( .A(n494), .B(KEYINPUT14), .ZN(n496) );
  NAND2_X1 U613 ( .A1(n496), .A2(G952), .ZN(n495) );
  XNOR2_X1 U614 ( .A(n495), .B(KEYINPUT90), .ZN(n686) );
  NOR2_X1 U615 ( .A1(G953), .A2(n686), .ZN(n602) );
  NAND2_X1 U616 ( .A1(G902), .A2(n496), .ZN(n600) );
  NOR2_X1 U617 ( .A1(n746), .A2(n600), .ZN(n497) );
  XOR2_X1 U618 ( .A(KEYINPUT104), .B(n497), .Z(n498) );
  NOR2_X1 U619 ( .A1(G900), .A2(n498), .ZN(n499) );
  XOR2_X1 U620 ( .A(KEYINPUT105), .B(n499), .Z(n500) );
  NOR2_X1 U621 ( .A1(n602), .A2(n500), .ZN(n562) );
  XNOR2_X1 U622 ( .A(KEYINPUT21), .B(n503), .ZN(n670) );
  NOR2_X1 U623 ( .A1(n562), .A2(n670), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(KEYINPUT70), .ZN(n514) );
  XNOR2_X1 U625 ( .A(G128), .B(G140), .ZN(n505) );
  XNOR2_X1 U626 ( .A(n505), .B(KEYINPUT24), .ZN(n507) );
  XNOR2_X1 U627 ( .A(n743), .B(n508), .ZN(n726) );
  NAND2_X1 U628 ( .A1(n509), .A2(G217), .ZN(n511) );
  NAND2_X1 U629 ( .A1(n514), .A2(n669), .ZN(n552) );
  XNOR2_X1 U630 ( .A(KEYINPUT13), .B(G475), .ZN(n526) );
  XNOR2_X1 U631 ( .A(n516), .B(n515), .ZN(n517) );
  NAND2_X1 U632 ( .A1(n518), .A2(G214), .ZN(n519) );
  XNOR2_X1 U633 ( .A(n535), .B(G113), .ZN(n522) );
  XNOR2_X1 U634 ( .A(G143), .B(KEYINPUT11), .ZN(n520) );
  NOR2_X1 U635 ( .A1(G902), .A2(n724), .ZN(n525) );
  XOR2_X1 U636 ( .A(n527), .B(KEYINPUT7), .Z(n529) );
  XNOR2_X1 U637 ( .A(n529), .B(n528), .ZN(n530) );
  NAND2_X1 U638 ( .A1(G217), .A2(n531), .ZN(n532) );
  NOR2_X1 U639 ( .A1(n725), .A2(G902), .ZN(n533) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n557) );
  NOR2_X1 U641 ( .A1(n552), .A2(n557), .ZN(n534) );
  NAND2_X1 U642 ( .A1(G227), .A2(n746), .ZN(n538) );
  XNOR2_X1 U643 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U644 ( .A(n541), .B(n540), .ZN(n542) );
  NAND2_X1 U645 ( .A1(n667), .A2(n656), .ZN(n545) );
  NOR2_X1 U646 ( .A1(n588), .A2(n545), .ZN(n546) );
  XNOR2_X1 U647 ( .A(n546), .B(KEYINPUT43), .ZN(n547) );
  XOR2_X1 U648 ( .A(KEYINPUT41), .B(KEYINPUT111), .Z(n551) );
  NAND2_X1 U649 ( .A1(n656), .A2(n657), .ZN(n549) );
  XNOR2_X1 U650 ( .A(n549), .B(KEYINPUT110), .ZN(n661) );
  XOR2_X1 U651 ( .A(n357), .B(KEYINPUT100), .Z(n659) );
  NOR2_X1 U652 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U653 ( .A(KEYINPUT28), .B(n554), .Z(n555) );
  NOR2_X1 U654 ( .A1(n560), .A2(n555), .ZN(n581) );
  NAND2_X1 U655 ( .A1(n653), .A2(n581), .ZN(n556) );
  XOR2_X1 U656 ( .A(KEYINPUT109), .B(KEYINPUT40), .Z(n567) );
  INV_X1 U657 ( .A(n557), .ZN(n710) );
  NOR2_X1 U658 ( .A1(KEYINPUT75), .A2(n559), .ZN(n565) );
  INV_X1 U659 ( .A(KEYINPUT75), .ZN(n561) );
  NAND2_X1 U660 ( .A1(n569), .A2(n580), .ZN(n570) );
  XNOR2_X1 U661 ( .A(n570), .B(KEYINPUT107), .ZN(n573) );
  NAND2_X1 U662 ( .A1(n571), .A2(n576), .ZN(n572) );
  XNOR2_X1 U663 ( .A(n572), .B(KEYINPUT103), .ZN(n622) );
  NAND2_X1 U664 ( .A1(n573), .A2(n622), .ZN(n574) );
  NOR2_X1 U665 ( .A1(n576), .A2(n575), .ZN(n712) );
  XNOR2_X1 U666 ( .A(KEYINPUT98), .B(n712), .ZN(n595) );
  NAND2_X1 U667 ( .A1(KEYINPUT47), .A2(n660), .ZN(n577) );
  NAND2_X1 U668 ( .A1(n758), .A2(n577), .ZN(n579) );
  NAND2_X1 U669 ( .A1(n581), .A2(n605), .ZN(n585) );
  NAND2_X1 U670 ( .A1(KEYINPUT47), .A2(n585), .ZN(n582) );
  NAND2_X1 U671 ( .A1(n583), .A2(n582), .ZN(n584) );
  INV_X1 U672 ( .A(n585), .ZN(n708) );
  NOR2_X1 U673 ( .A1(KEYINPUT47), .A2(n660), .ZN(n586) );
  NAND2_X1 U674 ( .A1(n708), .A2(n586), .ZN(n587) );
  XNOR2_X1 U675 ( .A(KEYINPUT112), .B(n588), .ZN(n589) );
  NOR2_X1 U676 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U677 ( .A(n593), .B(KEYINPUT82), .ZN(n597) );
  AND2_X1 U678 ( .A1(n595), .A2(n594), .ZN(n718) );
  INV_X1 U679 ( .A(KEYINPUT44), .ZN(n626) );
  NAND2_X1 U680 ( .A1(n626), .A2(KEYINPUT86), .ZN(n618) );
  XOR2_X1 U681 ( .A(KEYINPUT67), .B(KEYINPUT72), .Z(n599) );
  XNOR2_X1 U682 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n598) );
  XNOR2_X1 U683 ( .A(n599), .B(n598), .ZN(n611) );
  INV_X1 U684 ( .A(G953), .ZN(n736) );
  NOR2_X1 U685 ( .A1(G898), .A2(n736), .ZN(n732) );
  INV_X1 U686 ( .A(n600), .ZN(n601) );
  NAND2_X1 U687 ( .A1(n732), .A2(n601), .ZN(n604) );
  INV_X1 U688 ( .A(n602), .ZN(n603) );
  NAND2_X1 U689 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U690 ( .A1(n606), .A2(n605), .ZN(n608) );
  XOR2_X1 U691 ( .A(KEYINPUT68), .B(KEYINPUT0), .Z(n607) );
  XNOR2_X2 U692 ( .A(n608), .B(n607), .ZN(n634) );
  NOR2_X1 U693 ( .A1(n670), .A2(n659), .ZN(n609) );
  NAND2_X1 U694 ( .A1(n634), .A2(n609), .ZN(n610) );
  NOR2_X1 U695 ( .A1(n450), .A2(n612), .ZN(n702) );
  OR2_X1 U696 ( .A1(n450), .A2(n667), .ZN(n613) );
  XNOR2_X1 U697 ( .A(KEYINPUT101), .B(n613), .ZN(n615) );
  NAND2_X1 U698 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U699 ( .A1(n616), .A2(n619), .ZN(n617) );
  XNOR2_X1 U700 ( .A(n617), .B(KEYINPUT32), .ZN(n755) );
  INV_X1 U701 ( .A(n634), .ZN(n631) );
  INV_X1 U702 ( .A(n619), .ZN(n627) );
  NOR2_X1 U703 ( .A1(n627), .A2(n620), .ZN(n621) );
  INV_X1 U704 ( .A(n754), .ZN(n625) );
  NAND2_X1 U705 ( .A1(n450), .A2(n627), .ZN(n628) );
  NOR2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n696) );
  NAND2_X1 U707 ( .A1(n407), .A2(n630), .ZN(n675) );
  NOR2_X1 U708 ( .A1(n631), .A2(n675), .ZN(n633) );
  XOR2_X1 U709 ( .A(KEYINPUT94), .B(KEYINPUT31), .Z(n632) );
  XNOR2_X1 U710 ( .A(n633), .B(n632), .ZN(n713) );
  NAND2_X1 U711 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U712 ( .A1(n636), .A2(n407), .ZN(n637) );
  XOR2_X1 U713 ( .A(KEYINPUT93), .B(n637), .Z(n698) );
  NOR2_X1 U714 ( .A1(n713), .A2(n698), .ZN(n638) );
  NOR2_X1 U715 ( .A1(n660), .A2(n638), .ZN(n639) );
  NOR2_X1 U716 ( .A1(n696), .A2(n639), .ZN(n640) );
  XNOR2_X1 U717 ( .A(n646), .B(KEYINPUT80), .ZN(n643) );
  AND2_X1 U718 ( .A1(KEYINPUT2), .A2(n643), .ZN(n644) );
  NAND2_X1 U719 ( .A1(n655), .A2(n644), .ZN(n647) );
  INV_X1 U720 ( .A(KEYINPUT2), .ZN(n645) );
  XNOR2_X1 U721 ( .A(KEYINPUT54), .B(KEYINPUT122), .ZN(n650) );
  XNOR2_X1 U722 ( .A(n648), .B(KEYINPUT55), .ZN(n649) );
  INV_X1 U723 ( .A(KEYINPUT56), .ZN(n651) );
  INV_X1 U724 ( .A(n653), .ZN(n679) );
  NOR2_X1 U725 ( .A1(n679), .A2(n665), .ZN(n654) );
  NOR2_X1 U726 ( .A1(G953), .A2(n654), .ZN(n690) );
  AND2_X1 U727 ( .A1(KEYINPUT2), .A2(n655), .ZN(n688) );
  NOR2_X1 U728 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n663) );
  NOR2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U731 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U732 ( .A1(n665), .A2(n664), .ZN(n682) );
  NAND2_X1 U733 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U734 ( .A(n668), .B(KEYINPUT50), .ZN(n674) );
  NAND2_X1 U735 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U736 ( .A(KEYINPUT49), .B(n671), .ZN(n672) );
  NOR2_X1 U737 ( .A1(n407), .A2(n672), .ZN(n673) );
  NAND2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n676) );
  NAND2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n678) );
  XOR2_X1 U740 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n677) );
  XNOR2_X1 U741 ( .A(n678), .B(n677), .ZN(n680) );
  NOR2_X1 U742 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U743 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U744 ( .A(n683), .B(KEYINPUT120), .ZN(n684) );
  XNOR2_X1 U745 ( .A(KEYINPUT52), .B(n684), .ZN(n685) );
  NOR2_X1 U746 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U748 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U749 ( .A1(n652), .A2(n691), .ZN(n694) );
  INV_X1 U750 ( .A(KEYINPUT121), .ZN(n692) );
  XNOR2_X1 U751 ( .A(n692), .B(KEYINPUT53), .ZN(n693) );
  XOR2_X1 U752 ( .A(G101), .B(n696), .Z(G3) );
  NAND2_X1 U753 ( .A1(n698), .A2(n710), .ZN(n697) );
  XNOR2_X1 U754 ( .A(n697), .B(G104), .ZN(G6) );
  XOR2_X1 U755 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n700) );
  NAND2_X1 U756 ( .A1(n698), .A2(n712), .ZN(n699) );
  XNOR2_X1 U757 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U758 ( .A(G107), .B(n701), .ZN(G9) );
  XOR2_X1 U759 ( .A(G110), .B(n702), .Z(n703) );
  XNOR2_X1 U760 ( .A(KEYINPUT114), .B(n703), .ZN(G12) );
  XOR2_X1 U761 ( .A(KEYINPUT29), .B(KEYINPUT116), .Z(n705) );
  NAND2_X1 U762 ( .A1(n708), .A2(n712), .ZN(n704) );
  XNOR2_X1 U763 ( .A(n705), .B(n704), .ZN(n707) );
  XOR2_X1 U764 ( .A(G128), .B(KEYINPUT115), .Z(n706) );
  XNOR2_X1 U765 ( .A(n707), .B(n706), .ZN(G30) );
  NAND2_X1 U766 ( .A1(n708), .A2(n710), .ZN(n709) );
  XNOR2_X1 U767 ( .A(n709), .B(G146), .ZN(G48) );
  NAND2_X1 U768 ( .A1(n713), .A2(n710), .ZN(n711) );
  XNOR2_X1 U769 ( .A(n711), .B(G113), .ZN(G15) );
  NAND2_X1 U770 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U771 ( .A(n714), .B(G116), .ZN(G18) );
  XNOR2_X1 U772 ( .A(n715), .B(KEYINPUT37), .ZN(n716) );
  XNOR2_X1 U773 ( .A(n716), .B(KEYINPUT118), .ZN(n717) );
  XNOR2_X1 U774 ( .A(G125), .B(n717), .ZN(G27) );
  XOR2_X1 U775 ( .A(G134), .B(n718), .Z(G36) );
  XOR2_X1 U776 ( .A(G140), .B(n719), .Z(G42) );
  XOR2_X1 U777 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n721) );
  NAND2_X1 U778 ( .A1(G469), .A2(n727), .ZN(n720) );
  NOR2_X1 U779 ( .A1(n730), .A2(n723), .ZN(G54) );
  NAND2_X1 U780 ( .A1(G217), .A2(n727), .ZN(n728) );
  XNOR2_X1 U781 ( .A(n726), .B(n728), .ZN(n729) );
  NOR2_X1 U782 ( .A1(n730), .A2(n729), .ZN(G66) );
  NOR2_X1 U783 ( .A1(n731), .A2(n732), .ZN(n741) );
  NAND2_X1 U784 ( .A1(G953), .A2(G224), .ZN(n733) );
  XNOR2_X1 U785 ( .A(KEYINPUT61), .B(n733), .ZN(n734) );
  NAND2_X1 U786 ( .A1(n734), .A2(G898), .ZN(n735) );
  XNOR2_X1 U787 ( .A(KEYINPUT124), .B(n735), .ZN(n739) );
  XOR2_X1 U788 ( .A(KEYINPUT125), .B(n737), .Z(n738) );
  NAND2_X1 U789 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U790 ( .A(n741), .B(n740), .ZN(G69) );
  XOR2_X1 U791 ( .A(n743), .B(KEYINPUT126), .Z(n744) );
  XOR2_X1 U792 ( .A(n742), .B(n744), .Z(n748) );
  XOR2_X1 U793 ( .A(n748), .B(n745), .Z(n747) );
  NAND2_X1 U794 ( .A1(n747), .A2(n746), .ZN(n752) );
  XNOR2_X1 U795 ( .A(G227), .B(n748), .ZN(n749) );
  NAND2_X1 U796 ( .A1(n749), .A2(G900), .ZN(n750) );
  NAND2_X1 U797 ( .A1(G953), .A2(n750), .ZN(n751) );
  NAND2_X1 U798 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U799 ( .A(KEYINPUT127), .B(n753), .Z(G72) );
  XNOR2_X1 U800 ( .A(G122), .B(n754), .ZN(G24) );
  XOR2_X1 U801 ( .A(G119), .B(n755), .Z(G21) );
  XNOR2_X1 U802 ( .A(n756), .B(G137), .ZN(G39) );
  XNOR2_X1 U803 ( .A(G131), .B(n757), .ZN(G33) );
  XOR2_X1 U804 ( .A(n758), .B(G143), .Z(n759) );
  XNOR2_X1 U805 ( .A(KEYINPUT117), .B(n759), .ZN(G45) );
endmodule

