//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1310, new_n1311, new_n1312, new_n1314, new_n1315,
    new_n1316, new_n1317, new_n1318, new_n1319, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383,
    new_n1384, new_n1385, new_n1386, new_n1387, new_n1388, new_n1389;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(KEYINPUT64), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n201), .B(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AND2_X1   g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(G58), .A2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G107), .ZN(new_n224));
  INV_X1    g0024(.A(G264), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n206), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n209), .B1(new_n211), .B2(new_n214), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT66), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n233), .B(new_n234), .Z(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(G274), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G33), .A2(G41), .ZN(new_n248));
  AOI21_X1  g0048(.A(new_n247), .B1(new_n210), .B2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n250), .B1(G41), .B2(G45), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n210), .A2(new_n248), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G238), .A3(new_n251), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT73), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n253), .A2(KEYINPUT73), .A3(new_n255), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  OAI21_X1  g0061(.A(KEYINPUT67), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT67), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G226), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(G1698), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n262), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT72), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G97), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n262), .A2(new_n268), .A3(G232), .A4(G1698), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n262), .A2(new_n268), .A3(KEYINPUT72), .A4(new_n270), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n273), .A2(new_n274), .A3(new_n275), .A4(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n254), .ZN(new_n278));
  AOI221_X4 g0078(.A(KEYINPUT13), .B1(new_n258), .B2(new_n259), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT13), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n277), .A2(new_n278), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n258), .A2(new_n259), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G169), .ZN(new_n285));
  OAI21_X1  g0085(.A(KEYINPUT14), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT14), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n287), .B(G169), .C1(new_n279), .C2(new_n283), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT74), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n289), .B1(new_n284), .B2(G179), .ZN(new_n290));
  INV_X1    g0090(.A(G179), .ZN(new_n291));
  NOR4_X1   g0091(.A1(new_n279), .A2(new_n283), .A3(KEYINPUT74), .A4(new_n291), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n286), .B(new_n288), .C1(new_n290), .C2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G1), .A2(G13), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G50), .ZN(new_n299));
  INV_X1    g0099(.A(G20), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n298), .A2(new_n299), .B1(new_n300), .B2(G68), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(G33), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(new_n222), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n296), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT11), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n305), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n250), .A2(G13), .A3(G20), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n216), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT12), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n309), .A2(new_n296), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n312), .B(G68), .C1(G1), .C2(new_n300), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n306), .A2(new_n307), .A3(new_n311), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n293), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n284), .A2(G190), .ZN(new_n317));
  INV_X1    g0117(.A(new_n314), .ZN(new_n318));
  OAI21_X1  g0118(.A(G200), .B1(new_n279), .B2(new_n283), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n262), .A2(new_n268), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n254), .B1(new_n323), .B2(new_n222), .ZN(new_n324));
  MUX2_X1   g0124(.A(G222), .B(G223), .S(G1698), .Z(new_n325));
  OAI21_X1  g0125(.A(new_n324), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n253), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n254), .A2(new_n251), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n327), .B1(G226), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G190), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(G200), .B2(new_n331), .ZN(new_n334));
  INV_X1    g0134(.A(new_n312), .ZN(new_n335));
  OAI21_X1  g0135(.A(G50), .B1(new_n300), .B2(G1), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n335), .A2(new_n336), .B1(G50), .B2(new_n308), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n203), .A2(G20), .ZN(new_n339));
  XOR2_X1   g0139(.A(KEYINPUT8), .B(G58), .Z(new_n340));
  INV_X1    g0140(.A(new_n302), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n340), .A2(new_n341), .B1(G150), .B2(new_n297), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n294), .A2(new_n295), .ZN(new_n344));
  OAI211_X1 g0144(.A(KEYINPUT71), .B(new_n338), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT71), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n344), .B1(new_n339), .B2(new_n342), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n346), .B1(new_n347), .B2(new_n337), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT9), .ZN(new_n349));
  AND3_X1   g0149(.A1(new_n345), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n349), .B1(new_n345), .B2(new_n348), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n334), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT10), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT10), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n334), .B(new_n354), .C1(new_n350), .C2(new_n351), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n323), .A2(G107), .ZN(new_n357));
  INV_X1    g0157(.A(G1698), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n262), .A2(new_n268), .A3(G232), .A4(new_n358), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n262), .A2(new_n268), .A3(G238), .A4(G1698), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n357), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT68), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT68), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n357), .A2(new_n363), .A3(new_n359), .A4(new_n360), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(new_n278), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT69), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n327), .B1(G244), .B2(new_n329), .ZN(new_n367));
  AND3_X1   g0167(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n366), .B1(new_n365), .B2(new_n367), .ZN(new_n369));
  OAI21_X1  g0169(.A(G190), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n365), .A2(new_n367), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT69), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(G200), .A3(new_n373), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n340), .A2(new_n297), .B1(G20), .B2(G77), .ZN(new_n375));
  XNOR2_X1  g0175(.A(KEYINPUT15), .B(G87), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n375), .A2(KEYINPUT70), .B1(new_n341), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(KEYINPUT70), .B2(new_n375), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n296), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n300), .A2(G1), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n381), .A2(new_n222), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n312), .A2(new_n382), .B1(new_n222), .B2(new_n309), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n370), .A2(new_n374), .A3(new_n380), .A4(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n291), .B1(new_n368), .B2(new_n369), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n372), .A2(new_n285), .A3(new_n373), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n380), .A2(new_n383), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n347), .A2(new_n337), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n331), .A2(G179), .ZN(new_n390));
  AOI211_X1 g0190(.A(new_n389), .B(new_n390), .C1(new_n285), .C2(new_n331), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n356), .A2(new_n384), .A3(new_n388), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n269), .A2(G1698), .ZN(new_n394));
  OAI221_X1 g0194(.A(new_n394), .B1(G223), .B2(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G87), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n254), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G232), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n253), .B1(new_n328), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n400), .A2(new_n285), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n397), .A2(new_n399), .A3(new_n291), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G58), .A2(G68), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(G20), .B1(new_n405), .B2(new_n212), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT76), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n297), .A2(G159), .ZN(new_n409));
  OAI211_X1 g0209(.A(KEYINPUT76), .B(G20), .C1(new_n405), .C2(new_n212), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  XNOR2_X1  g0211(.A(KEYINPUT3), .B(G33), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n300), .A2(KEYINPUT7), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT75), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n260), .B2(new_n261), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n265), .A2(KEYINPUT75), .A3(new_n267), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(new_n417), .A3(new_n300), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT7), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n414), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n411), .B(KEYINPUT16), .C1(new_n420), .C2(new_n216), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n422));
  AOI21_X1  g0222(.A(G20), .B1(new_n262), .B2(new_n268), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n423), .A2(KEYINPUT7), .B1(new_n412), .B2(new_n413), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n422), .B1(new_n424), .B2(G68), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n421), .B(new_n296), .C1(new_n425), .C2(KEYINPUT16), .ZN(new_n426));
  INV_X1    g0226(.A(new_n340), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n335), .A2(new_n381), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n428), .B1(new_n309), .B2(new_n427), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n403), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT18), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI211_X1 g0232(.A(KEYINPUT18), .B(new_n403), .C1(new_n426), .C2(new_n429), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n400), .A2(new_n332), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(G200), .B2(new_n400), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n426), .A2(new_n429), .A3(new_n436), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n437), .B(KEYINPUT17), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n393), .A2(new_n439), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n322), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G45), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(G1), .ZN(new_n444));
  NAND2_X1  g0244(.A1(KEYINPUT5), .A2(G41), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n444), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n448), .A2(G270), .A3(new_n254), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n250), .A2(G45), .ZN(new_n450));
  OR2_X1    g0250(.A1(KEYINPUT5), .A2(G41), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(new_n445), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n249), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT67), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n266), .B1(new_n265), .B2(new_n267), .ZN(new_n456));
  OAI21_X1  g0256(.A(G303), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G257), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n358), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n225), .A2(G1698), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n459), .B(new_n460), .C1(new_n260), .C2(new_n261), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n454), .B1(new_n462), .B2(new_n278), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G179), .ZN(new_n464));
  INV_X1    g0264(.A(G303), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n465), .B1(new_n262), .B2(new_n268), .ZN(new_n466));
  INV_X1    g0266(.A(new_n461), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n278), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n449), .A2(new_n453), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(KEYINPUT21), .A3(G169), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n464), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n309), .A2(G116), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n344), .B(new_n308), .C1(G1), .C2(new_n264), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(G116), .ZN(new_n475));
  AOI21_X1  g0275(.A(G20), .B1(new_n264), .B2(G97), .ZN(new_n476));
  INV_X1    g0276(.A(G283), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n476), .B1(new_n264), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G116), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G20), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n296), .A2(KEYINPUT80), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT80), .B1(new_n296), .B2(new_n480), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n478), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT20), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(KEYINPUT20), .B(new_n478), .C1(new_n481), .C2(new_n482), .ZN(new_n486));
  AOI211_X1 g0286(.A(KEYINPUT81), .B(new_n475), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT81), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n485), .A2(new_n486), .ZN(new_n489));
  INV_X1    g0289(.A(new_n475), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n472), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n296), .A2(new_n480), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT80), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n296), .A2(KEYINPUT80), .A3(new_n480), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(KEYINPUT20), .B1(new_n497), .B2(new_n478), .ZN(new_n498));
  INV_X1    g0298(.A(new_n486), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n490), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT81), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n489), .A2(new_n488), .A3(new_n490), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n470), .A2(G200), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n463), .A2(G190), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n501), .A2(new_n502), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n470), .A2(G169), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n506), .B1(new_n501), .B2(new_n502), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n492), .B(new_n505), .C1(new_n507), .C2(KEYINPUT21), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT82), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n506), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n491), .B2(new_n487), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT21), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n514), .A2(KEYINPUT82), .A3(new_n492), .A4(new_n505), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n308), .A2(G97), .ZN(new_n518));
  INV_X1    g0318(.A(new_n474), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n518), .B1(new_n519), .B2(G97), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT6), .ZN(new_n522));
  INV_X1    g0322(.A(G97), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n522), .A2(new_n523), .A3(G107), .ZN(new_n524));
  XNOR2_X1  g0324(.A(G97), .B(G107), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n524), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n526), .A2(new_n300), .B1(new_n222), .B2(new_n298), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n323), .A2(new_n300), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n414), .B1(new_n529), .B2(new_n419), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n528), .B1(new_n530), .B2(new_n224), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n521), .B1(new_n531), .B2(new_n296), .ZN(new_n532));
  OAI211_X1 g0332(.A(G244), .B(new_n358), .C1(new_n260), .C2(new_n261), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT4), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n533), .A2(new_n534), .B1(G33), .B2(G283), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n358), .A2(G244), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n536), .A2(new_n534), .B1(new_n219), .B2(new_n358), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n537), .A2(new_n262), .A3(new_n268), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n278), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT77), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n448), .A2(new_n541), .A3(G257), .A4(new_n254), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n448), .A2(G257), .A3(new_n254), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n543), .A2(KEYINPUT77), .B1(new_n249), .B2(new_n452), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n540), .A2(G190), .A3(new_n542), .A4(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(KEYINPUT77), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n546), .A2(new_n453), .A3(new_n542), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n254), .B1(new_n535), .B2(new_n538), .ZN(new_n548));
  OAI21_X1  g0348(.A(G200), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n532), .A2(KEYINPUT78), .A3(new_n545), .A4(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT78), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n540), .A2(G179), .A3(new_n542), .A4(new_n544), .ZN(new_n552));
  OAI21_X1  g0352(.A(G169), .B1(new_n547), .B2(new_n548), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n527), .B1(new_n424), .B2(G107), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n520), .B1(new_n555), .B2(new_n344), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n551), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n545), .A2(new_n549), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(new_n556), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n550), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n309), .A2(KEYINPUT25), .A3(new_n224), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT83), .ZN(new_n562));
  XNOR2_X1  g0362(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT84), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n309), .A2(new_n224), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT25), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI211_X1 g0367(.A(KEYINPUT84), .B(KEYINPUT25), .C1(new_n309), .C2(new_n224), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI22_X1  g0369(.A1(new_n563), .A2(new_n569), .B1(new_n224), .B2(new_n474), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NOR3_X1   g0371(.A1(new_n218), .A2(KEYINPUT22), .A3(G20), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n262), .A2(new_n268), .A3(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n300), .B(G87), .C1(new_n260), .C2(new_n261), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT22), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT24), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G33), .A2(G116), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n578), .A2(G20), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT23), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n300), .B2(G107), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n224), .A2(KEYINPUT23), .A3(G20), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n576), .A2(new_n577), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n577), .B1(new_n576), .B2(new_n583), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n296), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n571), .A2(new_n587), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n452), .A2(new_n278), .A3(new_n225), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(G294), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n264), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(G250), .A2(G1698), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n458), .B2(G1698), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n592), .B1(new_n594), .B2(new_n412), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n278), .B1(new_n595), .B2(KEYINPUT85), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n219), .A2(new_n358), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n458), .A2(G1698), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n597), .B(new_n598), .C1(new_n260), .C2(new_n261), .ZN(new_n599));
  INV_X1    g0399(.A(new_n592), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT85), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n453), .B(new_n590), .C1(new_n596), .C2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT86), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(new_n605), .A3(G169), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n254), .B1(new_n601), .B2(new_n602), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n595), .A2(KEYINPUT85), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n589), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(G179), .A3(new_n453), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n605), .B1(new_n604), .B2(G169), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n588), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(G200), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n604), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n609), .A2(new_n332), .A3(new_n453), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n616), .A3(KEYINPUT87), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n576), .A2(new_n583), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT24), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n584), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n570), .B1(new_n620), .B2(new_n296), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT87), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n604), .A2(new_n622), .A3(new_n614), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n617), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT19), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n300), .B1(new_n274), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(G97), .A2(G107), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n218), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n300), .B(G68), .C1(new_n260), .C2(new_n261), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n625), .B1(new_n302), .B2(new_n523), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n296), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n312), .B(new_n377), .C1(G1), .C2(new_n264), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n376), .A2(new_n309), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n217), .A2(new_n358), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n223), .A2(G1698), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n637), .B(new_n638), .C1(new_n260), .C2(new_n261), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n254), .B1(new_n639), .B2(new_n578), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n254), .A2(G274), .A3(new_n444), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n219), .B1(new_n250), .B2(G45), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n254), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n285), .B1(new_n640), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n639), .A2(new_n578), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n278), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n249), .A2(new_n444), .B1(new_n254), .B2(new_n642), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(new_n291), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n636), .A2(new_n645), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(G200), .B1(new_n640), .B2(new_n644), .ZN(new_n651));
  NOR2_X1   g0451(.A1(G238), .A2(G1698), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(new_n223), .B2(G1698), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n653), .A2(new_n412), .B1(G33), .B2(G116), .ZN(new_n654));
  OAI211_X1 g0454(.A(G190), .B(new_n648), .C1(new_n654), .C2(new_n254), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n632), .A2(new_n296), .B1(new_n309), .B2(new_n376), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n519), .A2(G87), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n651), .A2(new_n655), .A3(new_n656), .A4(new_n657), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n650), .A2(new_n658), .A3(KEYINPUT79), .ZN(new_n659));
  AOI21_X1  g0459(.A(KEYINPUT79), .B1(new_n650), .B2(new_n658), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n613), .A2(new_n624), .A3(new_n661), .ZN(new_n662));
  NOR4_X1   g0462(.A1(new_n442), .A2(new_n517), .A3(new_n560), .A4(new_n662), .ZN(G372));
  INV_X1    g0463(.A(new_n438), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n320), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n664), .B1(new_n315), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT90), .ZN(new_n668));
  INV_X1    g0468(.A(new_n434), .ZN(new_n669));
  OR3_X1    g0469(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n668), .B1(new_n667), .B2(new_n669), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(new_n356), .A3(new_n671), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n672), .A2(new_n392), .ZN(new_n673));
  INV_X1    g0473(.A(new_n560), .ZN(new_n674));
  INV_X1    g0474(.A(new_n650), .ZN(new_n675));
  XOR2_X1   g0475(.A(new_n651), .B(KEYINPUT88), .Z(new_n676));
  NAND2_X1  g0476(.A1(new_n656), .A2(new_n657), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n640), .A2(new_n644), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n677), .B1(G190), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n675), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n624), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n514), .A2(new_n613), .A3(new_n492), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n674), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n554), .A2(new_n556), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n661), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT26), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT89), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n532), .B1(new_n688), .B2(new_n554), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT26), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT89), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n689), .A2(new_n680), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n687), .A2(new_n650), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n441), .B1(new_n683), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n673), .A2(new_n694), .ZN(G369));
  NAND3_X1  g0495(.A1(new_n250), .A2(new_n300), .A3(G13), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G213), .A3(new_n698), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT91), .Z(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G343), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n704), .B1(new_n502), .B2(new_n501), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n517), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n705), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n514), .B2(new_n492), .ZN(new_n708));
  OAI21_X1  g0508(.A(G330), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n613), .A2(new_n624), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n621), .B2(new_n704), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n613), .B2(new_n704), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n703), .B1(new_n514), .B2(new_n492), .ZN(new_n715));
  INV_X1    g0515(.A(new_n613), .ZN(new_n716));
  AOI22_X1  g0516(.A1(new_n715), .A2(new_n711), .B1(new_n716), .B2(new_n704), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n714), .A2(new_n717), .ZN(G399));
  NOR2_X1   g0518(.A1(new_n628), .A2(G116), .ZN(new_n719));
  XOR2_X1   g0519(.A(new_n719), .B(KEYINPUT92), .Z(new_n720));
  INV_X1    g0520(.A(new_n207), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G41), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n720), .A2(new_n250), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n214), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(new_n722), .ZN(new_n725));
  XOR2_X1   g0525(.A(new_n725), .B(KEYINPUT28), .Z(new_n726));
  INV_X1    g0526(.A(KEYINPUT29), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT96), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n554), .A2(new_n688), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n729), .A2(new_n691), .A3(new_n556), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n690), .B1(new_n730), .B2(new_n680), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n661), .A2(new_n685), .A3(new_n690), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n650), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n728), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n689), .A2(new_n680), .A3(new_n691), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT26), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n736), .A2(KEYINPUT96), .A3(new_n650), .A4(new_n732), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n560), .A2(KEYINPUT97), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT97), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n550), .B(new_n739), .C1(new_n557), .C2(new_n559), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n738), .A2(new_n682), .A3(new_n681), .A4(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n734), .A2(new_n737), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n727), .B1(new_n742), .B2(new_n704), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n704), .B1(new_n683), .B2(new_n693), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(KEYINPUT29), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT93), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(KEYINPUT30), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n463), .A2(new_n609), .A3(G179), .A4(new_n678), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n547), .A2(new_n548), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n748), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n291), .B1(new_n640), .B2(new_n644), .ZN(new_n753));
  OAI21_X1  g0553(.A(KEYINPUT94), .B1(new_n463), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT94), .ZN(new_n755));
  AOI21_X1  g0555(.A(G179), .B1(new_n647), .B2(new_n648), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n470), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n754), .A2(new_n751), .A3(new_n604), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n607), .A2(new_n608), .ZN(new_n759));
  AND3_X1   g0559(.A1(new_n759), .A2(new_n590), .A3(new_n678), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n470), .A2(new_n291), .ZN(new_n761));
  INV_X1    g0561(.A(new_n748), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n760), .A2(new_n761), .A3(new_n750), .A4(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n752), .A2(new_n758), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n703), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT31), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n764), .A2(KEYINPUT31), .A3(new_n703), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n662), .A2(new_n560), .A3(new_n703), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n769), .B1(new_n516), .B2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G330), .ZN(new_n772));
  OAI21_X1  g0572(.A(KEYINPUT95), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n516), .A2(new_n770), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n767), .A2(new_n768), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT95), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n776), .A2(new_n777), .A3(G330), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n746), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n726), .B1(new_n781), .B2(G1), .ZN(G364));
  OAI21_X1  g0582(.A(new_n210), .B1(new_n300), .B2(G169), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n783), .A2(KEYINPUT99), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(KEYINPUT99), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n300), .A2(new_n332), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n787), .A2(G179), .A3(G200), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G179), .A2(G200), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n300), .B1(new_n790), .B2(G190), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n789), .A2(G326), .B1(new_n792), .B2(G294), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n787), .A2(new_n291), .A3(G200), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n793), .B(new_n323), .C1(new_n465), .C2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n300), .A2(G190), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n796), .A2(new_n291), .A3(G200), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n796), .A2(new_n790), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n798), .A2(G283), .B1(new_n799), .B2(G329), .ZN(new_n800));
  INV_X1    g0600(.A(G322), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n291), .A2(G200), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n787), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n332), .A2(G20), .A3(G179), .A4(G200), .ZN(new_n804));
  XOR2_X1   g0604(.A(KEYINPUT33), .B(G317), .Z(new_n805));
  OAI221_X1 g0605(.A(new_n800), .B1(new_n801), .B2(new_n803), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n802), .A2(new_n796), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n807), .A2(KEYINPUT100), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(KEYINPUT100), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n795), .B(new_n806), .C1(G311), .C2(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT101), .ZN(new_n812));
  INV_X1    g0612(.A(new_n794), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G87), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(new_n299), .B2(new_n788), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n323), .B(new_n815), .C1(G97), .C2(new_n792), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n810), .A2(G77), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n799), .A2(G159), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT32), .Z(new_n819));
  NAND2_X1  g0619(.A1(new_n798), .A2(G107), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n216), .B2(new_n804), .ZN(new_n821));
  INV_X1    g0621(.A(new_n803), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n821), .B1(G58), .B2(new_n822), .ZN(new_n823));
  AND4_X1   g0623(.A1(new_n816), .A2(new_n817), .A3(new_n819), .A4(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n786), .B1(new_n812), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n300), .A2(G13), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n250), .B1(new_n826), .B2(G45), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n722), .ZN(new_n829));
  NOR2_X1   g0629(.A1(G13), .A2(G33), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(G20), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n786), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n416), .A2(new_n417), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n721), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(G45), .B2(new_n214), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(G45), .B2(new_n245), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n323), .A2(new_n721), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  XOR2_X1   g0640(.A(G355), .B(KEYINPUT98), .Z(new_n841));
  OAI22_X1  g0641(.A1(new_n840), .A2(new_n841), .B1(G116), .B2(new_n207), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n833), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n825), .A2(new_n829), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n706), .A2(new_n708), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n844), .B1(new_n845), .B2(new_n832), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n710), .A2(new_n829), .ZN(new_n847));
  OR3_X1    g0647(.A1(new_n706), .A2(G330), .A3(new_n708), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G396));
  AND3_X1   g0650(.A1(new_n687), .A2(new_n650), .A3(new_n692), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n674), .A2(new_n682), .A3(new_n681), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n703), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n388), .A2(new_n703), .ZN(new_n854));
  INV_X1    g0654(.A(new_n387), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n384), .B1(new_n855), .B2(new_n704), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n854), .B1(new_n856), .B2(new_n388), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n665), .A2(new_n704), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n368), .A2(new_n369), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n387), .B1(new_n860), .B2(G200), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n861), .A2(new_n370), .B1(new_n387), .B2(new_n703), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n859), .B1(new_n862), .B2(new_n665), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n744), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n858), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n829), .B1(new_n779), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n779), .B2(new_n865), .ZN(new_n867));
  INV_X1    g0667(.A(new_n829), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n786), .A2(new_n830), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n868), .B1(new_n869), .B2(new_n222), .ZN(new_n870));
  INV_X1    g0670(.A(new_n786), .ZN(new_n871));
  INV_X1    g0671(.A(new_n804), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n822), .A2(G294), .B1(G283), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n798), .A2(G87), .ZN(new_n874));
  INV_X1    g0674(.A(G311), .ZN(new_n875));
  INV_X1    g0675(.A(new_n799), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n873), .B(new_n874), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  AOI22_X1  g0677(.A1(G107), .A2(new_n813), .B1(new_n789), .B2(G303), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n878), .B(new_n323), .C1(new_n523), .C2(new_n791), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n877), .B(new_n879), .C1(G116), .C2(new_n810), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n822), .A2(G143), .B1(G150), .B2(new_n872), .ZN(new_n881));
  INV_X1    g0681(.A(G137), .ZN(new_n882));
  INV_X1    g0682(.A(new_n810), .ZN(new_n883));
  INV_X1    g0683(.A(G159), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n881), .B1(new_n882), .B2(new_n788), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT34), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n813), .A2(G50), .B1(new_n792), .B2(G58), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n798), .A2(G68), .B1(new_n799), .B2(G132), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n887), .A2(new_n835), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n880), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  OAI221_X1 g0690(.A(new_n870), .B1(new_n871), .B2(new_n890), .C1(new_n857), .C2(new_n831), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n867), .A2(new_n891), .ZN(G384));
  NAND2_X1  g0692(.A1(new_n525), .A2(new_n522), .ZN(new_n893));
  INV_X1    g0693(.A(new_n524), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT35), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n211), .A2(new_n479), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n895), .B2(KEYINPUT35), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT102), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n899), .B2(new_n898), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT36), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n724), .A2(G77), .A3(new_n404), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n299), .A2(G68), .ZN(new_n904));
  AOI211_X1 g0704(.A(new_n250), .B(G13), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT105), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n434), .A2(new_n700), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n411), .B1(new_n420), .B2(new_n216), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT16), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n344), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n912), .A2(KEYINPUT103), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n421), .B1(new_n912), .B2(KEYINPUT103), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n429), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n403), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n915), .A2(new_n700), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n917), .A2(new_n918), .A3(new_n437), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT37), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n426), .A2(new_n429), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n916), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n700), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT37), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n922), .A2(new_n923), .A3(new_n924), .A4(new_n437), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT104), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n426), .A2(new_n429), .A3(new_n436), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n928), .A2(new_n430), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n929), .A2(KEYINPUT104), .A3(new_n924), .A4(new_n923), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n920), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n918), .B1(new_n434), .B2(new_n438), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n932), .A2(KEYINPUT38), .A3(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT38), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n919), .A2(KEYINPUT37), .B1(new_n927), .B2(new_n930), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n936), .B1(new_n937), .B2(new_n933), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n859), .B1(new_n744), .B2(new_n863), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n703), .A2(new_n314), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n315), .A2(new_n320), .A3(new_n941), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n314), .B(new_n703), .C1(new_n293), .C2(new_n321), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n907), .B(new_n909), .C1(new_n939), .C2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT39), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n937), .A2(new_n936), .A3(new_n933), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n929), .A2(new_n923), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(KEYINPUT37), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n931), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n923), .B1(new_n434), .B2(new_n438), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT38), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n947), .B1(new_n948), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n315), .A2(new_n703), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n935), .A2(new_n938), .A3(KEYINPUT39), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n946), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n858), .A2(new_n859), .B1(new_n942), .B2(new_n943), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n935), .A2(new_n938), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n908), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n963), .A2(new_n907), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n960), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n441), .B1(new_n745), .B2(new_n743), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n673), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n966), .B(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n944), .A2(new_n776), .A3(new_n857), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n970), .B1(new_n939), .B2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n971), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n927), .A2(new_n930), .B1(KEYINPUT37), .B2(new_n949), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n936), .B1(new_n974), .B2(new_n952), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n935), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n973), .A2(KEYINPUT40), .A3(new_n976), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n972), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n442), .B2(new_n771), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n978), .A2(new_n441), .A3(new_n776), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n980), .A2(G330), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n969), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n250), .B2(new_n826), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n969), .A2(new_n982), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n906), .B1(new_n984), .B2(new_n985), .ZN(G367));
  INV_X1    g0786(.A(new_n836), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n987), .A2(new_n238), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n833), .B1(new_n207), .B2(new_n376), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n990), .A2(new_n868), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n810), .A2(G50), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n876), .A2(new_n882), .B1(new_n884), .B2(new_n804), .ZN(new_n993));
  INV_X1    g0793(.A(G150), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n797), .A2(new_n222), .B1(new_n803), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n323), .B1(new_n813), .B2(G58), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n789), .A2(G143), .B1(new_n792), .B2(G68), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n992), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n834), .B1(new_n875), .B2(new_n788), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(G107), .B2(new_n792), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n797), .A2(new_n523), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n803), .A2(new_n465), .B1(new_n591), .B2(new_n804), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n1002), .B(new_n1003), .C1(G317), .C2(new_n799), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1001), .B(new_n1004), .C1(new_n477), .C2(new_n883), .ZN(new_n1005));
  AOI21_X1  g0805(.A(KEYINPUT112), .B1(new_n813), .B2(G116), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT46), .Z(new_n1007));
  OAI21_X1  g0807(.A(new_n999), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT47), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n786), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n703), .A2(new_n677), .ZN(new_n1012));
  MUX2_X1   g0812(.A(new_n675), .B(new_n680), .S(new_n1012), .Z(new_n1013));
  INV_X1    g0813(.A(new_n832), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n991), .B1(new_n1010), .B2(new_n1011), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT45), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n738), .B(new_n740), .C1(new_n532), .C2(new_n704), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n730), .A2(new_n703), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT110), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1019), .A2(new_n717), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1020), .B1(new_n1019), .B2(new_n717), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1016), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1023), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1025), .A2(KEYINPUT45), .A3(new_n1021), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT44), .ZN(new_n1027));
  OR3_X1    g0827(.A1(new_n1019), .A2(new_n1027), .A3(new_n717), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1027), .B1(new_n1019), .B2(new_n717), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1024), .A2(new_n1026), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n714), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT111), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n715), .A2(new_n711), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n713), .A2(new_n715), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n709), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1035), .B1(new_n713), .B2(new_n715), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1038), .B(G330), .C1(new_n706), .C2(new_n708), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1040), .A2(new_n780), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n714), .A2(new_n1024), .A3(new_n1026), .A4(new_n1030), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1034), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1033), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n781), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n722), .B(KEYINPUT41), .Z(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n828), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1019), .A2(new_n711), .A3(new_n715), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT42), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1049), .B(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT108), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1019), .B(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n685), .B1(new_n1053), .B2(new_n716), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1051), .B1(new_n1054), .B2(new_n703), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT107), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1056), .A2(KEYINPUT43), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(KEYINPUT43), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1013), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1019), .B(KEYINPUT108), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n714), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT109), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1055), .A2(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1059), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1049), .B(KEYINPUT42), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n684), .B1(new_n1060), .B2(new_n613), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1065), .B1(new_n1066), .B2(new_n704), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1013), .A2(KEYINPUT43), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1064), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1063), .A2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1063), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1015), .B1(new_n1048), .B2(new_n1075), .ZN(G387));
  AOI22_X1  g0876(.A1(new_n810), .A2(G303), .B1(G317), .B2(new_n822), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n789), .A2(G322), .B1(G311), .B2(new_n872), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1078), .A2(KEYINPUT113), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(KEYINPUT113), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1077), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT48), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n813), .A2(G294), .B1(new_n792), .B2(G283), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT49), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n797), .A2(new_n479), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1090), .B(new_n835), .C1(G326), .C2(new_n799), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1088), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n876), .A2(new_n994), .B1(new_n427), .B2(new_n804), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1002), .B(new_n1093), .C1(G50), .C2(new_n822), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n834), .B1(G159), .B2(new_n789), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n813), .A2(G77), .B1(new_n792), .B2(new_n377), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n810), .A2(G68), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n871), .B1(new_n1092), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n987), .B1(new_n235), .B2(G45), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n720), .B2(new_n839), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n427), .A2(G50), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT50), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n443), .B1(new_n216), .B2(new_n222), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n720), .B(new_n1104), .C1(new_n1103), .C2(new_n1102), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n1101), .A2(new_n1105), .B1(G107), .B2(new_n207), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n868), .B(new_n1099), .C1(new_n833), .C2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1107), .A2(KEYINPUT114), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n713), .A2(new_n1014), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1107), .A2(KEYINPUT114), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1040), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1110), .A2(new_n1111), .B1(new_n1112), .B2(new_n828), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1041), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n722), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1112), .A2(new_n781), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1113), .B1(new_n1115), .B2(new_n1116), .ZN(G393));
  NAND2_X1  g0917(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1118), .A2(new_n1042), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n828), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n987), .A2(new_n242), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n833), .B1(new_n523), .B2(new_n207), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n829), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n874), .B1(new_n299), .B2(new_n804), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(G143), .B2(new_n799), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n788), .A2(new_n994), .B1(new_n803), .B2(new_n884), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT51), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n791), .A2(new_n222), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1128), .B(new_n834), .C1(G68), .C2(new_n813), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n810), .A2(new_n340), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1125), .A2(new_n1127), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n883), .A2(new_n591), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n323), .B1(new_n479), .B2(new_n791), .C1(new_n477), .C2(new_n794), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n820), .B1(new_n465), .B2(new_n804), .C1(new_n801), .C2(new_n876), .ZN(new_n1134));
  OR3_X1    g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n789), .A2(G317), .B1(new_n822), .B2(G311), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT52), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1131), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1123), .B1(new_n1138), .B2(new_n786), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n1053), .B2(new_n1014), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n722), .B1(new_n1119), .B2(new_n1041), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1120), .B(new_n1140), .C1(new_n1141), .C2(new_n1142), .ZN(G390));
  AOI21_X1  g0943(.A(new_n772), .B1(new_n774), .B2(new_n775), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n944), .A2(new_n1144), .A3(new_n857), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n773), .A2(new_n778), .A3(new_n857), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n942), .A2(new_n943), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1145), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n940), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n773), .A2(new_n778), .A3(new_n857), .A4(new_n944), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n856), .A2(new_n388), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n742), .A2(new_n704), .A3(new_n1151), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1152), .A2(new_n859), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n863), .B1(new_n1144), .B2(KEYINPUT116), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT116), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n771), .B2(new_n772), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n944), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n1148), .A2(new_n1149), .B1(new_n1154), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n441), .A2(new_n1144), .ZN(new_n1160));
  AND4_X1   g0960(.A1(new_n392), .A2(new_n672), .A3(new_n967), .A4(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT117), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1159), .A2(new_n1161), .A3(KEYINPUT117), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT115), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n956), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n976), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1147), .B1(new_n859), .B2(new_n1152), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n955), .A2(new_n957), .B1(new_n945), .B2(new_n1168), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1167), .B(new_n1145), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n955), .A2(new_n957), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n945), .A2(new_n1168), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1152), .A2(new_n859), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n944), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n956), .B1(new_n935), .B2(new_n975), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1176), .A2(new_n1180), .A3(new_n1150), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1173), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1176), .A2(new_n1180), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1167), .B1(new_n1183), .B2(new_n1145), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1166), .A2(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1174), .A2(new_n1175), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1145), .ZN(new_n1188));
  OAI21_X1  g0988(.A(KEYINPUT115), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1189), .A2(new_n1181), .A3(new_n1173), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1190), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1186), .A2(new_n1191), .A3(new_n722), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1174), .A2(new_n830), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n869), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1194), .A2(new_n340), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n797), .A2(new_n216), .B1(new_n803), .B2(new_n479), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n876), .A2(new_n591), .B1(new_n224), .B2(new_n804), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(new_n810), .C2(G97), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1128), .B1(G283), .B2(new_n789), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1198), .A2(new_n323), .A3(new_n814), .A4(new_n1199), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT118), .Z(new_n1201));
  AOI22_X1  g1001(.A1(new_n799), .A2(G125), .B1(new_n872), .B2(G137), .ZN(new_n1202));
  INV_X1    g1002(.A(G132), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1202), .B1(new_n299), .B2(new_n797), .C1(new_n1203), .C2(new_n803), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n794), .A2(new_n994), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1204), .B1(KEYINPUT53), .B2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n791), .A2(new_n884), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1208), .B(new_n323), .C1(G128), .C2(new_n789), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(KEYINPUT54), .B(G143), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT53), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n810), .A2(new_n1211), .B1(new_n1205), .B2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1207), .A2(new_n1209), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1201), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT119), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n871), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n868), .B(new_n1195), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1193), .A2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n1190), .B2(new_n827), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1192), .A2(new_n1224), .ZN(G378));
  NAND3_X1  g1025(.A1(new_n972), .A2(G330), .A3(new_n977), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n356), .A2(new_n392), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n345), .A2(new_n348), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n700), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1227), .B(new_n1229), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1226), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1234), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1236), .A2(G330), .A3(new_n972), .A4(new_n977), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n966), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n959), .A2(new_n964), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1240), .A2(new_n1237), .A3(new_n1235), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n828), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n868), .B1(new_n869), .B2(new_n299), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(G77), .A2(new_n813), .B1(new_n789), .B2(G116), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1245), .B(new_n834), .C1(new_n216), .C2(new_n791), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n798), .A2(G58), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT120), .ZN(new_n1248));
  INV_X1    g1048(.A(G41), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1249), .B1(new_n224), .B2(new_n803), .C1(new_n876), .C2(new_n477), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1246), .A2(new_n1248), .A3(new_n1250), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n810), .A2(new_n377), .B1(G97), .B2(new_n872), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1252), .A2(KEYINPUT121), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(KEYINPUT121), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1251), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT58), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1258));
  INV_X1    g1058(.A(G128), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n803), .A2(new_n1259), .B1(new_n1203), .B2(new_n804), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(G125), .B2(new_n789), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n813), .A2(new_n1211), .B1(new_n792), .B2(G150), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1261), .B(new_n1262), .C1(new_n883), .C2(new_n882), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1263), .A2(KEYINPUT59), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(KEYINPUT59), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n264), .B(new_n1249), .C1(new_n797), .C2(new_n884), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(G124), .B2(new_n799), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1264), .A2(new_n1265), .A3(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1258), .A2(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1249), .B1(new_n834), .B2(new_n264), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1257), .B(new_n1269), .C1(new_n299), .C2(new_n1270), .ZN(new_n1271));
  OAI221_X1 g1071(.A(new_n1244), .B1(new_n871), .B2(new_n1271), .C1(new_n1236), .C2(new_n831), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1243), .A2(new_n1272), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n1159), .A2(KEYINPUT117), .A3(new_n1161), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT117), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1161), .B1(new_n1276), .B2(new_n1190), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT57), .B1(new_n1277), .B2(new_n1242), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n672), .A2(new_n967), .A3(new_n392), .A4(new_n1160), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(new_n1166), .B2(new_n1185), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1240), .A2(new_n1237), .A3(new_n1235), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n1235), .A2(new_n1237), .B1(new_n960), .B2(new_n965), .ZN(new_n1282));
  OAI21_X1  g1082(.A(KEYINPUT57), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n722), .B1(new_n1280), .B2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1273), .B1(new_n1278), .B2(new_n1284), .ZN(G375));
  OAI22_X1  g1085(.A1(new_n803), .A2(new_n882), .B1(new_n1210), .B2(new_n804), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n813), .A2(G159), .B1(new_n792), .B2(G50), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1287), .B(new_n835), .C1(new_n1259), .C2(new_n876), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n1288), .B(new_n1248), .C1(G150), .C2(new_n810), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1289), .B(KEYINPUT122), .ZN(new_n1290));
  AOI211_X1 g1090(.A(new_n1286), .B(new_n1290), .C1(G132), .C2(new_n789), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(new_n822), .A2(G283), .B1(G116), .B2(new_n872), .ZN(new_n1292));
  OAI221_X1 g1092(.A(new_n1292), .B1(new_n222), .B2(new_n797), .C1(new_n465), .C2(new_n876), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(G97), .A2(new_n813), .B1(new_n789), .B2(G294), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1294), .B(new_n323), .C1(new_n376), .C2(new_n791), .ZN(new_n1295));
  AOI211_X1 g1095(.A(new_n1293), .B(new_n1295), .C1(G107), .C2(new_n810), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n786), .B1(new_n1291), .B2(new_n1296), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1297), .B(new_n829), .C1(G68), .C2(new_n1194), .ZN(new_n1298));
  XOR2_X1   g1098(.A(new_n1298), .B(KEYINPUT123), .Z(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(new_n831), .B2(new_n944), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1159), .A2(new_n828), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT124), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1300), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1302), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  OAI221_X1 g1106(.A(new_n1279), .B1(new_n1158), .B2(new_n1154), .C1(new_n1149), .C2(new_n1148), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1276), .A2(new_n1047), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1306), .A2(new_n1308), .ZN(G381));
  INV_X1    g1109(.A(G390), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1310), .A2(new_n1306), .A3(new_n1308), .A4(new_n1311), .ZN(new_n1312));
  OR4_X1    g1112(.A1(G387), .A2(G375), .A3(G378), .A4(new_n1312), .ZN(G407));
  INV_X1    g1113(.A(new_n722), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1314), .B1(new_n1276), .B2(new_n1190), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1223), .B1(new_n1315), .B2(new_n1186), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n702), .A2(G213), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1319));
  OAI211_X1 g1119(.A(G407), .B(G213), .C1(G375), .C2(new_n1319), .ZN(G409));
  OAI211_X1 g1120(.A(G378), .B(new_n1273), .C1(new_n1278), .C2(new_n1284), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1277), .A2(new_n1047), .A3(new_n1242), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1243), .A2(new_n1272), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1316), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1321), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1317), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1318), .A2(G2897), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT60), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n722), .B1(new_n1307), .B2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1330), .ZN(new_n1331));
  NOR3_X1   g1131(.A1(new_n1274), .A2(new_n1275), .A3(new_n1329), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1307), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1331), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(G384), .B1(new_n1334), .B2(new_n1306), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1164), .A2(KEYINPUT60), .A3(new_n1165), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1330), .B1(new_n1336), .B2(new_n1307), .ZN(new_n1337));
  INV_X1    g1137(.A(G384), .ZN(new_n1338));
  NOR3_X1   g1138(.A1(new_n1337), .A2(new_n1338), .A3(new_n1305), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1328), .B1(new_n1335), .B2(new_n1339), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1334), .A2(new_n1306), .A3(G384), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1338), .B1(new_n1337), .B2(new_n1305), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1341), .A2(new_n1342), .A3(new_n1327), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1340), .A2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(KEYINPUT61), .B1(new_n1326), .B2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1347));
  AOI211_X1 g1147(.A(new_n1318), .B(new_n1347), .C1(new_n1321), .C2(new_n1324), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT62), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1347), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1325), .A2(new_n1317), .A3(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1352), .A2(KEYINPUT62), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1346), .A2(new_n1350), .A3(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(G387), .A2(new_n1310), .ZN(new_n1355));
  XNOR2_X1  g1155(.A(G393), .B(new_n849), .ZN(new_n1356));
  OAI211_X1 g1156(.A(G390), .B(new_n1015), .C1(new_n1048), .C2(new_n1075), .ZN(new_n1357));
  AND3_X1   g1157(.A1(new_n1355), .A2(new_n1356), .A3(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1356), .B1(new_n1355), .B2(new_n1357), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1358), .A2(new_n1359), .ZN(new_n1360));
  INV_X1    g1160(.A(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1354), .A2(new_n1361), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT63), .ZN(new_n1363));
  NOR2_X1   g1163(.A1(new_n1347), .A2(new_n1363), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1325), .A2(new_n1317), .A3(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(KEYINPUT126), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1365), .A2(new_n1366), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1318), .B1(new_n1321), .B2(new_n1324), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(new_n1368), .A2(KEYINPUT126), .A3(new_n1364), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1367), .A2(new_n1369), .ZN(new_n1370));
  INV_X1    g1170(.A(KEYINPUT61), .ZN(new_n1371));
  OAI211_X1 g1171(.A(new_n1360), .B(new_n1371), .C1(new_n1368), .C2(new_n1344), .ZN(new_n1372));
  INV_X1    g1172(.A(new_n1372), .ZN(new_n1373));
  INV_X1    g1173(.A(KEYINPUT125), .ZN(new_n1374));
  OAI21_X1  g1174(.A(new_n1374), .B1(new_n1348), .B2(KEYINPUT63), .ZN(new_n1375));
  NAND3_X1  g1175(.A1(new_n1352), .A2(KEYINPUT125), .A3(new_n1363), .ZN(new_n1376));
  NAND4_X1  g1176(.A1(new_n1370), .A2(new_n1373), .A3(new_n1375), .A4(new_n1376), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1362), .A2(new_n1377), .ZN(G405));
  OR2_X1    g1178(.A1(new_n1361), .A2(KEYINPUT127), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(G375), .A2(new_n1316), .ZN(new_n1380));
  INV_X1    g1180(.A(new_n1380), .ZN(new_n1381));
  INV_X1    g1181(.A(new_n1321), .ZN(new_n1382));
  NOR3_X1   g1182(.A1(new_n1381), .A2(new_n1382), .A3(new_n1351), .ZN(new_n1383));
  INV_X1    g1183(.A(new_n1383), .ZN(new_n1384));
  AOI21_X1  g1184(.A(new_n1347), .B1(new_n1380), .B2(new_n1321), .ZN(new_n1385));
  INV_X1    g1185(.A(new_n1385), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1361), .A2(KEYINPUT127), .ZN(new_n1387));
  NAND4_X1  g1187(.A1(new_n1379), .A2(new_n1384), .A3(new_n1386), .A4(new_n1387), .ZN(new_n1388));
  OAI211_X1 g1188(.A(KEYINPUT127), .B(new_n1361), .C1(new_n1383), .C2(new_n1385), .ZN(new_n1389));
  NAND2_X1  g1189(.A1(new_n1388), .A2(new_n1389), .ZN(G402));
endmodule


