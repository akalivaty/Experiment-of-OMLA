//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n808, new_n810, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n202));
  AND2_X1   g001(.A1(G211gat), .A2(G218gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G211gat), .A2(G218gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n206), .B(new_n207), .C1(KEYINPUT22), .C2(new_n203), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(KEYINPUT22), .B2(new_n203), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(new_n205), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT29), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(KEYINPUT3), .ZN(new_n212));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  INV_X1    g012(.A(G155gat), .ZN(new_n214));
  INV_X1    g013(.A(G162gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G141gat), .B(G148gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n213), .B(new_n216), .C1(new_n217), .C2(KEYINPUT2), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n213), .A2(KEYINPUT2), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT79), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n216), .A2(new_n213), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT79), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n213), .A2(new_n222), .A3(KEYINPUT2), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n220), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT78), .ZN(new_n225));
  INV_X1    g024(.A(G148gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(G141gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(G141gat), .ZN(new_n228));
  INV_X1    g027(.A(G141gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(KEYINPUT78), .A3(G148gat), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n227), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n218), .B1(new_n224), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n202), .B1(new_n212), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n208), .A2(new_n210), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n232), .A2(KEYINPUT3), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n236), .B1(new_n237), .B2(KEYINPUT29), .ZN(new_n238));
  OAI211_X1 g037(.A(KEYINPUT83), .B(new_n232), .C1(new_n211), .C2(KEYINPUT3), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n234), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(G228gat), .A3(G233gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(G228gat), .A2(G233gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n227), .A2(new_n228), .A3(new_n230), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n243), .A2(new_n221), .A3(new_n223), .A4(new_n220), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT80), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n244), .A2(new_n245), .A3(new_n218), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n245), .B1(new_n244), .B2(new_n218), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n238), .B(new_n242), .C1(new_n248), .C2(new_n212), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n241), .A2(G22gat), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(G22gat), .B1(new_n241), .B2(new_n249), .ZN(new_n251));
  XNOR2_X1  g050(.A(G78gat), .B(G106gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT31), .B(G50gat), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n252), .B(new_n253), .Z(new_n254));
  OAI22_X1  g053(.A1(new_n250), .A2(new_n251), .B1(KEYINPUT84), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n241), .A2(new_n249), .ZN(new_n256));
  INV_X1    g055(.A(G22gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n254), .B(KEYINPUT84), .Z(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n241), .A2(G22gat), .A3(new_n249), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT28), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT27), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G183gat), .ZN(new_n266));
  INV_X1    g065(.A(G183gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT27), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT70), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT70), .B1(new_n267), .B2(KEYINPUT27), .ZN(new_n270));
  INV_X1    g069(.A(G190gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n264), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n267), .A2(KEYINPUT27), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n265), .A2(G183gat), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n266), .A2(new_n268), .A3(KEYINPUT71), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n264), .A2(G190gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT26), .ZN(new_n282));
  INV_X1    g081(.A(G169gat), .ZN(new_n283));
  INV_X1    g082(.A(G176gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n286));
  AND3_X1   g085(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n285), .B(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT72), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n289), .A2(new_n293), .A3(new_n290), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n281), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  AND2_X1   g094(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n296));
  NOR2_X1   g095(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n290), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT69), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT69), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n303), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n298), .A2(new_n300), .A3(new_n302), .A4(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT23), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(new_n287), .B2(new_n288), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT67), .ZN(new_n308));
  AND2_X1   g107(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n309));
  NOR2_X1   g108(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n310));
  OAI22_X1  g109(.A1(new_n309), .A2(new_n310), .B1(G169gat), .B2(G176gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT67), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n306), .B(new_n312), .C1(new_n287), .C2(new_n288), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n305), .A2(new_n308), .A3(new_n311), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT25), .ZN(new_n315));
  NAND2_X1  g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT65), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n311), .A2(new_n320), .A3(new_n306), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT66), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT66), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n311), .A2(new_n320), .A3(new_n323), .A4(new_n306), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT24), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n290), .B1(new_n299), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT25), .B1(new_n326), .B2(new_n301), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n322), .A2(new_n324), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n295), .A2(new_n315), .A3(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G127gat), .B(G134gat), .ZN(new_n330));
  XOR2_X1   g129(.A(G113gat), .B(G120gat), .Z(new_n331));
  INV_X1    g130(.A(KEYINPUT1), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G120gat), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT74), .B1(new_n334), .B2(G113gat), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n336));
  INV_X1    g135(.A(G113gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n337), .A3(G120gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n334), .A2(KEYINPUT73), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT73), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G120gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n335), .B(new_n338), .C1(new_n342), .C2(new_n337), .ZN(new_n343));
  OR2_X1    g142(.A1(KEYINPUT75), .A2(KEYINPUT1), .ZN(new_n344));
  NAND2_X1  g143(.A1(KEYINPUT75), .A2(KEYINPUT1), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n330), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n333), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n329), .A2(new_n348), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n324), .A2(new_n327), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n322), .A2(new_n350), .B1(new_n314), .B2(KEYINPUT25), .ZN(new_n351));
  INV_X1    g150(.A(new_n330), .ZN(new_n352));
  XNOR2_X1  g151(.A(G113gat), .B(G120gat), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n352), .B1(KEYINPUT1), .B2(new_n353), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n339), .A2(new_n341), .A3(G113gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n335), .A2(new_n338), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n354), .B1(new_n357), .B2(new_n346), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n351), .A2(new_n358), .A3(new_n295), .ZN(new_n359));
  INV_X1    g158(.A(G227gat), .ZN(new_n360));
  INV_X1    g159(.A(G233gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n349), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT32), .ZN(new_n364));
  XOR2_X1   g163(.A(G15gat), .B(G43gat), .Z(new_n365));
  XNOR2_X1  g164(.A(G71gat), .B(G99gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT33), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n368), .B1(new_n363), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n362), .B1(new_n349), .B2(new_n359), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT34), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI211_X1 g172(.A(KEYINPUT34), .B(new_n362), .C1(new_n349), .C2(new_n359), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n370), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n370), .A2(new_n373), .A3(new_n374), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n364), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OR3_X1    g177(.A1(new_n370), .A2(new_n373), .A3(new_n374), .ZN(new_n379));
  INV_X1    g178(.A(new_n364), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(new_n380), .A3(new_n375), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT35), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n263), .A2(new_n378), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G8gat), .B(G36gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(G64gat), .B(G92gat), .ZN(new_n385));
  XOR2_X1   g184(.A(new_n384), .B(new_n385), .Z(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n389), .A2(KEYINPUT29), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n390), .B1(new_n351), .B2(new_n295), .ZN(new_n391));
  AND4_X1   g190(.A1(new_n295), .A2(new_n315), .A3(new_n328), .A4(new_n388), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n236), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n393), .A2(KEYINPUT76), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT76), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n395), .B(new_n236), .C1(new_n391), .C2(new_n392), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n329), .B1(KEYINPUT29), .B2(new_n389), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n351), .A2(new_n295), .A3(new_n388), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n235), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n387), .B1(new_n394), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n393), .A2(KEYINPUT76), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n402), .A2(new_n386), .A3(new_n396), .A4(new_n399), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n401), .A2(KEYINPUT77), .A3(KEYINPUT30), .A4(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT77), .B(KEYINPUT30), .ZN(new_n405));
  OR2_X1    g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT85), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n404), .A2(KEYINPUT85), .A3(new_n406), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n383), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G1gat), .B(G29gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT0), .ZN(new_n412));
  XNOR2_X1  g211(.A(G57gat), .B(G85gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT5), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n233), .A2(new_n348), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n358), .A2(new_n232), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n416), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n232), .A2(KEYINPUT80), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n244), .A2(new_n245), .A3(new_n218), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n348), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT81), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n425), .A2(new_n426), .A3(KEYINPUT4), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n426), .B1(new_n425), .B2(KEYINPUT4), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n417), .A2(KEYINPUT4), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n348), .B1(KEYINPUT3), .B2(new_n232), .ZN(new_n431));
  INV_X1    g230(.A(new_n237), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n420), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n422), .B1(new_n430), .B2(new_n434), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n246), .A2(new_n247), .A3(new_n358), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n417), .A2(KEYINPUT4), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n421), .B1(new_n431), .B2(new_n432), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n416), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n415), .B1(new_n435), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT6), .ZN(new_n444));
  INV_X1    g243(.A(new_n422), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT81), .B1(new_n436), .B2(new_n437), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n425), .A2(new_n426), .A3(KEYINPUT4), .ZN(new_n447));
  INV_X1    g246(.A(new_n429), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n445), .B1(new_n449), .B2(new_n441), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n441), .A2(new_n416), .ZN(new_n451));
  INV_X1    g250(.A(new_n417), .ZN(new_n452));
  MUX2_X1   g251(.A(new_n425), .B(new_n452), .S(KEYINPUT4), .Z(new_n453));
  OAI21_X1  g252(.A(new_n415), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n444), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT87), .B1(new_n443), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n443), .A2(KEYINPUT82), .A3(KEYINPUT6), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT82), .ZN(new_n458));
  INV_X1    g257(.A(new_n442), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n414), .B1(new_n450), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n458), .B1(new_n460), .B2(new_n444), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT87), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n425), .A2(KEYINPUT4), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n429), .B1(new_n463), .B2(KEYINPUT81), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n434), .B1(new_n464), .B2(new_n447), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n442), .B(new_n415), .C1(new_n465), .C2(new_n445), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n460), .A2(new_n462), .A3(new_n444), .A4(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n456), .A2(new_n457), .A3(new_n461), .A4(new_n467), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n381), .A2(new_n378), .ZN(new_n469));
  INV_X1    g268(.A(new_n451), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n414), .B1(new_n470), .B2(new_n440), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT6), .B1(new_n435), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n460), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n461), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n404), .A2(new_n406), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n469), .A2(new_n474), .A3(new_n263), .A4(new_n475), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n410), .A2(new_n468), .B1(new_n476), .B2(KEYINPUT35), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n399), .A2(new_n393), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT38), .B1(new_n478), .B2(KEYINPUT37), .ZN(new_n479));
  XNOR2_X1  g278(.A(KEYINPUT88), .B(KEYINPUT37), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n402), .A2(new_n396), .A3(new_n399), .A4(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n481), .A3(new_n387), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT89), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n479), .A2(new_n481), .A3(KEYINPUT89), .A4(new_n387), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n484), .A2(new_n485), .A3(new_n403), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n443), .A2(new_n455), .A3(KEYINPUT87), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n462), .B1(new_n472), .B2(new_n460), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n457), .A2(new_n461), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n486), .A2(KEYINPUT90), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT90), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n484), .A2(new_n485), .A3(new_n403), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n492), .B1(new_n468), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT37), .B1(new_n394), .B2(new_n400), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n495), .A2(new_n387), .A3(new_n481), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT38), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT91), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n491), .A2(new_n494), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n263), .ZN(new_n501));
  INV_X1    g300(.A(new_n409), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n502), .A2(new_n407), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n440), .A2(new_n433), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT39), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n505), .A3(new_n421), .ZN(new_n506));
  INV_X1    g305(.A(new_n419), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n505), .B1(new_n507), .B2(new_n420), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n438), .A2(new_n439), .B1(new_n432), .B2(new_n431), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n508), .B1(new_n509), .B2(new_n420), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n506), .A2(new_n510), .A3(KEYINPUT40), .A4(new_n415), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT86), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n510), .A2(new_n415), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT40), .B1(new_n513), .B2(new_n506), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n512), .A2(new_n443), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n501), .B1(new_n503), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n381), .A2(new_n378), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT36), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n474), .A2(new_n475), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n501), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n477), .B1(new_n517), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT98), .ZN(new_n526));
  XNOR2_X1  g325(.A(G113gat), .B(G141gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G169gat), .B(G197gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n531), .B(KEYINPUT12), .Z(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534));
  XOR2_X1   g333(.A(new_n534), .B(KEYINPUT97), .Z(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G15gat), .B(G22gat), .ZN(new_n537));
  INV_X1    g336(.A(G1gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT16), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(G1gat), .B2(new_n537), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n541), .A2(G8gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(G8gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT17), .ZN(new_n545));
  XNOR2_X1  g344(.A(G43gat), .B(G50gat), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n546), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n547));
  XOR2_X1   g346(.A(G43gat), .B(G50gat), .Z(new_n548));
  INV_X1    g347(.A(KEYINPUT15), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT93), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT93), .ZN(new_n551));
  NOR3_X1   g350(.A1(new_n546), .A2(new_n551), .A3(KEYINPUT15), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n547), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT14), .ZN(new_n556));
  INV_X1    g355(.A(G29gat), .ZN(new_n557));
  INV_X1    g356(.A(G36gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT94), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n556), .A2(new_n557), .A3(new_n558), .A4(KEYINPUT94), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n555), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OR2_X1    g362(.A1(new_n563), .A2(KEYINPUT95), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT95), .ZN(new_n565));
  AOI211_X1 g364(.A(new_n565), .B(new_n555), .C1(new_n561), .C2(new_n562), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n553), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(G43gat), .ZN(new_n569));
  INV_X1    g368(.A(G50gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(G43gat), .A2(G50gat), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT15), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n559), .A2(new_n554), .ZN(new_n574));
  NAND2_X1  g373(.A1(G29gat), .A2(G36gat), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n545), .B1(new_n568), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n544), .B1(new_n577), .B2(KEYINPUT96), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT96), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n579), .B1(new_n542), .B2(new_n543), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n580), .A2(KEYINPUT17), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n573), .A2(new_n575), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n551), .B1(new_n546), .B2(KEYINPUT15), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n548), .A2(KEYINPUT93), .A3(new_n549), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n563), .A2(KEYINPUT95), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n585), .B1(new_n586), .B2(new_n566), .ZN(new_n587));
  INV_X1    g386(.A(new_n576), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n581), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n536), .B1(new_n578), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT18), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n564), .A2(new_n567), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n576), .B1(new_n593), .B2(new_n585), .ZN(new_n594));
  INV_X1    g393(.A(new_n544), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n589), .A2(new_n544), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n535), .B(KEYINPUT13), .Z(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n591), .A2(new_n592), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT17), .B1(new_n587), .B2(new_n588), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n595), .B1(new_n602), .B2(new_n579), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n594), .B1(new_n580), .B2(KEYINPUT17), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n535), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT18), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n533), .B1(new_n601), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n600), .B1(new_n596), .B2(new_n597), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n608), .B1(new_n605), .B2(KEYINPUT18), .ZN(new_n609));
  AOI211_X1 g408(.A(new_n592), .B(new_n535), .C1(new_n603), .C2(new_n604), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n609), .A2(new_n610), .A3(new_n532), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n526), .B1(new_n607), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n532), .B1(new_n609), .B2(new_n610), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n591), .A2(new_n592), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n614), .A2(new_n606), .A3(new_n608), .A4(new_n533), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n613), .A2(new_n615), .A3(KEYINPUT98), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n618));
  AND2_X1   g417(.A1(G57gat), .A2(G64gat), .ZN(new_n619));
  NOR2_X1   g418(.A1(G57gat), .A2(G64gat), .ZN(new_n620));
  NOR3_X1   g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(G71gat), .ZN(new_n622));
  INV_X1    g421(.A(G78gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G71gat), .A2(G78gat), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT9), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n624), .B(new_n625), .C1(KEYINPUT99), .C2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n621), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n621), .A2(new_n627), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n631), .A2(KEYINPUT21), .ZN(new_n632));
  AND2_X1   g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(G127gat), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n544), .B1(KEYINPUT21), .B2(new_n631), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n635), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(new_n214), .ZN(new_n640));
  XNOR2_X1  g439(.A(G183gat), .B(G211gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n640), .B(new_n641), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n638), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G190gat), .B(G218gat), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT100), .ZN(new_n647));
  INV_X1    g446(.A(G85gat), .ZN(new_n648));
  INV_X1    g447(.A(G92gat), .ZN(new_n649));
  OAI21_X1  g448(.A(KEYINPUT7), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT7), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(G85gat), .A3(G92gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G99gat), .B(G106gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(G99gat), .A2(G106gat), .ZN(new_n655));
  AOI22_X1  g454(.A1(KEYINPUT8), .A2(new_n655), .B1(new_n648), .B2(new_n649), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n654), .B1(new_n653), .B2(new_n656), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n659), .A2(KEYINPUT17), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT41), .ZN(new_n661));
  NAND2_X1  g460(.A1(G232gat), .A2(G233gat), .ZN(new_n662));
  OAI22_X1  g461(.A1(new_n594), .A2(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n589), .A2(KEYINPUT17), .A3(new_n659), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n647), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G134gat), .B(G162gat), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n646), .A2(KEYINPUT100), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n662), .A2(new_n661), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n666), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n647), .B(new_n671), .C1(new_n663), .C2(new_n664), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n667), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n670), .B1(new_n667), .B2(new_n672), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  OAI22_X1  g476(.A1(new_n629), .A2(new_n630), .B1(new_n657), .B2(new_n658), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n653), .A2(new_n656), .ZN(new_n679));
  INV_X1    g478(.A(new_n654), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n624), .A2(new_n625), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n626), .A2(KEYINPUT99), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n619), .A2(new_n620), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n682), .B(new_n683), .C1(new_n684), .C2(new_n618), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n681), .A2(new_n685), .A3(new_n628), .A4(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n678), .A2(KEYINPUT101), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT101), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n631), .A2(new_n659), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT10), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT102), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n687), .A2(new_n692), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(G230gat), .A2(G233gat), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT10), .B1(new_n688), .B2(new_n690), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT102), .B1(new_n699), .B2(new_n695), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(G120gat), .B(G148gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(G176gat), .B(G204gat), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n702), .B(new_n703), .Z(new_n704));
  OAI211_X1 g503(.A(new_n701), .B(new_n704), .C1(new_n698), .C2(new_n691), .ZN(new_n705));
  INV_X1    g504(.A(new_n704), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n699), .A2(new_n695), .ZN(new_n707));
  INV_X1    g506(.A(new_n698), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n691), .A2(new_n698), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n706), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n705), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n644), .A2(new_n677), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n525), .A2(new_n617), .A3(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n474), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(new_n538), .ZN(G1324gat));
  INV_X1    g517(.A(new_n503), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT42), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n720), .A2(new_n721), .A3(G8gat), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT16), .B(G8gat), .Z(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT103), .ZN(new_n724));
  NOR2_X1   g523(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n724), .B(new_n725), .Z(new_n726));
  AOI21_X1  g525(.A(new_n722), .B1(new_n720), .B2(new_n726), .ZN(G1325gat));
  OAI21_X1  g526(.A(G15gat), .B1(new_n716), .B2(new_n520), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n518), .A2(G15gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n716), .B2(new_n729), .ZN(G1326gat));
  OR3_X1    g529(.A1(new_n716), .A2(KEYINPUT105), .A3(new_n263), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT105), .B1(new_n716), .B2(new_n263), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(KEYINPUT43), .B(G22gat), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n733), .B(new_n734), .Z(G1327gat));
  XNOR2_X1  g534(.A(new_n638), .B(new_n642), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n713), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(new_n677), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT106), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n525), .A2(new_n617), .A3(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n474), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n741), .A2(new_n557), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(KEYINPUT44), .B1(new_n524), .B2(new_n677), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(new_n674), .B2(new_n675), .ZN(new_n748));
  INV_X1    g547(.A(new_n675), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n749), .A2(KEYINPUT108), .A3(new_n673), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(KEYINPUT44), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT109), .B1(new_n524), .B2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n520), .A2(new_n522), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n757), .B1(new_n500), .B2(new_n516), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n756), .B(new_n753), .C1(new_n758), .C2(new_n477), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n746), .A2(new_n755), .A3(new_n759), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n613), .A2(KEYINPUT107), .A3(new_n615), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT107), .B1(new_n613), .B2(new_n615), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n737), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(G29gat), .B1(new_n765), .B2(new_n474), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT110), .B1(new_n745), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n743), .B(KEYINPUT45), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n769), .A2(new_n770), .A3(new_n766), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n771), .ZN(G1328gat));
  NOR3_X1   g571(.A1(new_n740), .A2(G36gat), .A3(new_n719), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT46), .ZN(new_n774));
  OAI21_X1  g573(.A(G36gat), .B1(new_n765), .B2(new_n719), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(G1329gat));
  INV_X1    g575(.A(new_n520), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n760), .A2(G43gat), .A3(new_n777), .A4(new_n764), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n569), .B1(new_n740), .B2(new_n518), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g580(.A1(new_n760), .A2(new_n501), .A3(new_n764), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n760), .A2(KEYINPUT112), .A3(new_n501), .A4(new_n764), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n784), .A2(G50gat), .A3(new_n785), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n740), .A2(G50gat), .A3(new_n263), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(KEYINPUT48), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n782), .A2(G50gat), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n788), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT48), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n787), .B1(new_n782), .B2(G50gat), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n795), .A2(KEYINPUT111), .A3(KEYINPUT48), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n789), .B1(new_n794), .B2(new_n796), .ZN(G1331gat));
  NAND2_X1  g596(.A1(new_n763), .A2(new_n712), .ZN(new_n798));
  NOR4_X1   g597(.A1(new_n524), .A2(new_n736), .A3(new_n676), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n742), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n503), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n803));
  XOR2_X1   g602(.A(KEYINPUT49), .B(G64gat), .Z(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n802), .B2(new_n804), .ZN(G1333gat));
  AOI21_X1  g604(.A(new_n622), .B1(new_n799), .B2(new_n777), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n518), .A2(G71gat), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n806), .B1(new_n799), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g608(.A1(new_n799), .A2(new_n501), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(G78gat), .ZN(G1335gat));
  INV_X1    g610(.A(new_n763), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(new_n644), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n525), .A2(KEYINPUT51), .A3(new_n676), .A4(new_n813), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n676), .B(new_n813), .C1(new_n758), .C2(new_n477), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(KEYINPUT113), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n818), .A2(KEYINPUT113), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n819), .A2(new_n820), .A3(new_n713), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n648), .A3(new_n742), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n798), .A2(new_n644), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n760), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(G85gat), .B1(new_n824), .B2(new_n474), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n822), .A2(new_n825), .ZN(G1336gat));
  OAI21_X1  g625(.A(G92gat), .B1(new_n824), .B2(new_n719), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n719), .A2(G92gat), .A3(new_n713), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT114), .B1(new_n818), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT52), .ZN(G1337gat));
  INV_X1    g630(.A(G99gat), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n821), .A2(new_n832), .A3(new_n469), .ZN(new_n833));
  OAI21_X1  g632(.A(G99gat), .B1(new_n824), .B2(new_n520), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(G1338gat));
  OAI21_X1  g634(.A(G106gat), .B1(new_n824), .B2(new_n263), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(KEYINPUT115), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n263), .A2(new_n713), .A3(G106gat), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n818), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n818), .A2(KEYINPUT116), .A3(new_n838), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT53), .B1(new_n837), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT115), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT53), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n836), .B(new_n846), .C1(KEYINPUT53), .C2(new_n839), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n844), .A2(new_n847), .ZN(G1339gat));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n849), .B(new_n698), .C1(new_n699), .C2(new_n695), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n706), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n849), .B1(new_n707), .B2(new_n708), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n701), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n705), .B1(new_n853), .B2(KEYINPUT55), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT55), .ZN(new_n855));
  AOI211_X1 g654(.A(new_n855), .B(new_n851), .C1(new_n701), .C2(new_n852), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n857), .B1(new_n761), .B2(new_n762), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n603), .A2(new_n535), .A3(new_n604), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n598), .B2(new_n600), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n531), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n712), .A2(new_n615), .A3(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n751), .B1(new_n858), .B2(new_n863), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n615), .A2(new_n861), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n751), .A2(new_n865), .A3(new_n857), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n736), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n715), .A2(new_n763), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n474), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n870), .A2(new_n263), .A3(new_n469), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n719), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n337), .A3(new_n812), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n501), .B1(new_n868), .B2(new_n869), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n875), .B(new_n876), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n503), .A2(new_n474), .A3(new_n518), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n617), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n881), .A2(KEYINPUT118), .A3(G113gat), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT118), .B1(new_n881), .B2(G113gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n874), .B1(new_n882), .B2(new_n883), .ZN(G1340gat));
  OAI21_X1  g683(.A(G120gat), .B1(new_n879), .B2(new_n713), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n712), .A2(new_n339), .A3(new_n341), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(new_n872), .B2(new_n886), .ZN(G1341gat));
  AOI21_X1  g686(.A(KEYINPUT119), .B1(new_n873), .B2(new_n644), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(G127gat), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n873), .A2(KEYINPUT119), .A3(new_n644), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n644), .A2(G127gat), .ZN(new_n891));
  AOI22_X1  g690(.A1(new_n889), .A2(new_n890), .B1(new_n880), .B2(new_n891), .ZN(G1342gat));
  INV_X1    g691(.A(G134gat), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n503), .A2(new_n677), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT120), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n871), .A2(new_n893), .A3(new_n896), .ZN(new_n897));
  XOR2_X1   g696(.A(new_n897), .B(KEYINPUT56), .Z(new_n898));
  OAI21_X1  g697(.A(G134gat), .B1(new_n879), .B2(new_n677), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1343gat));
  NOR2_X1   g699(.A1(new_n777), .A2(new_n474), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n719), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n868), .A2(new_n869), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(new_n263), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n617), .A2(new_n857), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n677), .B1(new_n906), .B2(new_n862), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n644), .B1(new_n907), .B2(new_n866), .ZN(new_n908));
  INV_X1    g707(.A(new_n869), .ZN(new_n909));
  OAI211_X1 g708(.A(KEYINPUT57), .B(new_n501), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n902), .B1(new_n905), .B2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(G141gat), .B1(new_n912), .B2(new_n763), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n870), .A2(new_n501), .A3(new_n520), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n914), .A2(new_n229), .A3(new_n719), .A4(new_n617), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT58), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n229), .B1(new_n911), .B2(new_n617), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n916), .A2(new_n917), .B1(new_n918), .B2(new_n919), .ZN(G1344gat));
  NAND4_X1  g719(.A1(new_n914), .A2(new_n226), .A3(new_n719), .A4(new_n712), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT121), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n923));
  INV_X1    g722(.A(new_n902), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n714), .A2(new_n617), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n857), .A2(new_n676), .A3(new_n865), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n862), .B1(new_n617), .B2(new_n857), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n927), .B2(new_n676), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n925), .B1(new_n928), .B2(new_n736), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n903), .B1(new_n929), .B2(new_n263), .ZN(new_n930));
  AOI211_X1 g729(.A(new_n903), .B(new_n263), .C1(new_n868), .C2(new_n869), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n931), .B2(KEYINPUT122), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n263), .B1(new_n868), .B2(new_n869), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n933), .A2(KEYINPUT122), .A3(KEYINPUT57), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n712), .B(new_n924), .C1(new_n932), .C2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n923), .B1(new_n935), .B2(G148gat), .ZN(new_n936));
  AOI211_X1 g735(.A(KEYINPUT59), .B(new_n226), .C1(new_n911), .C2(new_n712), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n922), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n922), .B(KEYINPUT123), .C1(new_n936), .C2(new_n937), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1345gat));
  OAI21_X1  g741(.A(G155gat), .B1(new_n912), .B2(new_n736), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n914), .A2(new_n214), .A3(new_n719), .A4(new_n644), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1346gat));
  OAI21_X1  g744(.A(G162gat), .B1(new_n912), .B2(new_n752), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n914), .A2(new_n215), .A3(new_n896), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1347gat));
  NAND2_X1  g747(.A1(new_n503), .A2(new_n474), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n949), .A2(new_n518), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n875), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(G169gat), .B1(new_n952), .B2(new_n812), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n877), .A2(new_n950), .ZN(new_n954));
  INV_X1    g753(.A(new_n617), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n955), .A2(new_n283), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n953), .B1(new_n954), .B2(new_n956), .ZN(G1348gat));
  AOI21_X1  g756(.A(new_n284), .B1(new_n954), .B2(new_n712), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT124), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n951), .A2(G176gat), .A3(new_n713), .ZN(new_n960));
  OR3_X1    g759(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n959), .B1(new_n958), .B2(new_n960), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1349gat));
  AND4_X1   g762(.A1(new_n277), .A2(new_n952), .A3(new_n278), .A4(new_n644), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n954), .A2(new_n644), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(G183gat), .ZN(new_n966));
  NAND2_X1  g765(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n966), .B(new_n967), .ZN(G1350gat));
  NAND3_X1  g767(.A1(new_n952), .A2(new_n271), .A3(new_n751), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n676), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n970), .B1(new_n971), .B2(G190gat), .ZN(new_n972));
  AOI211_X1 g771(.A(KEYINPUT61), .B(new_n271), .C1(new_n954), .C2(new_n676), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n969), .B1(new_n972), .B2(new_n973), .ZN(G1351gat));
  NOR2_X1   g773(.A1(new_n777), .A2(new_n949), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n933), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT126), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n977), .A2(G197gat), .A3(new_n763), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n978), .B(KEYINPUT127), .ZN(new_n979));
  OR2_X1    g778(.A1(new_n932), .A2(new_n934), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(new_n975), .ZN(new_n981));
  OAI21_X1  g780(.A(G197gat), .B1(new_n981), .B2(new_n955), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n979), .A2(new_n982), .ZN(G1352gat));
  NAND3_X1  g782(.A1(new_n980), .A2(new_n712), .A3(new_n975), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(G204gat), .ZN(new_n985));
  NOR3_X1   g784(.A1(new_n976), .A2(G204gat), .A3(new_n713), .ZN(new_n986));
  XNOR2_X1  g785(.A(new_n986), .B(KEYINPUT62), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n985), .A2(new_n987), .ZN(G1353gat));
  OR3_X1    g787(.A1(new_n977), .A2(G211gat), .A3(new_n736), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n980), .A2(new_n644), .A3(new_n975), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n990), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n991));
  AOI21_X1  g790(.A(KEYINPUT63), .B1(new_n990), .B2(G211gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(G1354gat));
  OAI21_X1  g792(.A(G218gat), .B1(new_n981), .B2(new_n677), .ZN(new_n994));
  OR2_X1    g793(.A1(new_n752), .A2(G218gat), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n994), .B1(new_n977), .B2(new_n995), .ZN(G1355gat));
endmodule


