

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U552 ( .A1(n562), .A2(G2104), .ZN(n914) );
  NOR2_X1 U553 ( .A1(G2104), .A2(n562), .ZN(n921) );
  XOR2_X1 U554 ( .A(n681), .B(n680), .Z(n520) );
  NAND2_X1 U555 ( .A1(n548), .A2(n550), .ZN(n694) );
  XNOR2_X1 U556 ( .A(n572), .B(n571), .ZN(G160) );
  AND2_X1 U557 ( .A1(n544), .A2(n525), .ZN(n543) );
  NOR2_X1 U558 ( .A1(n549), .A2(n554), .ZN(n640) );
  NAND2_X1 U559 ( .A1(n550), .A2(G2072), .ZN(n549) );
  XNOR2_X1 U560 ( .A(KEYINPUT96), .B(KEYINPUT29), .ZN(n680) );
  NAND2_X1 U561 ( .A1(n543), .A2(n524), .ZN(n539) );
  XNOR2_X1 U562 ( .A(n559), .B(KEYINPUT23), .ZN(n561) );
  XNOR2_X1 U563 ( .A(n643), .B(KEYINPUT95), .ZN(n675) );
  OR2_X1 U564 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U565 ( .A1(n675), .A2(n831), .ZN(n645) );
  NOR2_X1 U566 ( .A1(G1966), .A2(n724), .ZN(n704) );
  NOR2_X1 U567 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U568 ( .A1(n520), .A2(n521), .ZN(n535) );
  XNOR2_X1 U569 ( .A(KEYINPUT98), .B(KEYINPUT32), .ZN(n701) );
  NAND2_X1 U570 ( .A1(n557), .A2(n555), .ZN(n554) );
  NAND2_X1 U571 ( .A1(n556), .A2(KEYINPUT64), .ZN(n555) );
  INV_X1 U572 ( .A(n730), .ZN(n556) );
  NAND2_X1 U573 ( .A1(n553), .A2(n551), .ZN(n550) );
  AND2_X1 U574 ( .A1(n730), .A2(n552), .ZN(n551) );
  INV_X1 U575 ( .A(n729), .ZN(n553) );
  INV_X1 U576 ( .A(KEYINPUT64), .ZN(n552) );
  INV_X1 U577 ( .A(n554), .ZN(n548) );
  AND2_X1 U578 ( .A1(n539), .A2(n545), .ZN(n538) );
  NAND2_X1 U579 ( .A1(n540), .A2(n542), .ZN(n541) );
  NOR2_X1 U580 ( .A1(n546), .A2(KEYINPUT33), .ZN(n542) );
  XNOR2_X1 U581 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n564) );
  AND2_X1 U582 ( .A1(G2104), .A2(G2105), .ZN(n918) );
  NAND2_X1 U583 ( .A1(n527), .A2(n717), .ZN(n526) );
  AND2_X1 U584 ( .A1(n529), .A2(n727), .ZN(n528) );
  AND2_X1 U585 ( .A1(n570), .A2(n569), .ZN(n572) );
  XNOR2_X2 U586 ( .A(n563), .B(n564), .ZN(n547) );
  OR2_X1 U587 ( .A1(G301), .A2(n685), .ZN(n521) );
  NOR2_X1 U588 ( .A1(n693), .A2(n530), .ZN(n522) );
  AND2_X1 U589 ( .A1(n535), .A2(n534), .ZN(n523) );
  NAND2_X1 U590 ( .A1(n990), .A2(n546), .ZN(n524) );
  AND2_X1 U591 ( .A1(n1007), .A2(n710), .ZN(n525) );
  NAND2_X1 U592 ( .A1(n528), .A2(n526), .ZN(n760) );
  INV_X1 U593 ( .A(n728), .ZN(n527) );
  NAND2_X1 U594 ( .A1(n728), .A2(KEYINPUT101), .ZN(n529) );
  INV_X1 U595 ( .A(n693), .ZN(n534) );
  NAND2_X1 U596 ( .A1(n522), .A2(n535), .ZN(n533) );
  INV_X1 U597 ( .A(n700), .ZN(n530) );
  NAND2_X1 U598 ( .A1(n533), .A2(n531), .ZN(n702) );
  NAND2_X1 U599 ( .A1(n700), .A2(n532), .ZN(n531) );
  INV_X1 U600 ( .A(G286), .ZN(n532) );
  INV_X1 U601 ( .A(n720), .ZN(n540) );
  NAND2_X1 U602 ( .A1(n541), .A2(n536), .ZN(n714) );
  NAND2_X1 U603 ( .A1(n537), .A2(n538), .ZN(n536) );
  NAND2_X1 U604 ( .A1(n540), .A2(n543), .ZN(n537) );
  OR2_X1 U605 ( .A1(n990), .A2(n546), .ZN(n544) );
  INV_X1 U606 ( .A(KEYINPUT33), .ZN(n545) );
  INV_X1 U607 ( .A(KEYINPUT99), .ZN(n546) );
  NAND2_X1 U608 ( .A1(n547), .A2(G137), .ZN(n565) );
  NAND2_X1 U609 ( .A1(n547), .A2(G138), .ZN(n577) );
  NAND2_X1 U610 ( .A1(n547), .A2(G136), .ZN(n889) );
  NAND2_X1 U611 ( .A1(n547), .A2(G141), .ZN(n749) );
  NAND2_X1 U612 ( .A1(n547), .A2(G140), .ZN(n731) );
  NAND2_X1 U613 ( .A1(n547), .A2(G131), .ZN(n742) );
  NAND2_X1 U614 ( .A1(n547), .A2(G139), .ZN(n902) );
  NAND2_X1 U615 ( .A1(n547), .A2(G135), .ZN(n809) );
  NAND2_X1 U616 ( .A1(n547), .A2(G142), .ZN(n915) );
  NAND2_X1 U617 ( .A1(n729), .A2(KEYINPUT64), .ZN(n557) );
  AND2_X1 U618 ( .A1(n759), .A2(n758), .ZN(n558) );
  INV_X1 U619 ( .A(G2105), .ZN(n562) );
  INV_X1 U620 ( .A(KEYINPUT27), .ZN(n639) );
  INV_X1 U621 ( .A(KEYINPUT28), .ZN(n644) );
  NOR2_X1 U622 ( .A1(G651), .A2(n619), .ZN(n817) );
  INV_X1 U623 ( .A(KEYINPUT65), .ZN(n571) );
  NAND2_X1 U624 ( .A1(G101), .A2(n914), .ZN(n559) );
  INV_X1 U625 ( .A(KEYINPUT66), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(n570) );
  AND2_X1 U627 ( .A1(G125), .A2(n921), .ZN(n568) );
  NAND2_X1 U628 ( .A1(G113), .A2(n918), .ZN(n566) );
  NOR2_X1 U629 ( .A1(G2104), .A2(G2105), .ZN(n563) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U631 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U632 ( .A1(n918), .A2(G114), .ZN(n575) );
  NAND2_X1 U633 ( .A1(G102), .A2(n914), .ZN(n573) );
  XOR2_X1 U634 ( .A(KEYINPUT91), .B(n573), .Z(n574) );
  NAND2_X1 U635 ( .A1(n575), .A2(n574), .ZN(n579) );
  NAND2_X1 U636 ( .A1(G126), .A2(n921), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U638 ( .A1(n579), .A2(n578), .ZN(G164) );
  NOR2_X1 U639 ( .A1(G651), .A2(G543), .ZN(n822) );
  NAND2_X1 U640 ( .A1(n822), .A2(G91), .ZN(n580) );
  XOR2_X1 U641 ( .A(KEYINPUT71), .B(n580), .Z(n582) );
  XOR2_X1 U642 ( .A(KEYINPUT0), .B(G543), .Z(n619) );
  INV_X1 U643 ( .A(G651), .ZN(n584) );
  NOR2_X1 U644 ( .A1(n619), .A2(n584), .ZN(n823) );
  NAND2_X1 U645 ( .A1(n823), .A2(G78), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT72), .B(n583), .Z(n590) );
  NOR2_X1 U648 ( .A1(G543), .A2(n584), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT68), .B(n585), .Z(n586) );
  XNOR2_X1 U650 ( .A(KEYINPUT1), .B(n586), .ZN(n818) );
  NAND2_X1 U651 ( .A1(n818), .A2(G65), .ZN(n588) );
  NAND2_X1 U652 ( .A1(G53), .A2(n817), .ZN(n587) );
  AND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(G299) );
  NAND2_X1 U655 ( .A1(G52), .A2(n817), .ZN(n592) );
  NAND2_X1 U656 ( .A1(G64), .A2(n818), .ZN(n591) );
  NAND2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n598) );
  NAND2_X1 U658 ( .A1(n823), .A2(G77), .ZN(n593) );
  XNOR2_X1 U659 ( .A(n593), .B(KEYINPUT70), .ZN(n595) );
  NAND2_X1 U660 ( .A1(G90), .A2(n822), .ZN(n594) );
  NAND2_X1 U661 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U662 ( .A(KEYINPUT9), .B(n596), .Z(n597) );
  NOR2_X1 U663 ( .A1(n598), .A2(n597), .ZN(G171) );
  INV_X1 U664 ( .A(G171), .ZN(G301) );
  NAND2_X1 U665 ( .A1(G51), .A2(n817), .ZN(n600) );
  NAND2_X1 U666 ( .A1(G63), .A2(n818), .ZN(n599) );
  NAND2_X1 U667 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U668 ( .A(KEYINPUT6), .B(n601), .ZN(n608) );
  NAND2_X1 U669 ( .A1(n822), .A2(G89), .ZN(n602) );
  XNOR2_X1 U670 ( .A(n602), .B(KEYINPUT4), .ZN(n604) );
  NAND2_X1 U671 ( .A1(G76), .A2(n823), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U673 ( .A(KEYINPUT5), .B(n605), .Z(n606) );
  XNOR2_X1 U674 ( .A(KEYINPUT76), .B(n606), .ZN(n607) );
  NOR2_X1 U675 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U676 ( .A(KEYINPUT7), .B(n609), .Z(G168) );
  XOR2_X1 U677 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U678 ( .A1(G88), .A2(n822), .ZN(n611) );
  NAND2_X1 U679 ( .A1(G75), .A2(n823), .ZN(n610) );
  NAND2_X1 U680 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U681 ( .A1(G50), .A2(n817), .ZN(n613) );
  NAND2_X1 U682 ( .A1(G62), .A2(n818), .ZN(n612) );
  NAND2_X1 U683 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U684 ( .A1(n615), .A2(n614), .ZN(G166) );
  XOR2_X1 U685 ( .A(KEYINPUT92), .B(G166), .Z(G303) );
  NAND2_X1 U686 ( .A1(G49), .A2(n817), .ZN(n617) );
  NAND2_X1 U687 ( .A1(G74), .A2(G651), .ZN(n616) );
  NAND2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U689 ( .A1(n818), .A2(n618), .ZN(n622) );
  NAND2_X1 U690 ( .A1(G87), .A2(n619), .ZN(n620) );
  XOR2_X1 U691 ( .A(KEYINPUT83), .B(n620), .Z(n621) );
  NAND2_X1 U692 ( .A1(n622), .A2(n621), .ZN(G288) );
  XOR2_X1 U693 ( .A(KEYINPUT85), .B(KEYINPUT2), .Z(n624) );
  NAND2_X1 U694 ( .A1(G73), .A2(n823), .ZN(n623) );
  XNOR2_X1 U695 ( .A(n624), .B(n623), .ZN(n631) );
  NAND2_X1 U696 ( .A1(G48), .A2(n817), .ZN(n626) );
  NAND2_X1 U697 ( .A1(G61), .A2(n818), .ZN(n625) );
  NAND2_X1 U698 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U699 ( .A1(n822), .A2(G86), .ZN(n627) );
  XOR2_X1 U700 ( .A(KEYINPUT84), .B(n627), .Z(n628) );
  NOR2_X1 U701 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U702 ( .A1(n631), .A2(n630), .ZN(G305) );
  NAND2_X1 U703 ( .A1(G85), .A2(n822), .ZN(n633) );
  NAND2_X1 U704 ( .A1(G72), .A2(n823), .ZN(n632) );
  NAND2_X1 U705 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U706 ( .A1(G47), .A2(n817), .ZN(n634) );
  XNOR2_X1 U707 ( .A(KEYINPUT69), .B(n634), .ZN(n635) );
  NOR2_X1 U708 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U709 ( .A1(G60), .A2(n818), .ZN(n637) );
  NAND2_X1 U710 ( .A1(n638), .A2(n637), .ZN(G290) );
  NAND2_X1 U711 ( .A1(G160), .A2(G40), .ZN(n729) );
  NOR2_X1 U712 ( .A1(G164), .A2(G1384), .ZN(n730) );
  XNOR2_X1 U713 ( .A(n640), .B(n639), .ZN(n642) );
  XNOR2_X1 U714 ( .A(KEYINPUT94), .B(G1956), .ZN(n945) );
  AND2_X1 U715 ( .A1(n945), .A2(n694), .ZN(n641) );
  INV_X1 U716 ( .A(G299), .ZN(n831) );
  XNOR2_X1 U717 ( .A(n645), .B(n644), .ZN(n679) );
  NAND2_X1 U718 ( .A1(n818), .A2(G56), .ZN(n646) );
  XOR2_X1 U719 ( .A(KEYINPUT14), .B(n646), .Z(n653) );
  NAND2_X1 U720 ( .A1(G81), .A2(n822), .ZN(n647) );
  XNOR2_X1 U721 ( .A(n647), .B(KEYINPUT74), .ZN(n648) );
  XNOR2_X1 U722 ( .A(n648), .B(KEYINPUT12), .ZN(n650) );
  NAND2_X1 U723 ( .A1(G68), .A2(n823), .ZN(n649) );
  NAND2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U725 ( .A(KEYINPUT13), .B(n651), .Z(n652) );
  NOR2_X1 U726 ( .A1(n653), .A2(n652), .ZN(n655) );
  NAND2_X1 U727 ( .A1(n817), .A2(G43), .ZN(n654) );
  NAND2_X1 U728 ( .A1(n655), .A2(n654), .ZN(n1004) );
  INV_X1 U729 ( .A(n694), .ZN(n682) );
  NAND2_X1 U730 ( .A1(n682), .A2(G1996), .ZN(n656) );
  XNOR2_X1 U731 ( .A(n656), .B(KEYINPUT26), .ZN(n658) );
  NAND2_X1 U732 ( .A1(n694), .A2(G1341), .ZN(n657) );
  NAND2_X1 U733 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U734 ( .A1(n1004), .A2(n659), .ZN(n671) );
  NAND2_X1 U735 ( .A1(n817), .A2(G54), .ZN(n666) );
  NAND2_X1 U736 ( .A1(n823), .A2(G79), .ZN(n661) );
  NAND2_X1 U737 ( .A1(G66), .A2(n818), .ZN(n660) );
  NAND2_X1 U738 ( .A1(n661), .A2(n660), .ZN(n664) );
  NAND2_X1 U739 ( .A1(G92), .A2(n822), .ZN(n662) );
  XNOR2_X1 U740 ( .A(KEYINPUT75), .B(n662), .ZN(n663) );
  NOR2_X1 U741 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U742 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U743 ( .A(KEYINPUT15), .B(n667), .Z(n993) );
  NAND2_X1 U744 ( .A1(G2067), .A2(n682), .ZN(n669) );
  NAND2_X1 U745 ( .A1(n694), .A2(G1348), .ZN(n668) );
  NAND2_X1 U746 ( .A1(n669), .A2(n668), .ZN(n672) );
  NOR2_X1 U747 ( .A1(n993), .A2(n672), .ZN(n670) );
  OR2_X1 U748 ( .A1(n671), .A2(n670), .ZN(n674) );
  NAND2_X1 U749 ( .A1(n993), .A2(n672), .ZN(n673) );
  NAND2_X1 U750 ( .A1(n674), .A2(n673), .ZN(n677) );
  NAND2_X1 U751 ( .A1(n831), .A2(n675), .ZN(n676) );
  NAND2_X1 U752 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U753 ( .A1(n679), .A2(n678), .ZN(n681) );
  XOR2_X1 U754 ( .A(G2078), .B(KEYINPUT25), .Z(n970) );
  NAND2_X1 U755 ( .A1(n970), .A2(n682), .ZN(n684) );
  NAND2_X1 U756 ( .A1(n694), .A2(G1961), .ZN(n683) );
  NAND2_X1 U757 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U758 ( .A1(G301), .A2(n685), .ZN(n686) );
  XNOR2_X1 U759 ( .A(n686), .B(KEYINPUT97), .ZN(n691) );
  NAND2_X1 U760 ( .A1(n694), .A2(G8), .ZN(n724) );
  NOR2_X1 U761 ( .A1(n694), .A2(G2084), .ZN(n703) );
  NOR2_X1 U762 ( .A1(n704), .A2(n703), .ZN(n687) );
  NAND2_X1 U763 ( .A1(G8), .A2(n687), .ZN(n688) );
  XNOR2_X1 U764 ( .A(KEYINPUT30), .B(n688), .ZN(n689) );
  NOR2_X1 U765 ( .A1(n689), .A2(G168), .ZN(n690) );
  XNOR2_X1 U766 ( .A(n692), .B(KEYINPUT31), .ZN(n693) );
  INV_X1 U767 ( .A(G8), .ZN(n699) );
  NOR2_X1 U768 ( .A1(n694), .A2(G2090), .ZN(n696) );
  NOR2_X1 U769 ( .A1(G1971), .A2(n724), .ZN(n695) );
  NOR2_X1 U770 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U771 ( .A1(G303), .A2(n697), .ZN(n698) );
  OR2_X1 U772 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U773 ( .A(n702), .B(n701), .ZN(n708) );
  NAND2_X1 U774 ( .A1(n703), .A2(G8), .ZN(n706) );
  NOR2_X1 U775 ( .A1(n704), .A2(n523), .ZN(n705) );
  NAND2_X1 U776 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U777 ( .A1(n708), .A2(n707), .ZN(n720) );
  NOR2_X1 U778 ( .A1(G1976), .A2(G288), .ZN(n711) );
  NOR2_X1 U779 ( .A1(G303), .A2(G1971), .ZN(n709) );
  NOR2_X1 U780 ( .A1(n711), .A2(n709), .ZN(n990) );
  NAND2_X1 U781 ( .A1(G1976), .A2(G288), .ZN(n1007) );
  INV_X1 U782 ( .A(n724), .ZN(n710) );
  NAND2_X1 U783 ( .A1(n711), .A2(KEYINPUT33), .ZN(n712) );
  NOR2_X1 U784 ( .A1(n712), .A2(n724), .ZN(n713) );
  NOR2_X1 U785 ( .A1(n714), .A2(n713), .ZN(n716) );
  XOR2_X1 U786 ( .A(G1981), .B(KEYINPUT100), .Z(n715) );
  XNOR2_X1 U787 ( .A(G305), .B(n715), .ZN(n1002) );
  NAND2_X1 U788 ( .A1(n716), .A2(n1002), .ZN(n728) );
  INV_X1 U789 ( .A(KEYINPUT101), .ZN(n717) );
  NOR2_X1 U790 ( .A1(G2090), .A2(G303), .ZN(n718) );
  NAND2_X1 U791 ( .A1(G8), .A2(n718), .ZN(n719) );
  NAND2_X1 U792 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U793 ( .A1(n724), .A2(n721), .ZN(n726) );
  NOR2_X1 U794 ( .A1(G1981), .A2(G305), .ZN(n722) );
  XOR2_X1 U795 ( .A(n722), .B(KEYINPUT24), .Z(n723) );
  OR2_X1 U796 ( .A1(n724), .A2(n723), .ZN(n725) );
  AND2_X1 U797 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U798 ( .A1(n730), .A2(n729), .ZN(n772) );
  XNOR2_X1 U799 ( .A(G2067), .B(KEYINPUT37), .ZN(n770) );
  NAND2_X1 U800 ( .A1(G104), .A2(n914), .ZN(n732) );
  NAND2_X1 U801 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U802 ( .A(KEYINPUT34), .B(n733), .ZN(n738) );
  NAND2_X1 U803 ( .A1(G116), .A2(n918), .ZN(n735) );
  NAND2_X1 U804 ( .A1(G128), .A2(n921), .ZN(n734) );
  NAND2_X1 U805 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U806 ( .A(KEYINPUT35), .B(n736), .Z(n737) );
  NOR2_X1 U807 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U808 ( .A(KEYINPUT36), .B(n739), .ZN(n929) );
  NOR2_X1 U809 ( .A1(n770), .A2(n929), .ZN(n1032) );
  NAND2_X1 U810 ( .A1(n772), .A2(n1032), .ZN(n768) );
  NAND2_X1 U811 ( .A1(G95), .A2(n914), .ZN(n741) );
  NAND2_X1 U812 ( .A1(G119), .A2(n921), .ZN(n740) );
  NAND2_X1 U813 ( .A1(n741), .A2(n740), .ZN(n745) );
  NAND2_X1 U814 ( .A1(G107), .A2(n918), .ZN(n743) );
  NAND2_X1 U815 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U816 ( .A1(n745), .A2(n744), .ZN(n907) );
  INV_X1 U817 ( .A(G1991), .ZN(n761) );
  NOR2_X1 U818 ( .A1(n907), .A2(n761), .ZN(n755) );
  NAND2_X1 U819 ( .A1(G105), .A2(n914), .ZN(n746) );
  XNOR2_X1 U820 ( .A(n746), .B(KEYINPUT38), .ZN(n753) );
  NAND2_X1 U821 ( .A1(G117), .A2(n918), .ZN(n748) );
  NAND2_X1 U822 ( .A1(G129), .A2(n921), .ZN(n747) );
  NAND2_X1 U823 ( .A1(n748), .A2(n747), .ZN(n751) );
  XNOR2_X1 U824 ( .A(KEYINPUT93), .B(n749), .ZN(n750) );
  NOR2_X1 U825 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U826 ( .A1(n753), .A2(n752), .ZN(n911) );
  AND2_X1 U827 ( .A1(n911), .A2(G1996), .ZN(n754) );
  NOR2_X1 U828 ( .A1(n755), .A2(n754), .ZN(n1029) );
  INV_X1 U829 ( .A(n772), .ZN(n756) );
  NOR2_X1 U830 ( .A1(n1029), .A2(n756), .ZN(n764) );
  INV_X1 U831 ( .A(n764), .ZN(n757) );
  AND2_X1 U832 ( .A1(n768), .A2(n757), .ZN(n759) );
  XNOR2_X1 U833 ( .A(G1986), .B(G290), .ZN(n1009) );
  NAND2_X1 U834 ( .A1(n1009), .A2(n772), .ZN(n758) );
  NAND2_X1 U835 ( .A1(n760), .A2(n558), .ZN(n775) );
  NOR2_X1 U836 ( .A1(G1996), .A2(n911), .ZN(n1021) );
  AND2_X1 U837 ( .A1(n761), .A2(n907), .ZN(n1034) );
  NOR2_X1 U838 ( .A1(G1986), .A2(G290), .ZN(n762) );
  NOR2_X1 U839 ( .A1(n1034), .A2(n762), .ZN(n763) );
  NOR2_X1 U840 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U841 ( .A(n765), .B(KEYINPUT102), .ZN(n766) );
  NOR2_X1 U842 ( .A1(n1021), .A2(n766), .ZN(n767) );
  XNOR2_X1 U843 ( .A(KEYINPUT39), .B(n767), .ZN(n769) );
  NAND2_X1 U844 ( .A1(n769), .A2(n768), .ZN(n771) );
  NAND2_X1 U845 ( .A1(n770), .A2(n929), .ZN(n1038) );
  NAND2_X1 U846 ( .A1(n771), .A2(n1038), .ZN(n773) );
  NAND2_X1 U847 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U848 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U849 ( .A(n776), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U850 ( .A(G2451), .B(G2427), .ZN(n786) );
  XOR2_X1 U851 ( .A(KEYINPUT103), .B(G2443), .Z(n778) );
  XNOR2_X1 U852 ( .A(G2435), .B(G2438), .ZN(n777) );
  XNOR2_X1 U853 ( .A(n778), .B(n777), .ZN(n782) );
  XOR2_X1 U854 ( .A(G2454), .B(G2430), .Z(n780) );
  XNOR2_X1 U855 ( .A(G1341), .B(G1348), .ZN(n779) );
  XNOR2_X1 U856 ( .A(n780), .B(n779), .ZN(n781) );
  XOR2_X1 U857 ( .A(n782), .B(n781), .Z(n784) );
  XNOR2_X1 U858 ( .A(G2446), .B(KEYINPUT104), .ZN(n783) );
  XNOR2_X1 U859 ( .A(n784), .B(n783), .ZN(n785) );
  XNOR2_X1 U860 ( .A(n786), .B(n785), .ZN(n787) );
  AND2_X1 U861 ( .A1(n787), .A2(G14), .ZN(G401) );
  AND2_X1 U862 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U863 ( .A(G120), .ZN(G236) );
  INV_X1 U864 ( .A(G69), .ZN(G235) );
  INV_X1 U865 ( .A(G108), .ZN(G238) );
  NAND2_X1 U866 ( .A1(G7), .A2(G661), .ZN(n788) );
  XNOR2_X1 U867 ( .A(n788), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U868 ( .A(G223), .ZN(n860) );
  NAND2_X1 U869 ( .A1(n860), .A2(G567), .ZN(n789) );
  XNOR2_X1 U870 ( .A(n789), .B(KEYINPUT11), .ZN(n790) );
  XNOR2_X1 U871 ( .A(KEYINPUT73), .B(n790), .ZN(G234) );
  INV_X1 U872 ( .A(G860), .ZN(n796) );
  OR2_X1 U873 ( .A1(n1004), .A2(n796), .ZN(G153) );
  NAND2_X1 U874 ( .A1(G868), .A2(G301), .ZN(n792) );
  INV_X1 U875 ( .A(G868), .ZN(n838) );
  NAND2_X1 U876 ( .A1(n993), .A2(n838), .ZN(n791) );
  NAND2_X1 U877 ( .A1(n792), .A2(n791), .ZN(G284) );
  NOR2_X1 U878 ( .A1(G286), .A2(n838), .ZN(n793) );
  XOR2_X1 U879 ( .A(KEYINPUT77), .B(n793), .Z(n795) );
  NOR2_X1 U880 ( .A1(G868), .A2(G299), .ZN(n794) );
  NOR2_X1 U881 ( .A1(n795), .A2(n794), .ZN(G297) );
  NAND2_X1 U882 ( .A1(n796), .A2(G559), .ZN(n797) );
  INV_X1 U883 ( .A(n993), .ZN(n815) );
  NAND2_X1 U884 ( .A1(n797), .A2(n815), .ZN(n798) );
  XNOR2_X1 U885 ( .A(n798), .B(KEYINPUT78), .ZN(n799) );
  XNOR2_X1 U886 ( .A(KEYINPUT16), .B(n799), .ZN(G148) );
  NOR2_X1 U887 ( .A1(G868), .A2(n1004), .ZN(n802) );
  NAND2_X1 U888 ( .A1(G868), .A2(n815), .ZN(n800) );
  NOR2_X1 U889 ( .A1(G559), .A2(n800), .ZN(n801) );
  NOR2_X1 U890 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U891 ( .A(KEYINPUT79), .B(n803), .Z(G282) );
  XOR2_X1 U892 ( .A(KEYINPUT80), .B(KEYINPUT18), .Z(n805) );
  NAND2_X1 U893 ( .A1(G123), .A2(n921), .ZN(n804) );
  XNOR2_X1 U894 ( .A(n805), .B(n804), .ZN(n812) );
  NAND2_X1 U895 ( .A1(G99), .A2(n914), .ZN(n807) );
  NAND2_X1 U896 ( .A1(G111), .A2(n918), .ZN(n806) );
  NAND2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U898 ( .A(n808), .B(KEYINPUT81), .ZN(n810) );
  NAND2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U900 ( .A1(n812), .A2(n811), .ZN(n1033) );
  XNOR2_X1 U901 ( .A(n1033), .B(G2096), .ZN(n814) );
  INV_X1 U902 ( .A(G2100), .ZN(n813) );
  NAND2_X1 U903 ( .A1(n814), .A2(n813), .ZN(G156) );
  NAND2_X1 U904 ( .A1(n815), .A2(G559), .ZN(n836) );
  XNOR2_X1 U905 ( .A(n1004), .B(n836), .ZN(n816) );
  NOR2_X1 U906 ( .A1(n816), .A2(G860), .ZN(n828) );
  NAND2_X1 U907 ( .A1(G55), .A2(n817), .ZN(n820) );
  NAND2_X1 U908 ( .A1(G67), .A2(n818), .ZN(n819) );
  NAND2_X1 U909 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U910 ( .A(KEYINPUT82), .B(n821), .ZN(n827) );
  NAND2_X1 U911 ( .A1(G93), .A2(n822), .ZN(n825) );
  NAND2_X1 U912 ( .A1(G80), .A2(n823), .ZN(n824) );
  NAND2_X1 U913 ( .A1(n825), .A2(n824), .ZN(n826) );
  OR2_X1 U914 ( .A1(n827), .A2(n826), .ZN(n839) );
  XOR2_X1 U915 ( .A(n828), .B(n839), .Z(G145) );
  XOR2_X1 U916 ( .A(G166), .B(KEYINPUT19), .Z(n829) );
  XNOR2_X1 U917 ( .A(n1004), .B(n829), .ZN(n830) );
  XOR2_X1 U918 ( .A(n839), .B(n830), .Z(n833) );
  XNOR2_X1 U919 ( .A(G290), .B(n831), .ZN(n832) );
  XNOR2_X1 U920 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U921 ( .A(n834), .B(G305), .ZN(n835) );
  XNOR2_X1 U922 ( .A(n835), .B(G288), .ZN(n933) );
  XOR2_X1 U923 ( .A(n933), .B(n836), .Z(n837) );
  NAND2_X1 U924 ( .A1(G868), .A2(n837), .ZN(n841) );
  NAND2_X1 U925 ( .A1(n839), .A2(n838), .ZN(n840) );
  NAND2_X1 U926 ( .A1(n841), .A2(n840), .ZN(G295) );
  NAND2_X1 U927 ( .A1(G2078), .A2(G2084), .ZN(n842) );
  XOR2_X1 U928 ( .A(KEYINPUT20), .B(n842), .Z(n843) );
  NAND2_X1 U929 ( .A1(G2090), .A2(n843), .ZN(n844) );
  XNOR2_X1 U930 ( .A(KEYINPUT21), .B(n844), .ZN(n845) );
  NAND2_X1 U931 ( .A1(n845), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U932 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U933 ( .A1(G235), .A2(G236), .ZN(n846) );
  XOR2_X1 U934 ( .A(KEYINPUT88), .B(n846), .Z(n847) );
  NOR2_X1 U935 ( .A1(G238), .A2(n847), .ZN(n848) );
  NAND2_X1 U936 ( .A1(G57), .A2(n848), .ZN(n864) );
  NAND2_X1 U937 ( .A1(G567), .A2(n864), .ZN(n849) );
  XNOR2_X1 U938 ( .A(n849), .B(KEYINPUT89), .ZN(n856) );
  XOR2_X1 U939 ( .A(KEYINPUT22), .B(KEYINPUT86), .Z(n851) );
  NAND2_X1 U940 ( .A1(G132), .A2(G82), .ZN(n850) );
  XNOR2_X1 U941 ( .A(n851), .B(n850), .ZN(n852) );
  NAND2_X1 U942 ( .A1(n852), .A2(G96), .ZN(n853) );
  NOR2_X1 U943 ( .A1(G218), .A2(n853), .ZN(n854) );
  XNOR2_X1 U944 ( .A(KEYINPUT87), .B(n854), .ZN(n865) );
  AND2_X1 U945 ( .A1(G2106), .A2(n865), .ZN(n855) );
  NOR2_X1 U946 ( .A1(n856), .A2(n855), .ZN(G319) );
  NAND2_X1 U947 ( .A1(G483), .A2(G661), .ZN(n858) );
  INV_X1 U948 ( .A(G319), .ZN(n857) );
  NOR2_X1 U949 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U950 ( .A(n859), .B(KEYINPUT90), .ZN(n863) );
  NAND2_X1 U951 ( .A1(G36), .A2(n863), .ZN(G176) );
  NAND2_X1 U952 ( .A1(G2106), .A2(n860), .ZN(G217) );
  AND2_X1 U953 ( .A1(G15), .A2(G2), .ZN(n861) );
  NAND2_X1 U954 ( .A1(G661), .A2(n861), .ZN(G259) );
  NAND2_X1 U955 ( .A1(G3), .A2(G1), .ZN(n862) );
  NAND2_X1 U956 ( .A1(n863), .A2(n862), .ZN(G188) );
  INV_X1 U958 ( .A(G132), .ZN(G219) );
  INV_X1 U959 ( .A(G96), .ZN(G221) );
  INV_X1 U960 ( .A(G82), .ZN(G220) );
  NOR2_X1 U961 ( .A1(n865), .A2(n864), .ZN(G325) );
  INV_X1 U962 ( .A(G325), .ZN(G261) );
  XOR2_X1 U963 ( .A(KEYINPUT108), .B(G1981), .Z(n867) );
  XNOR2_X1 U964 ( .A(G1956), .B(G1966), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U966 ( .A(n868), .B(KEYINPUT41), .Z(n870) );
  XNOR2_X1 U967 ( .A(G1996), .B(G1991), .ZN(n869) );
  XNOR2_X1 U968 ( .A(n870), .B(n869), .ZN(n874) );
  XOR2_X1 U969 ( .A(G1976), .B(G1961), .Z(n872) );
  XNOR2_X1 U970 ( .A(G1986), .B(G1971), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U972 ( .A(n874), .B(n873), .Z(n876) );
  XNOR2_X1 U973 ( .A(KEYINPUT107), .B(G2474), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n876), .B(n875), .ZN(G229) );
  XOR2_X1 U975 ( .A(KEYINPUT106), .B(KEYINPUT105), .Z(n878) );
  XNOR2_X1 U976 ( .A(G2678), .B(KEYINPUT43), .ZN(n877) );
  XNOR2_X1 U977 ( .A(n878), .B(n877), .ZN(n882) );
  XOR2_X1 U978 ( .A(KEYINPUT42), .B(G2072), .Z(n880) );
  XNOR2_X1 U979 ( .A(G2067), .B(G2090), .ZN(n879) );
  XNOR2_X1 U980 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U981 ( .A(n882), .B(n881), .Z(n884) );
  XNOR2_X1 U982 ( .A(G2096), .B(G2100), .ZN(n883) );
  XNOR2_X1 U983 ( .A(n884), .B(n883), .ZN(n886) );
  XOR2_X1 U984 ( .A(G2078), .B(G2084), .Z(n885) );
  XNOR2_X1 U985 ( .A(n886), .B(n885), .ZN(G227) );
  NAND2_X1 U986 ( .A1(G100), .A2(n914), .ZN(n888) );
  NAND2_X1 U987 ( .A1(G112), .A2(n918), .ZN(n887) );
  NAND2_X1 U988 ( .A1(n888), .A2(n887), .ZN(n896) );
  XNOR2_X1 U989 ( .A(KEYINPUT110), .B(n889), .ZN(n893) );
  XOR2_X1 U990 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n891) );
  NAND2_X1 U991 ( .A1(G124), .A2(n921), .ZN(n890) );
  XNOR2_X1 U992 ( .A(n891), .B(n890), .ZN(n892) );
  NAND2_X1 U993 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U994 ( .A(KEYINPUT111), .B(n894), .Z(n895) );
  NOR2_X1 U995 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U996 ( .A(KEYINPUT112), .B(n897), .ZN(G162) );
  XOR2_X1 U997 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n909) );
  NAND2_X1 U998 ( .A1(n918), .A2(G115), .ZN(n898) );
  XOR2_X1 U999 ( .A(KEYINPUT115), .B(n898), .Z(n900) );
  NAND2_X1 U1000 ( .A1(n921), .A2(G127), .ZN(n899) );
  NAND2_X1 U1001 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(n901), .B(KEYINPUT47), .ZN(n903) );
  NAND2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(n906) );
  NAND2_X1 U1004 ( .A1(n914), .A2(G103), .ZN(n904) );
  XOR2_X1 U1005 ( .A(KEYINPUT114), .B(n904), .Z(n905) );
  NOR2_X1 U1006 ( .A1(n906), .A2(n905), .ZN(n1023) );
  XNOR2_X1 U1007 ( .A(n907), .B(n1023), .ZN(n908) );
  XNOR2_X1 U1008 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(G162), .B(n910), .ZN(n913) );
  XOR2_X1 U1010 ( .A(G160), .B(n911), .Z(n912) );
  XNOR2_X1 U1011 ( .A(n913), .B(n912), .ZN(n926) );
  NAND2_X1 U1012 ( .A1(G106), .A2(n914), .ZN(n916) );
  NAND2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(n917), .B(KEYINPUT45), .ZN(n920) );
  NAND2_X1 U1015 ( .A1(G118), .A2(n918), .ZN(n919) );
  NAND2_X1 U1016 ( .A1(n920), .A2(n919), .ZN(n924) );
  NAND2_X1 U1017 ( .A1(G130), .A2(n921), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(KEYINPUT113), .B(n922), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1020 ( .A(n926), .B(n925), .Z(n928) );
  XNOR2_X1 U1021 ( .A(G164), .B(n1033), .ZN(n927) );
  XNOR2_X1 U1022 ( .A(n928), .B(n927), .ZN(n930) );
  XNOR2_X1 U1023 ( .A(n930), .B(n929), .ZN(n931) );
  NOR2_X1 U1024 ( .A1(G37), .A2(n931), .ZN(G395) );
  XNOR2_X1 U1025 ( .A(G286), .B(G301), .ZN(n932) );
  XNOR2_X1 U1026 ( .A(n932), .B(n993), .ZN(n934) );
  XNOR2_X1 U1027 ( .A(n934), .B(n933), .ZN(n935) );
  NOR2_X1 U1028 ( .A1(G37), .A2(n935), .ZN(G397) );
  NOR2_X1 U1029 ( .A1(G229), .A2(G227), .ZN(n936) );
  XOR2_X1 U1030 ( .A(KEYINPUT49), .B(n936), .Z(n937) );
  NAND2_X1 U1031 ( .A1(G319), .A2(n937), .ZN(n938) );
  NOR2_X1 U1032 ( .A1(G401), .A2(n938), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(KEYINPUT116), .B(n939), .ZN(n941) );
  NOR2_X1 U1034 ( .A1(G395), .A2(G397), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(G225) );
  INV_X1 U1036 ( .A(G225), .ZN(G308) );
  INV_X1 U1037 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1038 ( .A(G1961), .B(G5), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(G1966), .B(G21), .ZN(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n954) );
  XOR2_X1 U1041 ( .A(G1348), .B(KEYINPUT59), .Z(n944) );
  XNOR2_X1 U1042 ( .A(G4), .B(n944), .ZN(n947) );
  XNOR2_X1 U1043 ( .A(G20), .B(n945), .ZN(n946) );
  NOR2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(G1341), .B(G19), .ZN(n949) );
  XNOR2_X1 U1046 ( .A(G1981), .B(G6), .ZN(n948) );
  NOR2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1049 ( .A(KEYINPUT60), .B(n952), .Z(n953) );
  NAND2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n961) );
  XNOR2_X1 U1051 ( .A(G1971), .B(G22), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(G23), .B(G1976), .ZN(n955) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n958) );
  XOR2_X1 U1054 ( .A(G1986), .B(G24), .Z(n957) );
  NAND2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1056 ( .A(KEYINPUT58), .B(n959), .ZN(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1058 ( .A(KEYINPUT61), .B(n962), .Z(n963) );
  NOR2_X1 U1059 ( .A1(G16), .A2(n963), .ZN(n964) );
  XOR2_X1 U1060 ( .A(KEYINPUT127), .B(n964), .Z(n988) );
  NOR2_X1 U1061 ( .A1(KEYINPUT55), .A2(G29), .ZN(n985) );
  XNOR2_X1 U1062 ( .A(G2090), .B(G35), .ZN(n980) );
  XNOR2_X1 U1063 ( .A(G1996), .B(G32), .ZN(n965) );
  XNOR2_X1 U1064 ( .A(n965), .B(KEYINPUT119), .ZN(n969) );
  XNOR2_X1 U1065 ( .A(G2067), .B(G26), .ZN(n967) );
  XNOR2_X1 U1066 ( .A(G33), .B(G2072), .ZN(n966) );
  NOR2_X1 U1067 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1068 ( .A1(n969), .A2(n968), .ZN(n973) );
  XNOR2_X1 U1069 ( .A(G27), .B(n970), .ZN(n971) );
  XNOR2_X1 U1070 ( .A(KEYINPUT118), .B(n971), .ZN(n972) );
  NOR2_X1 U1071 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1072 ( .A(KEYINPUT120), .B(n974), .ZN(n975) );
  NAND2_X1 U1073 ( .A1(n975), .A2(G28), .ZN(n977) );
  XNOR2_X1 U1074 ( .A(G25), .B(G1991), .ZN(n976) );
  NOR2_X1 U1075 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1076 ( .A(KEYINPUT53), .B(n978), .ZN(n979) );
  NOR2_X1 U1077 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1078 ( .A(KEYINPUT121), .B(n981), .Z(n984) );
  XOR2_X1 U1079 ( .A(G34), .B(KEYINPUT54), .Z(n982) );
  XNOR2_X1 U1080 ( .A(G2084), .B(n982), .ZN(n983) );
  NAND2_X1 U1081 ( .A1(n984), .A2(n983), .ZN(n1019) );
  NAND2_X1 U1082 ( .A1(n985), .A2(n1019), .ZN(n986) );
  NAND2_X1 U1083 ( .A1(G11), .A2(n986), .ZN(n987) );
  NOR2_X1 U1084 ( .A1(n988), .A2(n987), .ZN(n1018) );
  NAND2_X1 U1085 ( .A1(G303), .A2(G1971), .ZN(n989) );
  NAND2_X1 U1086 ( .A1(n990), .A2(n989), .ZN(n992) );
  XNOR2_X1 U1087 ( .A(G1956), .B(G299), .ZN(n991) );
  NOR2_X1 U1088 ( .A1(n992), .A2(n991), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(G1348), .B(n993), .ZN(n996) );
  XNOR2_X1 U1090 ( .A(G171), .B(G1961), .ZN(n994) );
  XNOR2_X1 U1091 ( .A(n994), .B(KEYINPUT123), .ZN(n995) );
  NOR2_X1 U1092 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1093 ( .A(n997), .B(KEYINPUT124), .ZN(n998) );
  NAND2_X1 U1094 ( .A1(n999), .A2(n998), .ZN(n1013) );
  XNOR2_X1 U1095 ( .A(G168), .B(G1966), .ZN(n1000) );
  XNOR2_X1 U1096 ( .A(n1000), .B(KEYINPUT122), .ZN(n1001) );
  NAND2_X1 U1097 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1098 ( .A(n1003), .B(KEYINPUT57), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(G1341), .B(KEYINPUT125), .ZN(n1005) );
  XNOR2_X1 U1100 ( .A(n1005), .B(n1004), .ZN(n1006) );
  NAND2_X1 U1101 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1102 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1103 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1105 ( .A(KEYINPUT126), .B(n1014), .Z(n1016) );
  XNOR2_X1 U1106 ( .A(G16), .B(KEYINPUT56), .ZN(n1015) );
  NAND2_X1 U1107 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1049) );
  INV_X1 U1109 ( .A(KEYINPUT55), .ZN(n1043) );
  OR2_X1 U1110 ( .A1(n1043), .A2(n1019), .ZN(n1047) );
  XOR2_X1 U1111 ( .A(G2090), .B(G162), .Z(n1020) );
  NOR2_X1 U1112 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1113 ( .A(KEYINPUT51), .B(n1022), .Z(n1028) );
  XOR2_X1 U1114 ( .A(G2072), .B(n1023), .Z(n1025) );
  XOR2_X1 U1115 ( .A(G164), .B(G2078), .Z(n1024) );
  NOR2_X1 U1116 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1117 ( .A(KEYINPUT50), .B(n1026), .ZN(n1027) );
  NAND2_X1 U1118 ( .A1(n1028), .A2(n1027), .ZN(n1041) );
  XNOR2_X1 U1119 ( .A(G160), .B(G2084), .ZN(n1030) );
  NAND2_X1 U1120 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1121 ( .A1(n1032), .A2(n1031), .ZN(n1036) );
  NOR2_X1 U1122 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1123 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XNOR2_X1 U1124 ( .A(KEYINPUT117), .B(n1037), .ZN(n1039) );
  NAND2_X1 U1125 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NOR2_X1 U1126 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  XNOR2_X1 U1127 ( .A(n1042), .B(KEYINPUT52), .ZN(n1044) );
  NAND2_X1 U1128 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  NAND2_X1 U1129 ( .A1(G29), .A2(n1045), .ZN(n1046) );
  NAND2_X1 U1130 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  NOR2_X1 U1131 ( .A1(n1049), .A2(n1048), .ZN(n1050) );
  XNOR2_X1 U1132 ( .A(KEYINPUT62), .B(n1050), .ZN(G311) );
  INV_X1 U1133 ( .A(G311), .ZN(G150) );
endmodule

