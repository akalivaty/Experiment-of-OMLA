//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n797, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018;
  INV_X1    g000(.A(G120gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G113gat), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G120gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n207));
  XNOR2_X1  g006(.A(G127gat), .B(G134gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT68), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n206), .B(new_n207), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G134gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G127gat), .ZN(new_n212));
  INV_X1    g011(.A(G127gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G134gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n209), .A2(new_n207), .ZN(new_n216));
  XNOR2_X1  g015(.A(G113gat), .B(G120gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n210), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT24), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT24), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(G183gat), .A3(G190gat), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT66), .B(G190gat), .ZN(new_n226));
  INV_X1    g025(.A(G183gat), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT67), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT66), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G190gat), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n230), .A2(new_n232), .A3(KEYINPUT67), .A4(new_n227), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n225), .B1(new_n228), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NOR3_X1   g036(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT25), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G169gat), .A2(G176gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT64), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(G169gat), .A3(G176gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT65), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n241), .A2(new_n243), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n239), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT23), .ZN(new_n249));
  INV_X1    g048(.A(G169gat), .ZN(new_n250));
  INV_X1    g049(.A(G176gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n236), .ZN(new_n253));
  NOR2_X1   g052(.A1(G183gat), .A2(G190gat), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n244), .B(new_n253), .C1(new_n224), .C2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n235), .A2(new_n248), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n258));
  OR3_X1    g057(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n244), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n220), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT27), .B(G183gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n226), .A2(new_n262), .A3(KEYINPUT28), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT28), .B1(new_n226), .B2(new_n262), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n261), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n219), .B1(new_n257), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n253), .A2(new_n244), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n254), .B1(new_n221), .B2(new_n223), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n256), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n230), .A2(new_n232), .A3(new_n227), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n224), .B1(new_n273), .B2(new_n233), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n256), .B1(new_n252), .B2(new_n236), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n241), .A2(new_n243), .A3(new_n246), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n246), .B1(new_n241), .B2(new_n243), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n270), .B1(new_n274), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n219), .ZN(new_n280));
  INV_X1    g079(.A(new_n263), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n220), .B(new_n260), .C1(new_n281), .C2(new_n264), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n283), .ZN(new_n284));
  AND2_X1   g083(.A1(G227gat), .A2(G233gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(KEYINPUT34), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n284), .A2(KEYINPUT70), .A3(new_n285), .ZN(new_n291));
  XNOR2_X1  g090(.A(G15gat), .B(G43gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(G71gat), .B(G99gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n280), .B1(new_n279), .B2(new_n282), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n285), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n294), .B1(new_n297), .B2(KEYINPUT32), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT33), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  OR2_X1    g099(.A1(new_n294), .A2(new_n299), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n297), .A2(KEYINPUT32), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT69), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n297), .A2(KEYINPUT69), .A3(KEYINPUT32), .A4(new_n301), .ZN(new_n305));
  AOI221_X4 g104(.A(new_n291), .B1(new_n298), .B2(new_n300), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n291), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n305), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n298), .A2(new_n300), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n290), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT32), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n312), .B1(new_n284), .B2(new_n285), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT69), .B1(new_n313), .B2(new_n301), .ZN(new_n314));
  INV_X1    g113(.A(new_n305), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n309), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(new_n291), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n308), .A2(new_n307), .A3(new_n309), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n318), .A3(new_n289), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n311), .A2(KEYINPUT36), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT36), .B1(new_n311), .B2(new_n319), .ZN(new_n321));
  XOR2_X1   g120(.A(G78gat), .B(G106gat), .Z(new_n322));
  XNOR2_X1  g121(.A(new_n322), .B(KEYINPUT78), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT31), .B(G50gat), .ZN(new_n324));
  XOR2_X1   g123(.A(new_n323), .B(new_n324), .Z(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT2), .ZN(new_n328));
  OR2_X1    g127(.A1(G141gat), .A2(G148gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(G141gat), .A2(G148gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AND2_X1   g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT73), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G155gat), .ZN(new_n335));
  INV_X1    g134(.A(G162gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT73), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n338), .A3(new_n327), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n331), .A2(new_n334), .A3(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n332), .A2(new_n333), .ZN(new_n341));
  AND2_X1   g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(G141gat), .A2(G148gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n341), .A2(new_n344), .A3(new_n338), .A4(new_n328), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n340), .A2(new_n345), .A3(KEYINPUT74), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n340), .A2(new_n345), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G211gat), .B(G218gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G211gat), .A2(G218gat), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT22), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(KEYINPUT71), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G197gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G204gat), .ZN(new_n356));
  INV_X1    g155(.A(G204gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G197gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n354), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(KEYINPUT71), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n351), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  OR2_X1    g161(.A1(new_n360), .A2(KEYINPUT71), .ZN(new_n363));
  XNOR2_X1  g162(.A(G197gat), .B(G204gat), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n363), .A2(new_n350), .A3(new_n354), .A4(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT29), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n346), .B(new_n349), .C1(new_n366), .C2(KEYINPUT3), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n362), .A2(new_n365), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT3), .B1(new_n340), .B2(new_n345), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n369), .B1(KEYINPUT29), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G228gat), .A2(G233gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n367), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n340), .A2(new_n345), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(new_n366), .B2(KEYINPUT3), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT80), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT80), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n378), .B(new_n375), .C1(new_n366), .C2(KEYINPUT3), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n377), .A2(new_n379), .A3(new_n371), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n372), .B(KEYINPUT79), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n374), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT81), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n326), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(G22gat), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n382), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n386), .B1(new_n382), .B2(new_n383), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n385), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n380), .A2(new_n381), .ZN(new_n391));
  INV_X1    g190(.A(new_n374), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n383), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(G22gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(new_n384), .A3(new_n387), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G1gat), .B(G29gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT0), .ZN(new_n398));
  XNOR2_X1  g197(.A(G57gat), .B(G85gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n398), .A2(new_n399), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT77), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n375), .A2(new_n219), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n340), .A2(new_n345), .A3(KEYINPUT74), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT74), .B1(new_n340), .B2(new_n345), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n405), .B1(new_n408), .B2(new_n219), .ZN(new_n409));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(KEYINPUT75), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n404), .B(KEYINPUT5), .C1(new_n409), .C2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n349), .A2(new_n219), .A3(new_n346), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n280), .A2(new_n347), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT5), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT77), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n349), .A2(KEYINPUT3), .A3(new_n346), .ZN(new_n419));
  INV_X1    g218(.A(new_n370), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n219), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT4), .B1(new_n375), .B2(new_n219), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT4), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n280), .A2(new_n423), .A3(new_n347), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT76), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n422), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n415), .A2(KEYINPUT76), .A3(KEYINPUT4), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n421), .A2(new_n426), .A3(new_n412), .A4(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n413), .A2(new_n418), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n422), .A2(new_n424), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n421), .A2(new_n417), .A3(new_n412), .A4(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n403), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT6), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n429), .A2(new_n431), .A3(new_n403), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n432), .A2(KEYINPUT6), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(G226gat), .ZN(new_n439));
  INV_X1    g238(.A(G233gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT72), .B1(new_n257), .B2(new_n266), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT72), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n279), .A2(new_n444), .A3(new_n282), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n442), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  AOI211_X1 g245(.A(KEYINPUT29), .B(new_n441), .C1(new_n279), .C2(new_n282), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n368), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G8gat), .B(G36gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(G64gat), .B(G92gat), .ZN(new_n450));
  XOR2_X1   g249(.A(new_n449), .B(new_n450), .Z(new_n451));
  NOR2_X1   g250(.A1(new_n441), .A2(KEYINPUT29), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n443), .A2(new_n445), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n279), .A2(new_n441), .A3(new_n282), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(new_n369), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n448), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT30), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n448), .A2(new_n455), .ZN(new_n459));
  INV_X1    g258(.A(new_n451), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n448), .A2(KEYINPUT30), .A3(new_n451), .A4(new_n455), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n458), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n396), .B1(new_n438), .B2(new_n464), .ZN(new_n465));
  NOR3_X1   g264(.A1(new_n320), .A2(new_n321), .A3(new_n465), .ZN(new_n466));
  AOI211_X1 g265(.A(new_n434), .B(new_n403), .C1(new_n429), .C2(new_n431), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n435), .A2(new_n434), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n403), .A2(KEYINPUT82), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT82), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n401), .A2(new_n402), .A3(new_n470), .ZN(new_n471));
  OR2_X1    g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n472), .B1(new_n429), .B2(new_n431), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n467), .B1(new_n468), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n459), .A2(KEYINPUT37), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT85), .B(KEYINPUT37), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n448), .A2(new_n455), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n460), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT38), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n369), .B1(new_n446), .B2(new_n447), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n453), .A2(new_n368), .A3(new_n454), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(KEYINPUT37), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT38), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n483), .A2(new_n478), .A3(new_n484), .A4(new_n460), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n475), .A2(new_n456), .A3(new_n480), .A4(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT40), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n421), .A2(new_n430), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n411), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT39), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n490), .B1(new_n409), .B2(new_n412), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n487), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AOI211_X1 g291(.A(KEYINPUT39), .B(new_n412), .C1(new_n421), .C2(new_n430), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT83), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n469), .A2(new_n471), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n488), .A2(new_n490), .A3(new_n411), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT83), .B1(new_n497), .B2(new_n472), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n492), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n494), .B1(new_n493), .B2(new_n495), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n472), .A3(KEYINPUT83), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n500), .A2(new_n501), .B1(new_n489), .B2(new_n491), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n499), .B(new_n474), .C1(new_n502), .C2(KEYINPUT40), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT84), .B1(new_n503), .B2(new_n464), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n502), .A2(KEYINPUT40), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT84), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n500), .A2(new_n501), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n473), .B1(new_n507), .B2(new_n492), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n505), .A2(new_n506), .A3(new_n463), .A4(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n486), .A2(new_n504), .A3(new_n509), .A4(new_n396), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n463), .B1(new_n436), .B2(new_n437), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n306), .A2(new_n310), .A3(new_n290), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n289), .B1(new_n317), .B2(new_n318), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n511), .B(new_n396), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT35), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n394), .A2(new_n387), .A3(new_n384), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n384), .B1(new_n394), .B2(new_n387), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n518), .B1(new_n311), .B2(new_n319), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT35), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT86), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(new_n475), .B2(new_n463), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n435), .A2(new_n434), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n437), .B1(new_n523), .B2(new_n473), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n464), .A2(new_n524), .A3(KEYINPUT86), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n519), .A2(new_n520), .A3(new_n522), .A4(new_n525), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n466), .A2(new_n510), .B1(new_n515), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G113gat), .B(G141gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(G197gat), .ZN(new_n529));
  XOR2_X1   g328(.A(KEYINPUT11), .B(G169gat), .Z(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT87), .B(KEYINPUT12), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n531), .B(new_n532), .Z(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n534));
  INV_X1    g333(.A(G29gat), .ZN(new_n535));
  INV_X1    g334(.A(G36gat), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(new_n536), .A3(KEYINPUT14), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT14), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(G29gat), .B2(G36gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(G29gat), .A2(G36gat), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n537), .A2(new_n539), .A3(KEYINPUT15), .A4(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G43gat), .B(G50gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n542), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT15), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n543), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(G1gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT16), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n386), .A2(G15gat), .ZN(new_n552));
  INV_X1    g351(.A(G15gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(G22gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G15gat), .B(G22gat), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n555), .B1(G1gat), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(G8gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT89), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(new_n556), .B2(G1gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  OAI221_X1 g360(.A(new_n555), .B1(new_n559), .B2(G8gat), .C1(G1gat), .C2(new_n556), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT90), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n561), .A2(new_n562), .A3(KEYINPUT90), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n549), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT17), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n568), .B1(new_n549), .B2(KEYINPUT88), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n537), .A2(new_n540), .ZN(new_n570));
  INV_X1    g369(.A(new_n542), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n570), .A2(new_n571), .A3(KEYINPUT15), .A4(new_n539), .ZN(new_n572));
  AND2_X1   g371(.A1(new_n546), .A2(new_n547), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n572), .B1(new_n573), .B2(new_n544), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT88), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(new_n575), .A3(KEYINPUT17), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n567), .B1(new_n577), .B2(new_n563), .ZN(new_n578));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n534), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n574), .A2(new_n575), .A3(KEYINPUT17), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT17), .B1(new_n574), .B2(new_n575), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n563), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n566), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT90), .B1(new_n561), .B2(new_n562), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n574), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n583), .A2(KEYINPUT18), .A3(new_n579), .A4(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n579), .B(KEYINPUT13), .Z(new_n588));
  NOR3_X1   g387(.A1(new_n584), .A2(new_n585), .A3(new_n574), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n588), .B1(new_n589), .B2(new_n567), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n533), .B1(new_n580), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n583), .A2(new_n579), .A3(new_n586), .ZN(new_n593));
  INV_X1    g392(.A(new_n534), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n533), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n595), .A2(new_n596), .A3(new_n587), .A4(new_n590), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT92), .B1(new_n527), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n465), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n311), .A2(new_n319), .A3(KEYINPUT36), .ZN(new_n602));
  INV_X1    g401(.A(new_n321), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n510), .A2(new_n601), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n515), .A2(new_n526), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT92), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n606), .A2(new_n607), .A3(new_n598), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n600), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(G64gat), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n610), .A2(G57gat), .ZN(new_n611));
  INV_X1    g410(.A(G57gat), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(G64gat), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT9), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G71gat), .A2(G78gat), .ZN(new_n615));
  OR2_X1    g414(.A1(G71gat), .A2(G78gat), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT93), .B1(new_n610), .B2(G57gat), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT93), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n619), .A2(new_n612), .A3(G64gat), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n618), .B(new_n620), .C1(new_n612), .C2(G64gat), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT9), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n615), .B1(new_n616), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n617), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT94), .B(KEYINPUT21), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(G127gat), .ZN(new_n630));
  AOI211_X1 g429(.A(new_n585), .B(new_n584), .C1(KEYINPUT21), .C2(new_n625), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(new_n335), .ZN(new_n634));
  XNOR2_X1  g433(.A(G183gat), .B(G211gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n632), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G190gat), .B(G218gat), .ZN(new_n639));
  NAND2_X1  g438(.A1(G85gat), .A2(G92gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT7), .ZN(new_n641));
  INV_X1    g440(.A(G92gat), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT95), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT95), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(G92gat), .ZN(new_n645));
  INV_X1    g444(.A(G85gat), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n643), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT96), .ZN(new_n648));
  INV_X1    g447(.A(G99gat), .ZN(new_n649));
  INV_X1    g448(.A(G106gat), .ZN(new_n650));
  OAI21_X1  g449(.A(KEYINPUT8), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n647), .A2(new_n648), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n648), .B1(new_n647), .B2(new_n651), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n641), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G99gat), .B(G106gat), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n655), .B(new_n641), .C1(new_n652), .C2(new_n653), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n577), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n657), .A2(new_n574), .A3(new_n658), .ZN(new_n661));
  NAND3_X1  g460(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n639), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n577), .A2(new_n659), .ZN(new_n665));
  INV_X1    g464(.A(new_n639), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n665), .A2(new_n666), .A3(new_n661), .A4(new_n662), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n665), .A2(new_n661), .A3(new_n662), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT97), .B1(new_n669), .B2(new_n639), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(G134gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(new_n336), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n668), .B1(new_n670), .B2(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n664), .A2(KEYINPUT97), .A3(new_n667), .A4(new_n673), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(G230gat), .A2(G233gat), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n679), .B(KEYINPUT98), .Z(new_n680));
  INV_X1    g479(.A(new_n625), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n647), .A2(new_n651), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(KEYINPUT96), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n647), .A2(new_n648), .A3(new_n651), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n655), .B1(new_n685), .B2(new_n641), .ZN(new_n686));
  INV_X1    g485(.A(new_n658), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n681), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT10), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n657), .A2(new_n658), .A3(new_n625), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n657), .A2(KEYINPUT10), .A3(new_n658), .A4(new_n625), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n680), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n688), .A2(new_n690), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(new_n694), .B2(new_n680), .ZN(new_n695));
  XNOR2_X1  g494(.A(G120gat), .B(G148gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(G176gat), .B(G204gat), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n696), .B(new_n697), .Z(new_n698));
  OR2_X1    g497(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n691), .A2(new_n692), .ZN(new_n700));
  INV_X1    g499(.A(new_n680), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n694), .A2(new_n680), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(new_n703), .A3(new_n698), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n638), .A2(new_n678), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n609), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n438), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(new_n550), .ZN(G1324gat));
  INV_X1    g508(.A(KEYINPUT42), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n707), .A2(new_n464), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT16), .B(G8gat), .Z(new_n712));
  AOI21_X1  g511(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(G8gat), .B1(new_n707), .B2(new_n464), .ZN(new_n714));
  NOR2_X1   g513(.A1(KEYINPUT99), .A2(KEYINPUT42), .ZN(new_n715));
  MUX2_X1   g514(.A(KEYINPUT99), .B(new_n715), .S(new_n712), .Z(new_n716));
  AOI22_X1  g515(.A1(new_n713), .A2(new_n714), .B1(new_n711), .B2(new_n716), .ZN(G1325gat));
  NAND3_X1  g516(.A1(new_n603), .A2(KEYINPUT100), .A3(new_n602), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT100), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n320), .B2(new_n321), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(G15gat), .B1(new_n707), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n311), .A2(new_n319), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n553), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n723), .B1(new_n707), .B2(new_n725), .ZN(G1326gat));
  NOR2_X1   g525(.A1(new_n707), .A2(new_n396), .ZN(new_n727));
  XOR2_X1   g526(.A(KEYINPUT43), .B(G22gat), .Z(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1327gat));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n632), .B(new_n636), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n731), .A2(new_n677), .A3(new_n705), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT101), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n609), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n438), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n535), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n730), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  OR3_X1    g536(.A1(new_n734), .A2(new_n730), .A3(new_n736), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n527), .B2(new_n677), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n606), .A2(KEYINPUT44), .A3(new_n678), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n731), .B(KEYINPUT103), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n592), .A2(KEYINPUT102), .A3(new_n597), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT102), .B1(new_n592), .B2(new_n597), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n743), .A2(new_n705), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n742), .A2(new_n735), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT104), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G29gat), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n749), .A2(KEYINPUT104), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n737), .B(new_n738), .C1(new_n751), .C2(new_n752), .ZN(G1328gat));
  NOR2_X1   g552(.A1(new_n464), .A2(G36gat), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  OR3_X1    g554(.A1(new_n734), .A2(KEYINPUT46), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(KEYINPUT46), .B1(new_n734), .B2(new_n755), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n742), .A2(new_n463), .A3(new_n748), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n756), .B(new_n757), .C1(new_n536), .C2(new_n758), .ZN(G1329gat));
  NAND2_X1  g558(.A1(new_n603), .A2(new_n602), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n742), .A2(new_n760), .A3(new_n748), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G43gat), .ZN(new_n762));
  INV_X1    g561(.A(new_n734), .ZN(new_n763));
  INV_X1    g562(.A(new_n724), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(G43gat), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n762), .A2(new_n766), .A3(KEYINPUT47), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n742), .A2(new_n721), .A3(new_n748), .ZN(new_n768));
  AOI22_X1  g567(.A1(new_n768), .A2(G43gat), .B1(new_n763), .B2(new_n765), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n769), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g569(.A(G50gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n734), .B2(new_n396), .ZN(new_n772));
  NOR2_X1   g571(.A1(KEYINPUT105), .A2(KEYINPUT48), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n396), .A2(new_n771), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n740), .A2(new_n741), .A3(new_n748), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(KEYINPUT105), .A2(KEYINPUT48), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n772), .A2(new_n774), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n774), .B1(new_n772), .B2(new_n778), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(G1331gat));
  INV_X1    g580(.A(new_n705), .ZN(new_n782));
  NOR4_X1   g581(.A1(new_n638), .A2(new_n782), .A3(new_n746), .A4(new_n678), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n606), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n438), .B(KEYINPUT106), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XOR2_X1   g586(.A(KEYINPUT107), .B(G57gat), .Z(new_n788));
  XNOR2_X1  g587(.A(new_n787), .B(new_n788), .ZN(G1332gat));
  AOI211_X1 g588(.A(new_n464), .B(new_n784), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n790));
  NOR2_X1   g589(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n790), .B(new_n791), .ZN(G1333gat));
  OAI21_X1  g591(.A(G71gat), .B1(new_n784), .B2(new_n722), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n764), .A2(G71gat), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n784), .B2(new_n794), .ZN(new_n795));
  XOR2_X1   g594(.A(new_n795), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g595(.A1(new_n785), .A2(new_n518), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g597(.A1(new_n731), .A2(new_n746), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n606), .A2(new_n678), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n606), .A2(KEYINPUT51), .A3(new_n678), .A4(new_n799), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n782), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n804), .A2(new_n646), .A3(new_n735), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n799), .A2(new_n705), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n740), .A2(new_n741), .A3(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT108), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n740), .A2(new_n741), .A3(KEYINPUT108), .A4(new_n807), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n810), .A2(new_n735), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n805), .B1(new_n812), .B2(new_n646), .ZN(G1336gat));
  NAND2_X1  g612(.A1(new_n802), .A2(new_n803), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n464), .A2(G92gat), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(new_n705), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT109), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT109), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n804), .A2(new_n818), .A3(new_n815), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n740), .A2(new_n741), .A3(new_n463), .A4(new_n807), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n643), .A2(new_n645), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT52), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n817), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n810), .A2(new_n463), .A3(new_n811), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n824), .A2(new_n821), .B1(new_n804), .B2(new_n815), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(G1337gat));
  NAND3_X1  g626(.A1(new_n810), .A2(new_n721), .A3(new_n811), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT110), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT110), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n810), .A2(new_n830), .A3(new_n721), .A4(new_n811), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n829), .A2(G99gat), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n804), .A2(new_n649), .A3(new_n724), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(G1338gat));
  NAND4_X1  g633(.A1(new_n740), .A2(new_n741), .A3(new_n518), .A4(new_n807), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n650), .B1(new_n835), .B2(KEYINPUT113), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n836), .B1(KEYINPUT113), .B2(new_n835), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n518), .A2(new_n650), .A3(new_n705), .ZN(new_n838));
  XOR2_X1   g637(.A(new_n838), .B(KEYINPUT111), .Z(new_n839));
  AOI21_X1  g638(.A(KEYINPUT53), .B1(new_n814), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n810), .A2(new_n518), .A3(new_n811), .ZN(new_n842));
  XOR2_X1   g641(.A(new_n839), .B(KEYINPUT112), .Z(new_n843));
  AOI22_X1  g642(.A1(new_n842), .A2(G106gat), .B1(new_n814), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n841), .B1(new_n844), .B2(new_n845), .ZN(G1339gat));
  XNOR2_X1  g645(.A(new_n638), .B(KEYINPUT103), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT114), .ZN(new_n848));
  INV_X1    g647(.A(new_n691), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n692), .A2(new_n680), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n691), .A2(KEYINPUT114), .A3(new_n692), .A4(new_n680), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n851), .A2(new_n702), .A3(KEYINPUT54), .A4(new_n852), .ZN(new_n853));
  XOR2_X1   g652(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n854));
  AOI21_X1  g653(.A(new_n698), .B1(new_n693), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(KEYINPUT55), .A3(new_n855), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n856), .A2(new_n704), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT55), .B1(new_n853), .B2(new_n855), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI211_X1 g659(.A(KEYINPUT116), .B(KEYINPUT55), .C1(new_n853), .C2(new_n855), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n746), .B(new_n857), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT117), .B1(new_n578), .B2(new_n579), .ZN(new_n863));
  OR3_X1    g662(.A1(new_n589), .A2(new_n567), .A3(new_n588), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n578), .A2(KEYINPUT117), .A3(new_n579), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n531), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n705), .A2(new_n597), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n678), .B1(new_n862), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n856), .A2(new_n704), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n867), .A2(new_n675), .A3(new_n597), .A4(new_n676), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n853), .A2(new_n855), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT55), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT116), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n859), .ZN(new_n876));
  AOI211_X1 g675(.A(new_n870), .B(new_n871), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n847), .B1(new_n869), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n706), .A2(new_n747), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n518), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n880), .A2(new_n735), .A3(new_n464), .A4(new_n724), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n881), .A2(new_n204), .A3(new_n599), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n862), .A2(new_n868), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n877), .B1(new_n883), .B2(new_n677), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n879), .B1(new_n884), .B2(new_n743), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n519), .A3(new_n786), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n463), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n885), .A2(KEYINPUT118), .A3(new_n519), .A4(new_n786), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n746), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n882), .B1(new_n890), .B2(new_n204), .ZN(G1340gat));
  NOR3_X1   g690(.A1(new_n881), .A2(new_n202), .A3(new_n782), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n888), .A2(new_n705), .A3(new_n889), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(new_n202), .ZN(G1341gat));
  NOR3_X1   g693(.A1(new_n881), .A2(new_n213), .A3(new_n847), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n888), .A2(KEYINPUT119), .A3(new_n731), .A4(new_n889), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n896), .A2(new_n213), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n888), .A2(new_n889), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(new_n638), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n895), .B1(new_n897), .B2(new_n900), .ZN(G1342gat));
  NAND2_X1  g700(.A1(new_n678), .A2(new_n211), .ZN(new_n902));
  OR3_X1    g701(.A1(new_n899), .A2(KEYINPUT56), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(G134gat), .B1(new_n881), .B2(new_n677), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT56), .B1(new_n899), .B2(new_n902), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(G1343gat));
  NOR3_X1   g705(.A1(new_n760), .A2(new_n438), .A3(new_n463), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT57), .B1(new_n885), .B2(new_n518), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n518), .A2(KEYINPUT57), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(new_n870), .B2(new_n858), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n874), .A2(KEYINPUT120), .A3(new_n704), .A4(new_n856), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n598), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n678), .B1(new_n913), .B2(new_n868), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n638), .B1(new_n914), .B2(new_n877), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n909), .B1(new_n915), .B2(new_n879), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n598), .B(new_n907), .C1(new_n908), .C2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n915), .A2(new_n879), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n396), .B1(new_n878), .B2(new_n879), .ZN(new_n921));
  OAI22_X1  g720(.A1(new_n920), .A2(new_n909), .B1(new_n921), .B2(KEYINPUT57), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n922), .A2(KEYINPUT122), .A3(new_n598), .A4(new_n907), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n919), .A2(new_n923), .A3(G141gat), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n721), .A2(new_n463), .A3(new_n396), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n786), .A3(new_n885), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n599), .A2(G141gat), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT58), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n746), .B(new_n907), .C1(new_n908), .C2(new_n916), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n931), .A2(G141gat), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n925), .A2(new_n786), .A3(new_n885), .A4(new_n928), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT121), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT58), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n930), .A2(new_n935), .ZN(G1344gat));
  INV_X1    g735(.A(KEYINPUT57), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n937), .B1(new_n885), .B2(new_n518), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n907), .A2(new_n705), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n518), .A2(new_n937), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n706), .A2(new_n599), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n915), .B2(new_n941), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n938), .A2(new_n939), .A3(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(G148gat), .ZN(new_n944));
  OAI21_X1  g743(.A(KEYINPUT59), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n705), .B(new_n907), .C1(new_n908), .C2(new_n916), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n944), .A2(KEYINPUT59), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n947), .B1(new_n946), .B2(new_n948), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n945), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n927), .A2(new_n944), .A3(new_n705), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1345gat));
  NAND3_X1  g752(.A1(new_n922), .A2(new_n743), .A3(new_n907), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(G155gat), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n731), .A2(new_n335), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n926), .B2(new_n956), .ZN(G1346gat));
  NAND4_X1  g756(.A1(new_n922), .A2(G162gat), .A3(new_n678), .A4(new_n907), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n336), .B1(new_n926), .B2(new_n677), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n958), .A2(new_n959), .ZN(G1347gat));
  AOI21_X1  g759(.A(new_n735), .B1(new_n878), .B2(new_n879), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n519), .A2(new_n463), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(G169gat), .B1(new_n963), .B2(new_n746), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n786), .A2(new_n464), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n965), .A2(new_n764), .ZN(new_n966));
  AND4_X1   g765(.A1(KEYINPUT124), .A2(new_n885), .A3(new_n396), .A4(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(KEYINPUT124), .B1(new_n880), .B2(new_n966), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n599), .A2(new_n250), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n964), .B1(new_n969), .B2(new_n970), .ZN(G1348gat));
  NAND3_X1  g770(.A1(new_n963), .A2(new_n251), .A3(new_n705), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n967), .A2(new_n968), .A3(new_n782), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n972), .B1(new_n973), .B2(new_n251), .ZN(G1349gat));
  AOI21_X1  g773(.A(new_n227), .B1(new_n969), .B2(new_n743), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n961), .A2(new_n262), .A3(new_n731), .A4(new_n962), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n976), .B(new_n977), .ZN(new_n978));
  OAI21_X1  g777(.A(KEYINPUT60), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n976), .B(KEYINPUT125), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT60), .ZN(new_n981));
  NOR3_X1   g780(.A1(new_n967), .A2(new_n968), .A3(new_n847), .ZN(new_n982));
  OAI211_X1 g781(.A(new_n980), .B(new_n981), .C1(new_n227), .C2(new_n982), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n979), .A2(new_n983), .ZN(G1350gat));
  NAND3_X1  g783(.A1(new_n963), .A2(new_n226), .A3(new_n678), .ZN(new_n985));
  AOI211_X1 g784(.A(KEYINPUT61), .B(new_n229), .C1(new_n969), .C2(new_n678), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT61), .ZN(new_n987));
  INV_X1    g786(.A(new_n968), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n880), .A2(KEYINPUT124), .A3(new_n966), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n988), .A2(new_n678), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n987), .B1(new_n990), .B2(G190gat), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n985), .B1(new_n986), .B2(new_n991), .ZN(G1351gat));
  NOR3_X1   g791(.A1(new_n721), .A2(new_n464), .A3(new_n396), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n961), .A2(new_n993), .ZN(new_n994));
  NOR3_X1   g793(.A1(new_n994), .A2(G197gat), .A3(new_n747), .ZN(new_n995));
  XOR2_X1   g794(.A(new_n995), .B(KEYINPUT126), .Z(new_n996));
  NOR2_X1   g795(.A1(new_n938), .A2(new_n942), .ZN(new_n997));
  INV_X1    g796(.A(new_n965), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n997), .A2(new_n722), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g798(.A(G197gat), .B1(new_n999), .B2(new_n599), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n996), .A2(new_n1000), .ZN(G1352gat));
  NOR2_X1   g800(.A1(new_n782), .A2(G204gat), .ZN(new_n1002));
  INV_X1    g801(.A(new_n1002), .ZN(new_n1003));
  OR3_X1    g802(.A1(new_n994), .A2(KEYINPUT127), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g803(.A(KEYINPUT127), .B1(new_n994), .B2(new_n1003), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT62), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g807(.A(G204gat), .B1(new_n999), .B2(new_n782), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n1004), .A2(KEYINPUT62), .A3(new_n1005), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(G1353gat));
  OR3_X1    g810(.A1(new_n994), .A2(G211gat), .A3(new_n638), .ZN(new_n1012));
  NAND4_X1  g811(.A1(new_n997), .A2(new_n722), .A3(new_n731), .A4(new_n998), .ZN(new_n1013));
  AND3_X1   g812(.A1(new_n1013), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1014));
  AOI21_X1  g813(.A(KEYINPUT63), .B1(new_n1013), .B2(G211gat), .ZN(new_n1015));
  OAI21_X1  g814(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(G1354gat));
  OAI21_X1  g815(.A(G218gat), .B1(new_n999), .B2(new_n677), .ZN(new_n1017));
  OR2_X1    g816(.A1(new_n677), .A2(G218gat), .ZN(new_n1018));
  OAI21_X1  g817(.A(new_n1017), .B1(new_n994), .B2(new_n1018), .ZN(G1355gat));
endmodule


