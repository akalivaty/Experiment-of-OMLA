//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 1 1 0 0 0 1 0 1 1 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G13), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  AND2_X1   g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G20), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n202), .A2(G50), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G58), .A2(G232), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n222));
  AND4_X1   g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G68), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(KEYINPUT64), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT64), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G68), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G238), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n210), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(KEYINPUT1), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n215), .B1(new_n217), .B2(new_n218), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n230), .A2(new_n231), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT65), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n232), .A2(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G226), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G1), .A2(G13), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n209), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G150), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  OAI22_X1  g0059(.A1(new_n255), .A2(new_n256), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G50), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n209), .B1(new_n201), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n254), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT68), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g0065(.A(KEYINPUT68), .B(new_n254), .C1(new_n260), .C2(new_n262), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(new_n254), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n261), .B1(new_n208), .B2(G20), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n269), .A2(new_n270), .B1(new_n261), .B2(new_n268), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n265), .A2(new_n266), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(G1), .A3(G13), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(new_n277), .A3(G274), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n279), .B1(G226), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT3), .ZN(new_n285));
  INV_X1    g0085(.A(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  AOI21_X1  g0088(.A(G1698), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G222), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT3), .B(G33), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G223), .A3(G1698), .ZN(new_n292));
  AND2_X1   g0092(.A1(KEYINPUT3), .A2(G33), .ZN(new_n293));
  NOR2_X1   g0093(.A1(KEYINPUT3), .A2(G33), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G77), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n290), .A2(new_n292), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n277), .B1(new_n297), .B2(KEYINPUT67), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT67), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n290), .A2(new_n299), .A3(new_n292), .A4(new_n296), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n284), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n272), .B1(new_n301), .B2(G169), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n297), .A2(KEYINPUT67), .ZN(new_n303));
  INV_X1    g0103(.A(new_n277), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n303), .A2(new_n304), .A3(new_n300), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n283), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n306), .A2(G179), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(G200), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n301), .A2(G190), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT9), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n272), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n265), .A2(KEYINPUT9), .A3(new_n266), .A4(new_n271), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n309), .A2(new_n310), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT10), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n312), .A2(new_n313), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT10), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n316), .A2(new_n317), .A3(new_n310), .A4(new_n309), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n308), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n254), .ZN(new_n320));
  INV_X1    g0120(.A(new_n255), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n321), .A2(new_n258), .B1(G20), .B2(G77), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT15), .B(G87), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n323), .A2(new_n256), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n320), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n269), .ZN(new_n326));
  OAI21_X1  g0126(.A(G77), .B1(new_n209), .B2(G1), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n326), .A2(new_n327), .B1(G77), .B2(new_n267), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G244), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n278), .B1(new_n330), .B2(new_n281), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n291), .A2(G238), .A3(G1698), .ZN(new_n332));
  INV_X1    g0132(.A(G1698), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n291), .A2(G232), .A3(new_n333), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n332), .B(new_n334), .C1(new_n205), .C2(new_n291), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n331), .B1(new_n335), .B2(new_n304), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n329), .B(new_n338), .C1(G169), .C2(new_n336), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n336), .A2(G190), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n325), .A2(new_n328), .ZN(new_n341));
  INV_X1    g0141(.A(G200), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n340), .B(new_n341), .C1(new_n342), .C2(new_n336), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n319), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT69), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n319), .A2(KEYINPUT69), .A3(new_n344), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n258), .A2(G50), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT71), .ZN(new_n351));
  INV_X1    g0151(.A(G77), .ZN(new_n352));
  OAI22_X1  g0152(.A1(new_n228), .A2(new_n209), .B1(new_n352), .B2(new_n256), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n254), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT11), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n228), .B2(new_n267), .ZN(new_n358));
  OR3_X1    g0158(.A1(new_n267), .A2(KEYINPUT12), .A3(G68), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n224), .B1(new_n208), .B2(G20), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n358), .A2(new_n359), .B1(new_n269), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n354), .B2(new_n355), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n356), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n279), .B1(G238), .B2(new_n282), .ZN(new_n364));
  OAI211_X1 g0164(.A(G232), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n365));
  OAI211_X1 g0165(.A(G226), .B(new_n333), .C1(new_n293), .C2(new_n294), .ZN(new_n366));
  NAND2_X1  g0166(.A1(G33), .A2(G97), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT70), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n368), .A2(new_n369), .A3(new_n304), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n369), .B1(new_n368), .B2(new_n304), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n364), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT13), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT13), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n374), .B(new_n364), .C1(new_n370), .C2(new_n371), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G190), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n363), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n342), .B1(new_n373), .B2(new_n375), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n368), .A2(new_n304), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT70), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n368), .A2(new_n369), .A3(new_n304), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n374), .B1(new_n384), .B2(new_n364), .ZN(new_n385));
  INV_X1    g0185(.A(new_n375), .ZN(new_n386));
  OAI21_X1  g0186(.A(G169), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT14), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n373), .A2(G179), .A3(new_n375), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT14), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n390), .B(G169), .C1(new_n385), .C2(new_n386), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n363), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n380), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  INV_X1    g0195(.A(G159), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n259), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n201), .B1(new_n228), .B2(G58), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n398), .B1(new_n399), .B2(new_n209), .ZN(new_n400));
  XNOR2_X1  g0200(.A(KEYINPUT64), .B(G68), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n287), .A2(new_n209), .A3(new_n288), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n287), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n288), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n401), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n395), .B1(new_n400), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT7), .B1(new_n295), .B2(new_n209), .ZN(new_n408));
  INV_X1    g0208(.A(new_n405), .ZN(new_n409));
  OAI21_X1  g0209(.A(G68), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(G58), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n202), .B1(new_n401), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n397), .B1(new_n412), .B2(G20), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n410), .A2(new_n413), .A3(KEYINPUT16), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n407), .A2(new_n414), .A3(new_n254), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n255), .B1(new_n208), .B2(G20), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n416), .A2(new_n269), .B1(new_n268), .B2(new_n255), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  OAI211_X1 g0218(.A(G223), .B(new_n333), .C1(new_n293), .C2(new_n294), .ZN(new_n419));
  OAI211_X1 g0219(.A(G226), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G87), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n304), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n277), .A2(G232), .A3(new_n280), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n278), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT73), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT73), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n278), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n423), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G169), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n423), .A2(new_n426), .A3(G179), .A4(new_n428), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n418), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT18), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n429), .A2(G200), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n423), .A2(new_n426), .A3(G190), .A4(new_n428), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n437), .A2(KEYINPUT17), .A3(new_n415), .A4(new_n417), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n415), .A2(new_n417), .B1(new_n430), .B2(new_n431), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT18), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n415), .A2(new_n417), .A3(new_n436), .A4(new_n435), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT17), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n434), .A2(new_n438), .A3(new_n441), .A4(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n349), .A2(new_n394), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT21), .ZN(new_n448));
  OAI211_X1 g0248(.A(G257), .B(new_n333), .C1(new_n293), .C2(new_n294), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT78), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT78), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n291), .A2(new_n451), .A3(G257), .A4(new_n333), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(G264), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n287), .A2(G303), .A3(new_n288), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n277), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g0258(.A(KEYINPUT5), .B(G41), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n274), .A2(G1), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n459), .A2(new_n460), .B1(new_n216), .B2(new_n276), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G270), .ZN(new_n462));
  AND2_X1   g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  NOR2_X1   g0263(.A1(KEYINPUT5), .A2(G41), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g0265(.A1(G33), .A2(G41), .ZN(new_n466));
  OAI21_X1  g0266(.A(G274), .B1(new_n466), .B2(new_n253), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT75), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n208), .A2(G45), .ZN(new_n470));
  OR2_X1    g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  NAND2_X1  g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G274), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n474), .B1(new_n216), .B2(new_n276), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT75), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n462), .B1(new_n469), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n458), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G116), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n252), .A2(new_n253), .B1(G20), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G283), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n481), .B(new_n209), .C1(G33), .C2(new_n204), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n480), .A2(KEYINPUT20), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT20), .B1(new_n480), .B2(new_n482), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n267), .A2(G116), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n208), .A2(G33), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n320), .A2(new_n267), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n488), .B1(new_n490), .B2(new_n479), .ZN(new_n491));
  OAI21_X1  g0291(.A(G169), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n448), .B1(new_n478), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT80), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT80), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n495), .B(new_n448), .C1(new_n478), .C2(new_n492), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n486), .A2(new_n491), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n468), .B1(new_n465), .B2(new_n467), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n475), .A2(KEYINPUT75), .A3(new_n459), .A4(new_n460), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n501), .A2(G179), .A3(new_n462), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n498), .A2(new_n502), .A3(new_n458), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n499), .A2(new_n500), .B1(new_n461), .B2(G270), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n456), .B1(new_n452), .B2(new_n450), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n504), .B1(new_n505), .B2(new_n277), .ZN(new_n506));
  INV_X1    g0306(.A(G169), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n480), .A2(new_n482), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT20), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n483), .ZN(new_n511));
  AND4_X1   g0311(.A1(new_n253), .A2(new_n267), .A3(new_n252), .A4(new_n489), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n487), .B1(new_n512), .B2(G116), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n507), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n506), .A2(KEYINPUT21), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT79), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n506), .A2(new_n514), .A3(KEYINPUT79), .A4(KEYINPUT21), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n503), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n506), .A2(G200), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n520), .B(new_n498), .C1(new_n377), .C2(new_n506), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n497), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(G238), .B(new_n333), .C1(new_n293), .C2(new_n294), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G116), .ZN(new_n524));
  AND2_X1   g0324(.A1(G244), .A2(G1698), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n293), .B2(new_n294), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT76), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n523), .A2(new_n526), .A3(KEYINPUT76), .A4(new_n524), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(new_n304), .A3(new_n530), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n470), .A2(G250), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n277), .A2(new_n532), .B1(new_n475), .B2(new_n460), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n291), .A2(new_n209), .A3(G68), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT19), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n209), .B1(new_n367), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(G87), .B2(new_n206), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n536), .B1(new_n256), .B2(new_n204), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n540), .A2(new_n254), .B1(new_n268), .B2(new_n323), .ZN(new_n541));
  INV_X1    g0341(.A(new_n323), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n512), .A2(new_n542), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n534), .A2(new_n507), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n533), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n277), .B1(new_n527), .B2(new_n528), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(new_n530), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT77), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(new_n548), .A3(new_n337), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n531), .A2(new_n337), .A3(new_n533), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT77), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n544), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(G250), .B(new_n333), .C1(new_n293), .C2(new_n294), .ZN(new_n553));
  OAI211_X1 g0353(.A(G257), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G294), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(new_n304), .B1(new_n461), .B2(G264), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n557), .A2(new_n337), .A3(new_n501), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n501), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n507), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n209), .B(G87), .C1(new_n293), .C2(new_n294), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT22), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT22), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n291), .A2(new_n563), .A3(new_n209), .A4(G87), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n209), .A2(KEYINPUT23), .A3(G107), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT23), .ZN(new_n567));
  OAI22_X1  g0367(.A1(new_n566), .A2(KEYINPUT81), .B1(new_n567), .B2(new_n205), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n205), .A3(G20), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT81), .ZN(new_n570));
  AOI21_X1  g0370(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n571));
  OAI22_X1  g0371(.A1(new_n569), .A2(new_n570), .B1(new_n571), .B2(G20), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n565), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT24), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT24), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n565), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n320), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  XOR2_X1   g0378(.A(KEYINPUT82), .B(KEYINPUT25), .Z(new_n579));
  NOR2_X1   g0379(.A1(new_n267), .A2(G107), .ZN(new_n580));
  XNOR2_X1  g0380(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n490), .A2(new_n205), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n558), .B(new_n560), .C1(new_n578), .C2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n534), .A2(G200), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n512), .A2(G87), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n541), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n586), .B(new_n589), .C1(new_n377), .C2(new_n534), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n552), .A2(new_n585), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(G107), .B1(new_n408), .B2(new_n409), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n205), .A2(KEYINPUT6), .A3(G97), .ZN(new_n593));
  XOR2_X1   g0393(.A(G97), .B(G107), .Z(new_n594));
  OAI21_X1  g0394(.A(new_n593), .B1(new_n594), .B2(KEYINPUT6), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G20), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n258), .A2(G77), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n592), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n254), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n267), .A2(G97), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n512), .B2(G97), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(G244), .B(new_n333), .C1(new_n293), .C2(new_n294), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT4), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n330), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n291), .A2(new_n333), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n605), .A2(new_n481), .A3(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(G250), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT74), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT74), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n291), .A2(new_n611), .A3(G250), .A4(G1698), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n304), .B1(new_n608), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n499), .A2(new_n500), .B1(new_n461), .B2(G257), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n614), .A2(G179), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n507), .B1(new_n614), .B2(new_n615), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n602), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n565), .A2(new_n573), .A3(new_n576), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n576), .B1(new_n565), .B2(new_n573), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n254), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n559), .A2(G190), .ZN(new_n622));
  AOI21_X1  g0422(.A(G200), .B1(new_n557), .B2(new_n501), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n621), .B(new_n583), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n601), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(new_n598), .B2(new_n254), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n614), .A2(G190), .A3(new_n615), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n461), .A2(G257), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(new_n469), .B2(new_n476), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n289), .A2(new_n606), .B1(G33), .B2(G283), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n630), .A2(new_n605), .A3(new_n610), .A4(new_n612), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n629), .B1(new_n304), .B2(new_n631), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n626), .B(new_n627), .C1(new_n632), .C2(new_n342), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n618), .A2(new_n624), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n591), .A2(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n447), .A2(new_n522), .A3(new_n635), .ZN(G372));
  NAND2_X1  g0436(.A1(new_n315), .A2(new_n318), .ZN(new_n637));
  INV_X1    g0437(.A(new_n380), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n438), .A2(new_n444), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n391), .A2(new_n389), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n390), .B1(new_n376), .B2(G169), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n393), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n640), .B1(new_n339), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n439), .B(KEYINPUT18), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n637), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n308), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n447), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n618), .A2(new_n633), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n588), .B1(G190), .B2(new_n547), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n586), .A2(new_n652), .B1(new_n544), .B2(new_n550), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n651), .A2(KEYINPUT83), .A3(new_n624), .A4(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT83), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n544), .A2(new_n550), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n590), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n655), .B1(new_n634), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n497), .A2(new_n519), .A3(new_n585), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n654), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT84), .B1(new_n616), .B2(new_n617), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT84), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n614), .A2(G179), .A3(new_n615), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n662), .B(new_n663), .C1(new_n632), .C2(new_n507), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n661), .A2(new_n602), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT85), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n661), .A2(new_n664), .A3(KEYINPUT85), .A4(new_n602), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n667), .A2(new_n668), .A3(new_n653), .A4(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n656), .ZN(new_n671));
  INV_X1    g0471(.A(new_n617), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n626), .B1(new_n672), .B2(new_n663), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n673), .A2(new_n552), .A3(new_n590), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n671), .B1(new_n674), .B2(KEYINPUT26), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n660), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n649), .B1(new_n650), .B2(new_n677), .ZN(G369));
  INV_X1    g0478(.A(G330), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n498), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT86), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n497), .A2(new_n519), .A3(new_n521), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT87), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n690), .B2(new_n689), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n497), .A2(new_n519), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n688), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n679), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n685), .B1(new_n578), .B2(new_n584), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n585), .A2(new_n624), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n585), .A2(new_n686), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT88), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(KEYINPUT88), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n585), .A2(new_n685), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n685), .B1(new_n497), .B2(new_n519), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n705), .B1(new_n706), .B2(new_n697), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n704), .A2(new_n707), .ZN(G399));
  NOR2_X1   g0508(.A1(new_n212), .A2(G41), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G1), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n218), .B2(new_n710), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n556), .A2(new_n304), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n461), .A2(G264), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n502), .A2(new_n458), .A3(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(KEYINPUT30), .A3(new_n632), .A4(new_n547), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n453), .A2(new_n457), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n304), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n722), .A2(G179), .A3(new_n504), .A4(new_n557), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n614), .A2(new_n531), .A3(new_n615), .A4(new_n533), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n720), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n531), .A2(new_n533), .B1(new_n557), .B2(new_n501), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n614), .A2(new_n615), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n726), .A2(new_n337), .A3(new_n506), .A4(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n719), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n730));
  AOI21_X1  g0530(.A(KEYINPUT31), .B1(new_n729), .B2(new_n685), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n522), .A2(new_n635), .A3(new_n686), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n679), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n686), .B1(new_n660), .B2(new_n676), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n738), .A2(KEYINPUT29), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n657), .B1(new_n666), .B2(new_n665), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(KEYINPUT26), .A3(new_n669), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT89), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n742), .B1(new_n674), .B2(new_n668), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n740), .A2(new_n742), .A3(KEYINPUT26), .A4(new_n669), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n634), .A2(new_n657), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n671), .B1(new_n746), .B2(new_n659), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n744), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(KEYINPUT29), .A3(new_n686), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n736), .B1(new_n739), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n714), .B1(new_n750), .B2(G1), .ZN(G364));
  NOR2_X1   g0551(.A1(new_n211), .A2(G20), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n208), .B1(new_n752), .B2(G45), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n709), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n213), .A2(new_n291), .ZN(new_n756));
  INV_X1    g0556(.A(G355), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n756), .A2(new_n757), .B1(G116), .B2(new_n213), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n247), .A2(new_n274), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n213), .A2(new_n295), .ZN(new_n760));
  INV_X1    g0560(.A(new_n218), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n760), .B1(new_n274), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n758), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n253), .B1(G20), .B2(new_n507), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT90), .Z(new_n769));
  OAI21_X1  g0569(.A(new_n755), .B1(new_n763), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n337), .A2(new_n342), .A3(G190), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G294), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n209), .A2(G179), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n775), .A2(G190), .A3(G200), .ZN(new_n776));
  INV_X1    g0576(.A(G303), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n773), .A2(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G190), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT92), .Z(new_n781));
  AND2_X1   g0581(.A1(new_n781), .A2(G329), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n209), .A2(new_n337), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n779), .ZN(new_n784));
  INV_X1    g0584(.A(G311), .ZN(new_n785));
  INV_X1    g0585(.A(G322), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n783), .A2(G190), .A3(new_n342), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n295), .B1(new_n784), .B2(new_n785), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n783), .A2(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G190), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  XOR2_X1   g0591(.A(KEYINPUT33), .B(G317), .Z(new_n792));
  NOR2_X1   g0592(.A1(new_n789), .A2(new_n377), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G326), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n791), .A2(new_n792), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OR3_X1    g0596(.A1(new_n782), .A2(new_n788), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n775), .A2(new_n377), .A3(G200), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n778), .B(new_n797), .C1(G283), .C2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n801), .A2(KEYINPUT93), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(KEYINPUT93), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n291), .B1(new_n787), .B2(new_n411), .ZN(new_n804));
  INV_X1    g0604(.A(G87), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n791), .A2(new_n224), .B1(new_n805), .B2(new_n776), .ZN(new_n806));
  INV_X1    g0606(.A(new_n784), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n804), .B(new_n806), .C1(G77), .C2(new_n807), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n772), .B(KEYINPUT91), .Z(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G97), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n793), .A2(G50), .B1(new_n799), .B2(G107), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n780), .A2(new_n396), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT32), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n808), .A2(new_n810), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n802), .A2(new_n803), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n770), .B1(new_n815), .B2(new_n767), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n692), .A2(new_n694), .ZN(new_n817));
  INV_X1    g0617(.A(new_n766), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n695), .A2(new_n755), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n817), .A2(G330), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(G396));
  INV_X1    g0622(.A(KEYINPUT95), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n329), .A2(new_n685), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n344), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n339), .A2(new_n343), .A3(new_n824), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(KEYINPUT95), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n686), .B(new_n828), .C1(new_n660), .C2(new_n676), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n339), .A2(new_n686), .ZN(new_n830));
  AND3_X1   g0630(.A1(new_n825), .A2(new_n830), .A3(new_n827), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n829), .B1(new_n738), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n736), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n755), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n834), .B2(new_n833), .ZN(new_n836));
  INV_X1    g0636(.A(new_n767), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n765), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n755), .B1(G77), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n787), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n840), .A2(G143), .B1(new_n807), .B2(G159), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n841), .B1(new_n794), .B2(new_n842), .C1(new_n257), .C2(new_n791), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT34), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n781), .A2(G132), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n773), .A2(new_n411), .B1(new_n776), .B2(new_n261), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n295), .B(new_n847), .C1(G68), .C2(new_n799), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n843), .A2(new_n844), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT94), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n295), .B1(new_n784), .B2(new_n479), .C1(new_n774), .C2(new_n787), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n781), .B2(G311), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n790), .A2(G283), .B1(new_n793), .B2(G303), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n798), .A2(new_n805), .ZN(new_n856));
  INV_X1    g0656(.A(new_n776), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(G107), .B2(new_n857), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n854), .A2(new_n810), .A3(new_n855), .A4(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n851), .B1(new_n852), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n852), .B2(new_n859), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n839), .B1(new_n861), .B2(new_n767), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n832), .B2(new_n765), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n836), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(G384));
  NAND3_X1  g0665(.A1(new_n739), .A2(new_n447), .A3(new_n749), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n649), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT100), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n224), .B1(new_n404), .B2(new_n405), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n395), .B1(new_n400), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n870), .A2(new_n414), .A3(new_n254), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n417), .ZN(new_n872));
  INV_X1    g0672(.A(new_n683), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n445), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n418), .A2(new_n873), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n433), .A2(new_n877), .A3(new_n878), .A4(new_n442), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n872), .A2(new_n432), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n880), .A2(new_n874), .A3(new_n442), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n879), .B1(new_n881), .B2(new_n878), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n876), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n876), .A2(new_n882), .A3(KEYINPUT38), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n885), .A2(KEYINPUT39), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n433), .A2(new_n877), .A3(new_n442), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n683), .B1(new_n415), .B2(new_n417), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT99), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT37), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n888), .B(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n877), .B1(new_n645), .B2(new_n639), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n884), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT39), .B1(new_n894), .B2(new_n886), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n887), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n392), .A2(new_n393), .A3(new_n686), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n645), .A2(new_n873), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n393), .A2(new_n685), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n643), .A2(new_n638), .A3(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n393), .B(new_n685), .C1(new_n392), .C2(new_n380), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n339), .A2(new_n685), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT97), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n905), .B1(new_n829), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n885), .A2(new_n886), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n900), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT98), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n899), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI211_X1 g0712(.A(KEYINPUT98), .B(new_n900), .C1(new_n908), .C2(new_n909), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n868), .B(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n878), .B1(new_n877), .B2(KEYINPUT99), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(new_n888), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n445), .A2(new_n889), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT38), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n876), .A2(new_n882), .A3(KEYINPUT38), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n904), .A2(new_n734), .A3(new_n832), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT40), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n904), .A2(new_n734), .A3(new_n832), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT40), .B1(new_n885), .B2(new_n886), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n447), .B2(new_n734), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n831), .B1(new_n732), .B2(new_n733), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n929), .B(new_n904), .C1(new_n919), .C2(new_n920), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n930), .A2(KEYINPUT40), .B1(new_n924), .B2(new_n925), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n931), .A2(new_n650), .A3(new_n735), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n928), .A2(new_n932), .A3(new_n679), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n915), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n915), .A2(new_n933), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n934), .B(new_n935), .C1(new_n208), .C2(new_n752), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n595), .A2(KEYINPUT35), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n217), .A2(new_n479), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n595), .B2(KEYINPUT35), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT96), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n940), .B2(new_n939), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT36), .Z(new_n943));
  AOI211_X1 g0743(.A(new_n352), .B(new_n218), .C1(new_n228), .C2(G58), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n224), .A2(G50), .ZN(new_n945));
  OAI211_X1 g0745(.A(G1), .B(new_n211), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n936), .A2(new_n943), .A3(new_n946), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT101), .Z(G367));
  OAI221_X1 g0748(.A(new_n768), .B1(new_n213), .B2(new_n323), .C1(new_n243), .C2(new_n760), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n949), .A2(new_n755), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n588), .A2(new_n685), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n653), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n656), .B2(new_n951), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n787), .A2(new_n257), .B1(new_n784), .B2(new_n261), .ZN(new_n954));
  INV_X1    g0754(.A(new_n780), .ZN(new_n955));
  AOI211_X1 g0755(.A(new_n295), .B(new_n954), .C1(G137), .C2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n809), .A2(G68), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n790), .A2(G159), .B1(new_n793), .B2(G143), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n798), .A2(new_n352), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(G58), .B2(new_n857), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n956), .A2(new_n957), .A3(new_n958), .A4(new_n960), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n793), .A2(G311), .B1(G107), .B2(new_n772), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n962), .B1(new_n204), .B2(new_n798), .C1(new_n774), .C2(new_n791), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n840), .A2(G303), .B1(new_n955), .B2(G317), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT46), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n776), .B2(new_n479), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n857), .A2(KEYINPUT46), .A3(G116), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n291), .B1(new_n807), .B2(G283), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n964), .A2(new_n966), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n961), .B1(new_n963), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT47), .Z(new_n971));
  OAI221_X1 g0771(.A(new_n950), .B1(new_n953), .B2(new_n818), .C1(new_n837), .C2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n665), .A2(new_n686), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n651), .B1(new_n626), .B2(new_n686), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n706), .A2(new_n697), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT42), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n618), .B1(new_n976), .B2(new_n585), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n686), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n979), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT102), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n979), .A2(new_n982), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n953), .B(KEYINPUT43), .Z(new_n986));
  AOI22_X1  g0786(.A1(new_n983), .A2(new_n984), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n979), .A2(KEYINPUT102), .A3(new_n980), .A4(new_n982), .ZN(new_n988));
  AOI21_X1  g0788(.A(KEYINPUT103), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n983), .A2(new_n984), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n985), .A2(new_n986), .ZN(new_n991));
  AND4_X1   g0791(.A1(KEYINPUT103), .A2(new_n990), .A3(new_n988), .A4(new_n991), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n989), .A2(new_n992), .B1(new_n704), .B2(new_n976), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n987), .A2(new_n988), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT103), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n704), .A2(new_n976), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n987), .A2(KEYINPUT103), .A3(new_n988), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n993), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT104), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n701), .A2(new_n1001), .A3(new_n702), .ZN(new_n1002));
  AND2_X1   g0802(.A1(new_n707), .A2(new_n975), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1003), .A2(KEYINPUT45), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n707), .A2(new_n975), .A3(KEYINPUT45), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT44), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n707), .B2(new_n975), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n707), .A2(new_n975), .A3(new_n1006), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n1004), .A2(new_n1005), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1002), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1010), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1012), .A2(new_n1001), .A3(new_n701), .A4(new_n702), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n977), .B1(new_n699), .B2(new_n706), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n695), .B(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n750), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n709), .B(KEYINPUT41), .Z(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n754), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n972), .B1(new_n1000), .B2(new_n1021), .ZN(G387));
  OR2_X1    g0822(.A1(new_n699), .A2(new_n818), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n756), .A2(new_n711), .B1(G107), .B2(new_n213), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n240), .A2(new_n274), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n711), .ZN(new_n1026));
  AOI211_X1 g0826(.A(G45), .B(new_n1026), .C1(G68), .C2(G77), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n255), .A2(G50), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT50), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n760), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1024), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n755), .B1(new_n1031), .B2(new_n769), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n787), .A2(new_n261), .B1(new_n780), .B2(new_n257), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n295), .B(new_n1033), .C1(G68), .C2(new_n807), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n809), .A2(new_n542), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n790), .A2(new_n321), .B1(new_n799), .B2(G97), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n793), .A2(G159), .B1(new_n857), .B2(G77), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(G283), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n773), .A2(new_n1039), .B1(new_n776), .B2(new_n774), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n840), .A2(G317), .B1(new_n807), .B2(G303), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n794), .B2(new_n786), .C1(new_n785), .C2(new_n791), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT48), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1040), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n1043), .B2(new_n1042), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT49), .Z(new_n1046));
  OAI221_X1 g0846(.A(new_n295), .B1(new_n780), .B2(new_n795), .C1(new_n479), .C2(new_n798), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1038), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1032), .B1(new_n1048), .B2(new_n767), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1016), .A2(new_n754), .B1(new_n1023), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n750), .A2(new_n1016), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n709), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n750), .A2(new_n1016), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1050), .B1(new_n1052), .B2(new_n1053), .ZN(G393));
  XNOR2_X1  g0854(.A(new_n703), .B(new_n1010), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1052), .A2(new_n753), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n768), .B1(new_n204), .B2(new_n213), .C1(new_n250), .C2(new_n760), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n755), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n809), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1060), .A2(new_n352), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT51), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n794), .A2(new_n257), .B1(new_n396), .B2(new_n787), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n295), .B1(new_n955), .B2(G143), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n255), .B2(new_n784), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n856), .B1(G50), .B2(new_n790), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n401), .C2(new_n776), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G317), .A2(new_n793), .B1(new_n840), .B2(G311), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT52), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n791), .A2(new_n777), .B1(new_n798), .B2(new_n205), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n295), .B1(new_n780), .B2(new_n786), .C1(new_n774), .C2(new_n784), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n773), .A2(new_n479), .B1(new_n776), .B2(new_n1039), .ZN(new_n1075));
  OR3_X1    g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n1065), .A2(new_n1070), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1059), .B1(new_n1077), .B2(new_n767), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n975), .B2(new_n818), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1014), .A2(new_n709), .A3(new_n750), .A4(new_n1016), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1057), .A2(new_n1079), .A3(new_n1080), .ZN(G390));
  NAND3_X1  g0881(.A1(new_n929), .A2(G330), .A3(new_n904), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n908), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n896), .B1(new_n1084), .B2(new_n897), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n897), .B1(new_n919), .B2(new_n920), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n748), .A2(new_n686), .A3(new_n828), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n906), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1086), .B1(new_n1088), .B2(new_n904), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1083), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n885), .A2(KEYINPUT39), .A3(new_n886), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n921), .B2(KEYINPUT39), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n908), .B2(new_n898), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n905), .B1(new_n1087), .B2(new_n906), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1093), .B(new_n1082), .C1(new_n1094), .C2(new_n1086), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1090), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n754), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n755), .B1(new_n321), .B2(new_n838), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n794), .A2(new_n1039), .B1(new_n776), .B2(new_n805), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n791), .A2(new_n205), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n295), .B1(new_n784), .B2(new_n204), .C1(new_n479), .C2(new_n787), .ZN(new_n1101));
  NOR4_X1   g0901(.A1(new_n1061), .A2(new_n1099), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n781), .A2(G294), .B1(G68), .B2(new_n799), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT107), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT108), .ZN(new_n1106));
  INV_X1    g0906(.A(G132), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n291), .B1(new_n787), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(G128), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n794), .A2(new_n1109), .B1(new_n798), .B2(new_n261), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1108), .B(new_n1110), .C1(G137), .C2(new_n790), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(KEYINPUT54), .B(G143), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT106), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n781), .A2(G125), .B1(new_n807), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n776), .A2(new_n257), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT53), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n809), .A2(G159), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1111), .A2(new_n1114), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(KEYINPUT109), .B1(new_n1106), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1119), .A2(new_n837), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1106), .A2(KEYINPUT109), .A3(new_n1118), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1098), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n896), .B2(new_n765), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1097), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n447), .A2(new_n736), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n866), .A2(new_n649), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n929), .A2(G330), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n905), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n1082), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n829), .A2(new_n907), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n1088), .B2(new_n1129), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1126), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT105), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n1135), .A2(new_n1096), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n710), .B1(new_n1135), .B2(new_n1096), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1124), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(G378));
  INV_X1    g0939(.A(KEYINPUT116), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT115), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n637), .A2(new_n648), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n272), .A2(new_n873), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1144), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n319), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1142), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n319), .A2(new_n1146), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1144), .B(new_n308), .C1(new_n315), .C2(new_n318), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1142), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1141), .B1(new_n1148), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1145), .A2(new_n1147), .A3(new_n1142), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1151), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(new_n1155), .A3(KEYINPUT115), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n927), .A2(new_n1140), .A3(G330), .A4(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1148), .A2(new_n1152), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n931), .B2(new_n679), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n679), .B1(new_n923), .B2(new_n926), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1140), .B1(new_n1162), .B2(new_n1157), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1161), .A2(new_n914), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n1166), .A2(new_n1163), .B1(new_n913), .B2(new_n912), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1090), .A2(new_n1095), .A3(new_n1132), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n1126), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT117), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT57), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1165), .A2(new_n1167), .B1(new_n1126), .B2(new_n1169), .ZN(new_n1175));
  OAI21_X1  g0975(.A(KEYINPUT117), .B1(new_n1175), .B2(KEYINPUT57), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n710), .B1(new_n1175), .B2(KEYINPUT57), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1174), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n755), .B1(G50), .B2(new_n838), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1157), .A2(new_n765), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n790), .A2(G97), .B1(new_n799), .B2(G58), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n957), .B(new_n1181), .C1(new_n479), .C2(new_n794), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n787), .A2(new_n205), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT110), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n781), .A2(G283), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n857), .A2(G77), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n295), .A2(new_n273), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n542), .B2(new_n807), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .A4(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1182), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1191), .A2(KEYINPUT58), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1187), .B(new_n261), .C1(G33), .C2(G41), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1194), .A2(KEYINPUT111), .B1(KEYINPUT58), .B2(new_n1191), .ZN(new_n1195));
  AOI211_X1 g0995(.A(G33), .B(G41), .C1(new_n955), .C2(G124), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n809), .A2(G150), .B1(G125), .B2(new_n793), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT113), .Z(new_n1198));
  NAND2_X1  g0998(.A1(new_n1113), .A2(new_n857), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1199), .A2(KEYINPUT112), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(KEYINPUT112), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n787), .A2(new_n1109), .B1(new_n784), .B2(new_n842), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G132), .B2(new_n790), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1198), .A2(new_n1200), .A3(new_n1201), .A4(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT59), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT114), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1196), .B1(new_n396), .B2(new_n798), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1195), .B1(KEYINPUT111), .B2(new_n1194), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1179), .B(new_n1180), .C1(new_n767), .C2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n1168), .B2(new_n754), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1178), .A2(new_n1211), .ZN(G375));
  OR2_X1    g1012(.A1(new_n1126), .A2(new_n1132), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1213), .A2(new_n1020), .A3(new_n1133), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1132), .A2(new_n754), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n755), .B1(G68), .B2(new_n838), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n396), .A2(new_n776), .B1(new_n784), .B2(new_n257), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n781), .B2(G128), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n291), .B1(new_n798), .B2(new_n411), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT118), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1218), .B(new_n1220), .C1(new_n261), .C2(new_n1060), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT119), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n794), .A2(new_n1107), .B1(new_n842), .B2(new_n787), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n790), .B2(new_n1113), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n794), .A2(new_n774), .B1(new_n776), .B2(new_n204), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n959), .B(new_n1226), .C1(G116), .C2(new_n790), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n781), .A2(G303), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n295), .B1(new_n787), .B2(new_n1039), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(G107), .B2(new_n807), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1227), .A2(new_n1035), .A3(new_n1228), .A4(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1225), .A2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1216), .B1(new_n1232), .B2(new_n767), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n904), .B2(new_n765), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1214), .A2(new_n1215), .A3(new_n1234), .ZN(G381));
  INV_X1    g1035(.A(G390), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(G393), .A2(G396), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(new_n864), .A3(new_n1237), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1238), .A2(G387), .A3(G381), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1239), .A2(new_n1138), .A3(new_n1211), .A4(new_n1178), .ZN(G407));
  NAND2_X1  g1040(.A1(new_n684), .A2(G213), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(G375), .A2(G378), .A3(new_n1241), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(KEYINPUT120), .ZN(new_n1243));
  AND2_X1   g1043(.A1(G407), .A2(G213), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(KEYINPUT121), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT121), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1243), .A2(new_n1247), .A3(new_n1244), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(G409));
  NAND3_X1  g1049(.A1(new_n1178), .A2(G378), .A3(new_n1211), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1211), .B1(new_n1019), .B2(new_n1171), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1138), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(KEYINPUT122), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT122), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1251), .A2(new_n1254), .A3(new_n1138), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1250), .A2(new_n1253), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1215), .A2(new_n1234), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT60), .ZN(new_n1258));
  OR3_X1    g1058(.A1(new_n1126), .A2(new_n1132), .A3(new_n1258), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1259), .A2(new_n709), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1133), .A2(KEYINPUT60), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1213), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1257), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1263), .B(new_n864), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1256), .A2(new_n1241), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT62), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1256), .A2(new_n1241), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1263), .B(G384), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n684), .A2(G213), .A3(G2897), .ZN(new_n1269));
  XOR2_X1   g1069(.A(new_n1269), .B(KEYINPUT124), .Z(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1268), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1264), .A2(new_n1270), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1267), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT61), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT62), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1256), .A2(new_n1277), .A3(new_n1241), .A4(new_n1264), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1266), .A2(new_n1275), .A3(new_n1276), .A4(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT125), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G387), .A2(new_n1236), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G390), .B(new_n972), .C1(new_n1000), .C2(new_n1021), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(G393), .B(G396), .ZN(new_n1283));
  AND4_X1   g1083(.A1(new_n1280), .A2(new_n1281), .A3(new_n1282), .A4(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(KEYINPUT125), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(new_n1285), .A2(new_n1283), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1279), .A2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1276), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1289), .B1(new_n1265), .B2(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1256), .A2(KEYINPUT63), .A3(new_n1241), .A4(new_n1264), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1267), .A2(KEYINPUT123), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1274), .B1(new_n1267), .B2(KEYINPUT123), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1291), .B(new_n1292), .C1(new_n1293), .C2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1288), .A2(new_n1295), .ZN(G405));
  AND3_X1   g1096(.A1(new_n1178), .A2(G378), .A3(new_n1211), .ZN(new_n1297));
  AOI21_X1  g1097(.A(G378), .B1(new_n1178), .B2(new_n1211), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1264), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT126), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1264), .B(KEYINPUT126), .C1(new_n1297), .C2(new_n1298), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(G375), .A2(new_n1138), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1304), .A2(new_n1250), .A3(new_n1268), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT127), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1304), .A2(KEYINPUT127), .A3(new_n1250), .A4(new_n1268), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1303), .A2(new_n1309), .A3(new_n1287), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1287), .B1(new_n1303), .B2(new_n1309), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(G402));
endmodule


