//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 0 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G78gat), .B(G106gat), .ZN(new_n204));
  XOR2_X1   g003(.A(G197gat), .B(G204gat), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(KEYINPUT71), .A2(G211gat), .ZN(new_n207));
  AND2_X1   g006(.A1(KEYINPUT71), .A2(G211gat), .ZN(new_n208));
  AND2_X1   g007(.A1(KEYINPUT72), .A2(G218gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(KEYINPUT72), .A2(G218gat), .ZN(new_n210));
  OAI22_X1  g009(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT73), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT22), .ZN(new_n213));
  AND3_X1   g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n212), .B1(new_n211), .B2(new_n213), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n206), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G211gat), .B(G218gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT74), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT29), .ZN(new_n221));
  INV_X1    g020(.A(G155gat), .ZN(new_n222));
  INV_X1    g021(.A(G162gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(G155gat), .A2(G162gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G141gat), .B(G148gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n226), .B1(KEYINPUT2), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G148gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(G141gat), .ZN(new_n230));
  XOR2_X1   g029(.A(KEYINPUT79), .B(G148gat), .Z(new_n231));
  AOI21_X1  g030(.A(new_n230), .B1(new_n231), .B2(G141gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT2), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n224), .B1(new_n233), .B2(new_n225), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n228), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n221), .B1(new_n235), .B2(KEYINPUT3), .ZN(new_n236));
  OR2_X1    g035(.A1(KEYINPUT71), .A2(G211gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(KEYINPUT71), .A2(G211gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT72), .ZN(new_n239));
  INV_X1    g038(.A(G218gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(KEYINPUT72), .A2(G218gat), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n237), .A2(new_n238), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT73), .B1(new_n243), .B2(KEYINPUT22), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n219), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n247), .A3(new_n206), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n220), .A2(new_n236), .A3(new_n248), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n216), .A2(new_n217), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT29), .B1(new_n216), .B2(new_n217), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT3), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n235), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n249), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G228gat), .ZN(new_n255));
  INV_X1    g054(.A(G233gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n247), .B1(new_n246), .B2(new_n206), .ZN(new_n260));
  AOI211_X1 g059(.A(new_n219), .B(new_n205), .C1(new_n244), .C2(new_n245), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n221), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT3), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n253), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT84), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n257), .ZN(new_n266));
  NOR3_X1   g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT29), .B1(new_n220), .B2(new_n248), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n235), .B1(new_n268), .B2(KEYINPUT3), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n260), .A2(new_n261), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n258), .B1(new_n270), .B2(new_n236), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT84), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n259), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(G22gat), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n265), .B1(new_n264), .B2(new_n266), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n269), .A2(new_n271), .A3(KEYINPUT84), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G22gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(new_n278), .A3(new_n259), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n204), .B1(new_n280), .B2(KEYINPUT83), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT83), .ZN(new_n282));
  INV_X1    g081(.A(new_n204), .ZN(new_n283));
  AOI211_X1 g082(.A(new_n282), .B(new_n283), .C1(new_n274), .C2(new_n279), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n203), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  AOI221_X4 g084(.A(G22gat), .B1(new_n254), .B2(new_n258), .C1(new_n275), .C2(new_n276), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n278), .B1(new_n277), .B2(new_n259), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT83), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(new_n283), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n280), .A2(KEYINPUT83), .A3(new_n204), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(new_n290), .A3(new_n202), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n253), .A2(new_n263), .ZN(new_n293));
  XOR2_X1   g092(.A(KEYINPUT67), .B(G113gat), .Z(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G120gat), .ZN(new_n295));
  INV_X1    g094(.A(G120gat), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n296), .A2(G113gat), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n297), .A2(KEYINPUT66), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(KEYINPUT66), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n295), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(G127gat), .B(G134gat), .Z(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(KEYINPUT1), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT1), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n296), .A2(G113gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n303), .B1(new_n297), .B2(new_n304), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n300), .A2(new_n302), .B1(new_n305), .B2(new_n301), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n235), .A2(KEYINPUT3), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(new_n253), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT4), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n306), .A2(new_n253), .A3(KEYINPUT4), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n309), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT39), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n306), .A2(new_n253), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n321), .A2(new_n310), .A3(KEYINPUT80), .ZN(new_n322));
  OR3_X1    g121(.A1(new_n306), .A2(new_n253), .A3(KEYINPUT80), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n324), .A2(KEYINPUT86), .A3(new_n315), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT86), .B1(new_n324), .B2(new_n315), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n319), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT40), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT87), .ZN(new_n329));
  XOR2_X1   g128(.A(G57gat), .B(G85gat), .Z(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(KEYINPUT82), .ZN(new_n331));
  XOR2_X1   g130(.A(KEYINPUT81), .B(KEYINPUT0), .Z(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G1gat), .B(G29gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n335), .B1(new_n317), .B2(new_n318), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n327), .A2(new_n329), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n322), .A2(new_n316), .A3(new_n323), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT5), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(new_n316), .B2(new_n314), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n314), .A2(new_n316), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT5), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n335), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n337), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n329), .B1(new_n327), .B2(new_n336), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT65), .ZN(new_n347));
  NAND2_X1  g146(.A1(G169gat), .A2(G176gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(G169gat), .A2(G176gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n348), .B1(new_n349), .B2(KEYINPUT23), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n351), .A2(G169gat), .A3(G176gat), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n347), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n354), .A2(KEYINPUT24), .ZN(new_n355));
  INV_X1    g154(.A(G183gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(G190gat), .ZN(new_n357));
  INV_X1    g156(.A(G190gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G183gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n355), .B1(new_n360), .B2(KEYINPUT24), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n349), .A2(KEYINPUT23), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n351), .B1(G169gat), .B2(G176gat), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n362), .A2(KEYINPUT65), .A3(new_n363), .A4(new_n348), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n353), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  XOR2_X1   g164(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n366));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n352), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT24), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n368), .B1(new_n357), .B2(new_n359), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT25), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n369), .A2(new_n370), .A3(new_n355), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n365), .A2(new_n366), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n349), .A2(KEYINPUT26), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT26), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n348), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n373), .B(new_n354), .C1(new_n375), .C2(new_n349), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT28), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT27), .B(G183gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n377), .B1(new_n379), .B2(G190gat), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n378), .A2(KEYINPUT28), .A3(new_n358), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n376), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n221), .B1(new_n372), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT75), .ZN(new_n384));
  NAND2_X1  g183(.A1(G226gat), .A2(G233gat), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n384), .B1(new_n383), .B2(new_n385), .ZN(new_n387));
  INV_X1    g186(.A(new_n385), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n388), .B1(new_n372), .B2(new_n382), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n220), .A2(new_n248), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n386), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n365), .A2(new_n366), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n371), .A2(new_n367), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n382), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n385), .B1(new_n395), .B2(KEYINPUT29), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n390), .B1(new_n396), .B2(new_n389), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT76), .B1(new_n392), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(KEYINPUT75), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n389), .A2(new_n390), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT76), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n396), .A2(new_n389), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n270), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G8gat), .B(G36gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  XOR2_X1   g208(.A(new_n409), .B(KEYINPUT77), .Z(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n398), .A2(new_n406), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n402), .A2(new_n405), .A3(new_n409), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n402), .A2(new_n405), .A3(KEYINPUT30), .A4(new_n409), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT78), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n416), .A2(new_n417), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n412), .B(new_n415), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT85), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n412), .A2(new_n415), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT85), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n416), .B(new_n417), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n346), .A2(new_n421), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n335), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n341), .B1(KEYINPUT5), .B2(new_n338), .ZN(new_n428));
  INV_X1    g227(.A(new_n342), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n343), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n340), .A2(KEYINPUT6), .A3(new_n335), .A4(new_n342), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n398), .A2(KEYINPUT37), .A3(new_n406), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT37), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n402), .A2(new_n437), .A3(new_n405), .ZN(new_n438));
  INV_X1    g237(.A(new_n409), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT38), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n437), .B1(new_n404), .B2(new_n390), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n399), .A2(new_n389), .A3(new_n270), .A4(new_n400), .ZN(new_n443));
  AOI211_X1 g242(.A(KEYINPUT38), .B(new_n410), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n438), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n435), .A2(new_n413), .A3(new_n441), .A4(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n292), .A2(new_n426), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n395), .A2(new_n307), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n306), .B1(new_n372), .B2(new_n382), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(G227gat), .A2(G233gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(KEYINPUT68), .A3(KEYINPUT34), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT68), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n448), .A2(new_n449), .B1(G227gat), .B2(G233gat), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT34), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n450), .A2(new_n456), .A3(new_n451), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT69), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT69), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n455), .A2(new_n461), .A3(new_n456), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT32), .B1(new_n450), .B2(new_n451), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT33), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n466), .B1(new_n450), .B2(new_n451), .ZN(new_n467));
  XOR2_X1   g266(.A(G15gat), .B(G43gat), .Z(new_n468));
  XNOR2_X1  g267(.A(G71gat), .B(G99gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n465), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n470), .ZN(new_n472));
  OAI221_X1 g271(.A(KEYINPUT32), .B1(new_n466), .B2(new_n472), .C1(new_n450), .C2(new_n451), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n464), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n458), .A2(new_n463), .A3(new_n471), .A4(new_n473), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT36), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT70), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n475), .A2(new_n478), .A3(new_n476), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n464), .A2(KEYINPUT70), .A3(new_n474), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n477), .B1(new_n481), .B2(KEYINPUT36), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n434), .A2(new_n422), .A3(new_n424), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n285), .A2(new_n484), .A3(new_n291), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n447), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n423), .B1(new_n422), .B2(new_n424), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n420), .A2(KEYINPUT85), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n434), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT88), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT89), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT90), .B(KEYINPUT35), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n475), .A2(KEYINPUT89), .A3(new_n476), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n497), .B1(new_n285), .B2(new_n291), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n425), .A2(new_n421), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(KEYINPUT88), .A3(new_n434), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n491), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT35), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n285), .A2(new_n291), .B1(new_n480), .B2(new_n479), .ZN(new_n503));
  INV_X1    g302(.A(new_n484), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n486), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G229gat), .A2(G233gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(KEYINPUT94), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(KEYINPUT13), .ZN(new_n509));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT16), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(G1gat), .ZN(new_n512));
  INV_X1    g311(.A(G1gat), .ZN(new_n513));
  INV_X1    g312(.A(G15gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n514), .A2(G22gat), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n278), .A2(G15gat), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(G8gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT92), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT92), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n518), .A2(new_n521), .A3(G8gat), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT93), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n512), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(G8gat), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n510), .B(KEYINPUT93), .C1(new_n511), .C2(G1gat), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n524), .A2(new_n525), .A3(new_n517), .A4(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n520), .A2(new_n522), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G36gat), .ZN(new_n529));
  AND2_X1   g328(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n530));
  NOR2_X1   g329(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(G29gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n533), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n537));
  XNOR2_X1  g336(.A(G43gat), .B(G50gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n537), .A2(new_n538), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OR3_X1    g340(.A1(new_n528), .A2(new_n541), .A3(KEYINPUT97), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT97), .B1(new_n528), .B2(new_n541), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n541), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT96), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n509), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n528), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n541), .A2(KEYINPUT17), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT17), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n551), .B1(new_n539), .B2(new_n540), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n549), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n508), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n554), .A3(new_n545), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT18), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n553), .A2(KEYINPUT18), .A3(new_n554), .A4(new_n545), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n548), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n548), .A2(KEYINPUT95), .A3(new_n558), .ZN(new_n560));
  XNOR2_X1  g359(.A(G113gat), .B(G141gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(G169gat), .B(G197gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(KEYINPUT91), .B(KEYINPUT11), .Z(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT12), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n559), .A2(new_n560), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n509), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n545), .B(KEYINPUT96), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n542), .A2(new_n543), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n558), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n574), .B(new_n557), .C1(KEYINPUT95), .C2(new_n566), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n568), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT106), .ZN(new_n577));
  XNOR2_X1  g376(.A(G183gat), .B(G211gat), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(G127gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT9), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT101), .ZN(new_n584));
  XOR2_X1   g383(.A(G57gat), .B(G64gat), .Z(new_n585));
  NOR2_X1   g384(.A1(new_n585), .A2(KEYINPUT100), .ZN(new_n586));
  INV_X1    g385(.A(G57gat), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n587), .A2(G64gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT100), .ZN(new_n589));
  INV_X1    g388(.A(new_n581), .ZN(new_n590));
  NOR2_X1   g389(.A1(G71gat), .A2(G78gat), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OR3_X1    g391(.A1(new_n584), .A2(new_n586), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT99), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n585), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n587), .A2(G64gat), .ZN(new_n596));
  OR3_X1    g395(.A1(new_n596), .A2(new_n588), .A3(new_n594), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n595), .A2(new_n583), .A3(new_n597), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n590), .A2(KEYINPUT98), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n590), .A2(KEYINPUT98), .ZN(new_n600));
  NOR3_X1   g399(.A1(new_n599), .A2(new_n600), .A3(new_n591), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n593), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  OAI211_X1 g403(.A(G231gat), .B(G233gat), .C1(new_n604), .C2(KEYINPUT21), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT21), .ZN(new_n606));
  NAND2_X1  g405(.A1(G231gat), .A2(G233gat), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n603), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n580), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n605), .A2(new_n580), .A3(new_n608), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n579), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT102), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G155gat), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n549), .B1(new_n603), .B2(new_n606), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n618), .A2(KEYINPUT103), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(KEYINPUT103), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n610), .A2(new_n579), .A3(new_n611), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n619), .A2(new_n620), .A3(new_n617), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n613), .A2(new_n622), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n623), .ZN(new_n626));
  INV_X1    g425(.A(new_n624), .ZN(new_n627));
  OAI22_X1  g426(.A1(new_n626), .A2(new_n612), .B1(new_n627), .B2(new_n621), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(KEYINPUT104), .B(G92gat), .Z(new_n631));
  INV_X1    g430(.A(G85gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G85gat), .A2(G92gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT7), .ZN(new_n635));
  INV_X1    g434(.A(G99gat), .ZN(new_n636));
  INV_X1    g435(.A(G106gat), .ZN(new_n637));
  OAI21_X1  g436(.A(KEYINPUT8), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n633), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(G99gat), .B(G106gat), .Z(new_n640));
  OR2_X1    g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n643), .B1(new_n550), .B2(new_n552), .ZN(new_n644));
  NAND2_X1  g443(.A1(G232gat), .A2(G233gat), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT41), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n643), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n647), .B1(new_n648), .B2(new_n541), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G190gat), .B(G218gat), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(KEYINPUT105), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n645), .A2(new_n646), .ZN(new_n654));
  INV_X1    g453(.A(G134gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(new_n223), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n650), .A2(new_n651), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n652), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n653), .A2(new_n659), .A3(new_n652), .A4(new_n657), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n577), .B1(new_n630), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n629), .A2(new_n663), .A3(KEYINPUT106), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n643), .A2(new_n603), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n641), .A2(new_n593), .A3(new_n602), .A4(new_n642), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT10), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT107), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n648), .A2(new_n604), .A3(KEYINPUT10), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT107), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n668), .A2(new_n669), .A3(new_n674), .A4(new_n670), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n672), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(G230gat), .A2(G233gat), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n668), .A2(new_n669), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(G230gat), .A3(G233gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(G120gat), .B(G148gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(G176gat), .B(G204gat), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n681), .B(new_n682), .Z(new_n683));
  NAND3_X1  g482(.A1(new_n678), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n677), .B(KEYINPUT108), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n676), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n683), .B1(new_n688), .B2(new_n680), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n667), .A2(new_n691), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n506), .A2(new_n576), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n435), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(G1gat), .ZN(G1324gat));
  INV_X1    g494(.A(KEYINPUT42), .ZN(new_n696));
  INV_X1    g495(.A(new_n499), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT16), .B(G8gat), .Z(new_n698));
  NAND3_X1  g497(.A1(new_n693), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n506), .A2(new_n697), .A3(new_n576), .A4(new_n692), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(G8gat), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n696), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT109), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n699), .A2(new_n696), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n705), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT109), .B1(new_n707), .B2(new_n702), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(G1325gat));
  INV_X1    g508(.A(new_n693), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n710), .A2(new_n514), .A3(new_n483), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n494), .A2(new_n496), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n514), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n713), .A2(KEYINPUT110), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(KEYINPUT110), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n711), .B1(new_n714), .B2(new_n715), .ZN(G1326gat));
  INV_X1    g515(.A(new_n292), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n693), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT43), .B(G22gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1327gat));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  INV_X1    g520(.A(new_n291), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n202), .B1(new_n289), .B2(new_n290), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n504), .B(new_n481), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT35), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n491), .A2(new_n498), .A3(new_n500), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n485), .A2(new_n483), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n725), .A2(new_n726), .B1(new_n727), .B2(new_n447), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n721), .B1(new_n728), .B2(new_n663), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n506), .A2(KEYINPUT44), .A3(new_n664), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT111), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n576), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n568), .A2(new_n575), .A3(KEYINPUT111), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n630), .A2(new_n690), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n731), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(G29gat), .B1(new_n738), .B2(new_n434), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n568), .A2(new_n575), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n728), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n736), .A2(new_n663), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n741), .A2(new_n533), .A3(new_n435), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT45), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n739), .A2(new_n744), .ZN(G1328gat));
  NAND2_X1  g544(.A1(new_n741), .A2(new_n742), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n746), .A2(G36gat), .A3(new_n499), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT46), .ZN(new_n748));
  OAI21_X1  g547(.A(G36gat), .B1(new_n738), .B2(new_n499), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(G1329gat));
  INV_X1    g549(.A(G43gat), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n483), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n731), .A2(new_n737), .A3(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n754), .A2(KEYINPUT47), .ZN(new_n755));
  INV_X1    g554(.A(new_n712), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n756), .A3(new_n742), .ZN(new_n757));
  AOI22_X1  g556(.A1(new_n757), .A2(new_n751), .B1(new_n754), .B2(KEYINPUT47), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n753), .A2(new_n755), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n755), .B1(new_n753), .B2(new_n758), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(G1330gat));
  NAND4_X1  g560(.A1(new_n731), .A2(G50gat), .A3(new_n717), .A4(new_n737), .ZN(new_n762));
  INV_X1    g561(.A(G50gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(new_n746), .B2(new_n292), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT48), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT48), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n762), .A2(new_n767), .A3(new_n764), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(G1331gat));
  INV_X1    g568(.A(new_n735), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n667), .A2(new_n770), .A3(new_n690), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n506), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n434), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(new_n587), .ZN(G1332gat));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n506), .A2(KEYINPUT113), .A3(new_n771), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n697), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n780));
  XOR2_X1   g579(.A(KEYINPUT49), .B(G64gat), .Z(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n779), .B2(new_n781), .ZN(G1333gat));
  NAND4_X1  g581(.A1(new_n776), .A2(G71gat), .A3(new_n482), .A4(new_n777), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n772), .A2(new_n712), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(G71gat), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g585(.A1(new_n778), .A2(new_n717), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g587(.A1(new_n735), .A2(new_n630), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n735), .A2(KEYINPUT114), .A3(new_n630), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT115), .B1(new_n793), .B2(new_n691), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n795));
  AOI211_X1 g594(.A(new_n795), .B(new_n690), .C1(new_n791), .C2(new_n792), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n729), .A2(new_n730), .A3(new_n435), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT116), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(G85gat), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n798), .A2(KEYINPUT116), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n506), .A2(new_n664), .A3(new_n793), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n725), .A2(new_n726), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n663), .B1(new_n805), .B2(new_n486), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n806), .A2(KEYINPUT51), .A3(new_n793), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n435), .A2(new_n632), .A3(new_n691), .ZN(new_n810));
  OAI22_X1  g609(.A1(new_n800), .A2(new_n801), .B1(new_n809), .B2(new_n810), .ZN(G1336gat));
  NAND4_X1  g610(.A1(new_n729), .A2(new_n730), .A3(new_n697), .A4(new_n797), .ZN(new_n812));
  INV_X1    g611(.A(new_n631), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n499), .A2(G92gat), .A3(new_n690), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT51), .B1(new_n806), .B2(new_n793), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n791), .A2(new_n792), .ZN(new_n817));
  NOR4_X1   g616(.A1(new_n728), .A2(new_n803), .A3(new_n663), .A4(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n815), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(KEYINPUT117), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n821), .A3(KEYINPUT52), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n814), .B(new_n819), .C1(KEYINPUT117), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(G1337gat));
  AND3_X1   g624(.A1(new_n731), .A2(new_n482), .A3(new_n797), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n756), .A2(new_n636), .A3(new_n691), .ZN(new_n827));
  OAI22_X1  g626(.A1(new_n826), .A2(new_n636), .B1(new_n809), .B2(new_n827), .ZN(G1338gat));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT118), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(KEYINPUT118), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n292), .A2(G106gat), .A3(new_n690), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n831), .B1(new_n808), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n729), .A2(new_n730), .A3(new_n717), .A4(new_n797), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(G106gat), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n830), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n832), .B1(new_n816), .B2(new_n818), .ZN(new_n837));
  INV_X1    g636(.A(new_n831), .ZN(new_n838));
  AND4_X1   g637(.A1(new_n830), .A2(new_n835), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n836), .A2(new_n839), .ZN(G1339gat));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n672), .A2(new_n686), .A3(new_n673), .A4(new_n675), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n678), .A2(KEYINPUT54), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n676), .A2(new_n844), .A3(new_n687), .ZN(new_n845));
  INV_X1    g644(.A(new_n683), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n841), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(new_n684), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n678), .A2(KEYINPUT54), .A3(new_n842), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n850), .A2(KEYINPUT55), .A3(new_n846), .A4(new_n845), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n849), .A2(new_n733), .A3(new_n734), .A4(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n574), .A2(new_n557), .A3(new_n566), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n544), .A2(new_n547), .A3(new_n509), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n554), .B1(new_n553), .B2(new_n545), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n565), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n853), .B(new_n856), .C1(new_n685), .C2(new_n689), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n664), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n848), .A2(new_n684), .A3(new_n851), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n853), .A2(new_n661), .A3(new_n662), .A4(new_n856), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n630), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n665), .A2(new_n666), .A3(new_n690), .A4(new_n735), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n717), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n697), .A2(new_n434), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n864), .A2(new_n756), .A3(new_n865), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n866), .A2(KEYINPUT119), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(KEYINPUT119), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n576), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(G113gat), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n434), .B1(new_n862), .B2(new_n863), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n503), .A2(new_n499), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n770), .A2(new_n294), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT120), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n870), .A2(new_n876), .ZN(G1340gat));
  AOI21_X1  g676(.A(G120gat), .B1(new_n873), .B2(new_n691), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n867), .A2(new_n868), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n690), .A2(new_n296), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(G1341gat));
  NAND3_X1  g680(.A1(new_n867), .A2(new_n629), .A3(new_n868), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(G127gat), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n873), .A2(new_n580), .A3(new_n629), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(G1342gat));
  NAND3_X1  g684(.A1(new_n867), .A2(new_n664), .A3(new_n868), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(G134gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n873), .A2(new_n655), .A3(new_n664), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT56), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n888), .A2(KEYINPUT56), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(G1343gat));
  NAND2_X1  g690(.A1(new_n865), .A2(new_n483), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n857), .B1(new_n859), .B2(new_n740), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n861), .B1(new_n894), .B2(new_n663), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n863), .B1(new_n895), .B2(new_n629), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n292), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n896), .A2(KEYINPUT121), .A3(new_n898), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n862), .A2(new_n863), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT57), .B1(new_n904), .B2(new_n717), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n893), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(G141gat), .B1(new_n906), .B2(new_n740), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT58), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n292), .A2(new_n482), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n904), .A2(new_n435), .A3(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n871), .A2(KEYINPUT122), .A3(new_n910), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n913), .A2(new_n499), .A3(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n740), .A2(G141gat), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n770), .B(new_n893), .C1(new_n903), .C2(new_n905), .ZN(new_n918));
  INV_X1    g717(.A(new_n911), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n916), .A2(new_n499), .ZN(new_n920));
  AOI22_X1  g719(.A1(new_n918), .A2(G141gat), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI22_X1  g720(.A1(new_n909), .A2(new_n917), .B1(new_n921), .B2(new_n908), .ZN(G1344gat));
  AND2_X1   g721(.A1(new_n691), .A2(new_n231), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n913), .A2(new_n499), .A3(new_n914), .A4(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n924), .B(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n231), .A2(KEYINPUT59), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n927), .B1(new_n906), .B2(new_n690), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT59), .ZN(new_n929));
  INV_X1    g728(.A(new_n898), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n930), .B1(new_n862), .B2(new_n863), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n665), .A2(new_n740), .A3(new_n666), .A4(new_n690), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n932), .B1(new_n895), .B2(new_n629), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT57), .B1(new_n933), .B2(new_n717), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n892), .A2(new_n690), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n229), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n928), .B1(new_n929), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n926), .A2(new_n938), .ZN(G1345gat));
  NAND3_X1  g738(.A1(new_n915), .A2(new_n222), .A3(new_n629), .ZN(new_n940));
  OAI21_X1  g739(.A(G155gat), .B1(new_n906), .B2(new_n630), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1346gat));
  NOR3_X1   g741(.A1(new_n906), .A2(new_n223), .A3(new_n663), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n915), .A2(new_n664), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n943), .B1(new_n944), .B2(new_n223), .ZN(G1347gat));
  AOI21_X1  g744(.A(new_n435), .B1(new_n862), .B2(new_n863), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n503), .A2(new_n697), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n947), .A2(KEYINPUT124), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(KEYINPUT124), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(G169gat), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n951), .A2(new_n952), .A3(new_n770), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT125), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n697), .A2(new_n434), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n955), .A2(new_n712), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n864), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(new_n576), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n954), .B1(new_n958), .B2(G169gat), .ZN(new_n959));
  AOI211_X1 g758(.A(KEYINPUT125), .B(new_n952), .C1(new_n957), .C2(new_n576), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n953), .B1(new_n959), .B2(new_n960), .ZN(G1348gat));
  INV_X1    g760(.A(G176gat), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n951), .A2(new_n962), .A3(new_n691), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n957), .A2(new_n691), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n963), .B1(new_n964), .B2(new_n962), .ZN(G1349gat));
  NAND2_X1  g764(.A1(new_n957), .A2(new_n629), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G183gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n951), .A2(new_n378), .A3(new_n629), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(KEYINPUT60), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT60), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n967), .A2(new_n971), .A3(new_n968), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(G1350gat));
  NAND3_X1  g772(.A1(new_n951), .A2(new_n358), .A3(new_n664), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT61), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n957), .A2(new_n664), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n975), .B1(new_n976), .B2(G190gat), .ZN(new_n977));
  AOI211_X1 g776(.A(KEYINPUT61), .B(new_n358), .C1(new_n957), .C2(new_n664), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n974), .B1(new_n977), .B2(new_n978), .ZN(G1351gat));
  AND3_X1   g778(.A1(new_n946), .A2(new_n697), .A3(new_n910), .ZN(new_n980));
  AOI21_X1  g779(.A(G197gat), .B1(new_n980), .B2(new_n770), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n483), .A2(new_n434), .A3(new_n697), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(KEYINPUT126), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n935), .A2(new_n983), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n576), .A2(G197gat), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n981), .B1(new_n984), .B2(new_n985), .ZN(G1352gat));
  NAND2_X1  g785(.A1(new_n984), .A2(new_n691), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(G204gat), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n690), .A2(G204gat), .ZN(new_n989));
  AND2_X1   g788(.A1(new_n980), .A2(new_n989), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n991));
  OR2_X1    g790(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n990), .A2(new_n991), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n988), .A2(new_n992), .A3(new_n993), .ZN(G1353gat));
  NAND4_X1  g793(.A1(new_n980), .A2(new_n237), .A3(new_n238), .A4(new_n629), .ZN(new_n995));
  OAI211_X1 g794(.A(new_n629), .B(new_n983), .C1(new_n931), .C2(new_n934), .ZN(new_n996));
  AND3_X1   g795(.A1(new_n996), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n997));
  AOI21_X1  g796(.A(KEYINPUT63), .B1(new_n996), .B2(G211gat), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT127), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g800(.A(new_n995), .B(KEYINPUT127), .C1(new_n997), .C2(new_n998), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1001), .A2(new_n1002), .ZN(G1354gat));
  AOI21_X1  g802(.A(G218gat), .B1(new_n980), .B2(new_n664), .ZN(new_n1004));
  AOI21_X1  g803(.A(new_n663), .B1(new_n241), .B2(new_n242), .ZN(new_n1005));
  AOI21_X1  g804(.A(new_n1004), .B1(new_n984), .B2(new_n1005), .ZN(G1355gat));
endmodule


