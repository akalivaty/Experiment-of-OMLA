//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  INV_X1    g0010(.A(G232), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n202), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n212), .B(new_n216), .C1(G107), .C2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G97), .A2(G257), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n217), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT65), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(new_n203), .ZN(new_n223));
  NAND2_X1  g0023(.A1(KEYINPUT65), .A2(G68), .ZN(new_n224));
  AND2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AND2_X1   g0025(.A1(new_n225), .A2(G238), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n207), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(KEYINPUT64), .ZN(new_n230));
  INV_X1    g0030(.A(KEYINPUT64), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G20), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n202), .A2(new_n203), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n236), .A2(G50), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(new_n238));
  AOI211_X1 g0038(.A(new_n210), .B(new_n228), .C1(new_n235), .C2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n211), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT2), .B(G226), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G257), .ZN(new_n245));
  XOR2_X1   g0045(.A(KEYINPUT66), .B(G250), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n243), .B(new_n247), .Z(G358));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G68), .B(G77), .Z(new_n252));
  XNOR2_X1  g0052(.A(G50), .B(G58), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n229), .A2(new_n256), .A3(KEYINPUT68), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT68), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(G20), .B2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n260), .A2(G150), .B1(G20), .B2(new_n204), .ZN(new_n261));
  AOI21_X1  g0061(.A(KEYINPUT67), .B1(new_n202), .B2(KEYINPUT8), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT8), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G58), .ZN(new_n264));
  MUX2_X1   g0064(.A(KEYINPUT67), .B(new_n262), .S(new_n264), .Z(new_n265));
  AOI21_X1  g0065(.A(new_n256), .B1(new_n230), .B2(new_n232), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n261), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n234), .ZN(new_n270));
  INV_X1    g0070(.A(G1), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G13), .A3(G20), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n268), .A2(new_n270), .B1(new_n201), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n270), .B1(new_n271), .B2(G20), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G50), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT9), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT72), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n277), .B(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT3), .B(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G222), .A2(G1698), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G223), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n234), .B1(G33), .B2(G41), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n285), .B(new_n286), .C1(G77), .C2(new_n281), .ZN(new_n287));
  INV_X1    g0087(.A(new_n234), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G41), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n271), .B1(G41), .B2(G45), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G226), .ZN(new_n294));
  INV_X1    g0094(.A(G274), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n287), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G190), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n298), .A2(new_n299), .B1(KEYINPUT72), .B2(new_n278), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n280), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n298), .A2(G200), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n302), .B(new_n303), .C1(KEYINPUT73), .C2(KEYINPUT10), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n280), .A2(new_n303), .A3(new_n301), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n280), .A2(KEYINPUT73), .A3(new_n301), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT10), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n298), .A2(new_n309), .ZN(new_n310));
  XOR2_X1   g0110(.A(KEYINPUT69), .B(G179), .Z(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n277), .B(new_n310), .C1(new_n312), .C2(new_n298), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n281), .A2(G238), .A3(G1698), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n281), .A2(G232), .A3(new_n283), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT3), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G33), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G107), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n314), .A2(new_n315), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n296), .B1(new_n321), .B2(new_n286), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n293), .A2(G244), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n311), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n264), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n260), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT70), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT64), .B(G20), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G77), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n259), .A2(new_n257), .B1(new_n264), .B2(new_n327), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n230), .A2(new_n232), .A3(G77), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT70), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  XOR2_X1   g0136(.A(KEYINPUT15), .B(G87), .Z(new_n337));
  NAND2_X1  g0137(.A1(new_n266), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n333), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n270), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n273), .A2(new_n219), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n275), .A2(G77), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n324), .A2(new_n309), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n326), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n304), .A2(new_n308), .A3(new_n313), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n265), .A2(new_n272), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n275), .B2(new_n265), .ZN(new_n348));
  INV_X1    g0148(.A(G159), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(new_n257), .B2(new_n259), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n223), .A2(G58), .A3(new_n224), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n236), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n350), .B1(new_n352), .B2(G20), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n231), .A2(G20), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n229), .A2(KEYINPUT64), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT77), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n319), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n281), .A2(KEYINPUT77), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(G20), .B1(new_n316), .B2(new_n318), .ZN(new_n362));
  OAI21_X1  g0162(.A(G68), .B1(new_n362), .B2(new_n354), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n353), .B(KEYINPUT16), .C1(new_n361), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n270), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT7), .B1(new_n331), .B2(new_n281), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n319), .A2(new_n354), .A3(new_n229), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n225), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT16), .B1(new_n368), .B2(new_n353), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n348), .B1(new_n365), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n316), .A2(new_n318), .A3(G223), .A4(new_n283), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT78), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n281), .A2(KEYINPUT78), .A3(G223), .A4(new_n283), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n281), .A2(G226), .A3(G1698), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G33), .A2(G87), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n377), .B(KEYINPUT79), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n374), .A2(new_n375), .A3(new_n376), .A4(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n286), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n292), .A2(new_n211), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n380), .A2(G190), .A3(new_n297), .A4(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n380), .A2(new_n297), .A3(new_n382), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G200), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n371), .A2(KEYINPUT17), .A3(new_n383), .A4(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n368), .A2(new_n353), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT16), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n389), .A2(new_n270), .A3(new_n364), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n385), .A2(new_n390), .A3(new_n383), .A4(new_n348), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT17), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n380), .A2(new_n297), .A3(new_n382), .A4(new_n312), .ZN(new_n394));
  AOI211_X1 g0194(.A(new_n296), .B(new_n381), .C1(new_n379), .C2(new_n286), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n394), .B1(new_n395), .B2(new_n309), .ZN(new_n396));
  AND3_X1   g0196(.A1(new_n396), .A2(new_n370), .A3(KEYINPUT18), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT18), .B1(new_n396), .B2(new_n370), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n386), .B(new_n393), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT13), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n281), .A2(G226), .A3(new_n283), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G97), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n316), .A2(new_n318), .A3(G232), .A4(G1698), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n286), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n293), .A2(G238), .ZN(new_n407));
  AND4_X1   g0207(.A1(new_n401), .A2(new_n406), .A3(new_n407), .A4(new_n297), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n296), .B1(new_n405), .B2(new_n286), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n401), .B1(new_n409), .B2(new_n407), .ZN(new_n410));
  OAI21_X1  g0210(.A(G169), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT14), .ZN(new_n412));
  INV_X1    g0212(.A(new_n408), .ZN(new_n413));
  INV_X1    g0213(.A(new_n410), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(G179), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT14), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n416), .B(G169), .C1(new_n408), .C2(new_n410), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n412), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n260), .A2(G50), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n419), .B1(new_n225), .B2(new_n229), .C1(new_n267), .C2(new_n219), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n270), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT11), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n421), .A2(KEYINPUT11), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT12), .B1(new_n225), .B2(new_n272), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT75), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT75), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n426), .B(KEYINPUT12), .C1(new_n225), .C2(new_n272), .ZN(new_n427));
  OR3_X1    g0227(.A1(new_n272), .A2(KEYINPUT12), .A3(G68), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n425), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n275), .A2(G68), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT76), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT76), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n429), .A2(new_n433), .A3(new_n430), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n422), .A2(new_n423), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n418), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(G200), .B1(new_n408), .B2(new_n410), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT74), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n413), .A2(G190), .A3(new_n414), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT74), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(G200), .C1(new_n408), .C2(new_n410), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n435), .A2(new_n439), .A3(new_n440), .A4(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n400), .A2(new_n437), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G200), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n445), .B1(new_n322), .B2(new_n323), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT71), .B1(new_n343), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n324), .A2(G200), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n339), .A2(new_n270), .B1(new_n219), .B2(new_n273), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT71), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n448), .A2(new_n449), .A3(new_n450), .A4(new_n342), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n325), .A2(G190), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n447), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n346), .A2(new_n444), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n233), .A2(new_n281), .A3(G87), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT22), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT22), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n233), .A2(new_n281), .A3(new_n459), .A4(G87), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(KEYINPUT23), .A2(G107), .ZN(new_n462));
  OR2_X1    g0262(.A1(KEYINPUT80), .A2(G116), .ZN(new_n463));
  NAND2_X1  g0263(.A1(KEYINPUT80), .A2(G116), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(G33), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT23), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(KEYINPUT23), .A2(G107), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n467), .A2(new_n229), .B1(new_n331), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n461), .A2(new_n462), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT24), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT24), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n461), .A2(new_n469), .A3(new_n472), .A4(new_n462), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n270), .ZN(new_n475));
  INV_X1    g0275(.A(new_n270), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n476), .B(new_n272), .C1(G1), .C2(new_n256), .ZN(new_n477));
  INV_X1    g0277(.A(G107), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n272), .A2(G107), .ZN(new_n481));
  XNOR2_X1  g0281(.A(new_n481), .B(KEYINPUT25), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n475), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n316), .A2(new_n318), .A3(G257), .A4(G1698), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT84), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n281), .A2(KEYINPUT84), .A3(G257), .A4(G1698), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G294), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n281), .A2(G250), .A3(new_n283), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n486), .A2(new_n487), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n286), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n271), .A2(G45), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(new_n295), .ZN(new_n493));
  XNOR2_X1  g0293(.A(KEYINPUT5), .B(G41), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(G45), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(G1), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n286), .B1(new_n497), .B2(new_n494), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G264), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n491), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n500), .A2(G169), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G179), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n483), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(G97), .A2(G107), .ZN(new_n506));
  AND2_X1   g0306(.A1(KEYINPUT81), .A2(G87), .ZN(new_n507));
  NOR2_X1   g0307(.A1(KEYINPUT81), .A2(G87), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AND3_X1   g0309(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n509), .B1(new_n331), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n233), .A2(new_n281), .A3(G68), .ZN(new_n512));
  INV_X1    g0312(.A(G97), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n331), .A2(new_n256), .A3(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n511), .B(new_n512), .C1(new_n514), .C2(KEYINPUT19), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n270), .ZN(new_n516));
  INV_X1    g0316(.A(new_n477), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n337), .ZN(new_n518));
  INV_X1    g0318(.A(new_n337), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n273), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n516), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  OR2_X1    g0321(.A1(G238), .A2(G1698), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n220), .A2(G1698), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n316), .A2(new_n522), .A3(new_n318), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n465), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n286), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n497), .B1(new_n288), .B2(new_n289), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n493), .B1(new_n527), .B2(G250), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n311), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n309), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n521), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n515), .A2(new_n270), .B1(new_n273), .B2(new_n519), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n529), .A2(G200), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n526), .A2(G190), .A3(new_n528), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n517), .A2(G87), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n534), .A2(new_n535), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n533), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n505), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n491), .A2(new_n299), .A3(new_n495), .A4(new_n499), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(new_n500), .B2(G200), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n475), .A2(new_n543), .A3(new_n480), .A4(new_n482), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n517), .A2(G116), .ZN(new_n545));
  AND2_X1   g0345(.A1(KEYINPUT80), .A2(G116), .ZN(new_n546));
  NOR2_X1   g0346(.A1(KEYINPUT80), .A2(G116), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n273), .ZN(new_n550));
  XNOR2_X1  g0350(.A(new_n550), .B(KEYINPUT82), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G283), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n256), .A2(G97), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n552), .B(new_n553), .C1(new_n355), .C2(new_n356), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT83), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT83), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n233), .A2(new_n556), .A3(new_n552), .A4(new_n553), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n270), .B1(new_n548), .B2(new_n229), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT20), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT20), .ZN(new_n562));
  AOI211_X1 g0362(.A(new_n562), .B(new_n559), .C1(new_n555), .C2(new_n557), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n545), .B(new_n551), .C1(new_n561), .C2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n281), .A2(G264), .A3(G1698), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n319), .A2(G303), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n316), .A2(new_n318), .A3(G257), .A4(new_n283), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n286), .ZN(new_n569));
  INV_X1    g0369(.A(G41), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT5), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT5), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(G41), .ZN(new_n573));
  AND4_X1   g0373(.A1(G274), .A2(new_n497), .A3(new_n571), .A4(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n498), .B2(G270), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n576), .A2(new_n309), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n564), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT21), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n569), .A2(new_n575), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(KEYINPUT21), .A3(G169), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n569), .A2(new_n575), .A3(G179), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n578), .A2(new_n579), .B1(new_n564), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n316), .A2(new_n318), .A3(G244), .A4(new_n283), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT4), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n281), .A2(KEYINPUT4), .A3(G244), .A4(new_n283), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n281), .A2(G250), .A3(G1698), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n552), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n286), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n571), .A2(new_n573), .ZN(new_n593));
  OAI211_X1 g0393(.A(G257), .B(new_n290), .C1(new_n593), .C2(new_n492), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n495), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n309), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n272), .A2(G97), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT6), .ZN(new_n600));
  AND2_X1   g0400(.A1(G97), .A2(G107), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n600), .B1(new_n601), .B2(new_n506), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n478), .A2(KEYINPUT6), .A3(G97), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n604), .A2(new_n331), .B1(G77), .B2(new_n260), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n366), .A2(G107), .A3(new_n367), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n599), .B1(new_n607), .B2(new_n270), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n477), .A2(new_n513), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n587), .A2(new_n588), .A3(new_n552), .A4(new_n590), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n595), .B1(new_n611), .B2(new_n286), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n608), .A2(new_n610), .B1(new_n311), .B2(new_n612), .ZN(new_n613));
  AOI211_X1 g0413(.A(new_n299), .B(new_n595), .C1(new_n286), .C2(new_n611), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n445), .B1(new_n592), .B2(new_n596), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI211_X1 g0416(.A(new_n599), .B(new_n609), .C1(new_n607), .C2(new_n270), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n598), .A2(new_n613), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n564), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n576), .A2(G190), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n619), .B(new_n620), .C1(new_n445), .C2(new_n576), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n544), .A2(new_n584), .A3(new_n618), .A4(new_n621), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n456), .A2(new_n541), .A3(new_n622), .ZN(G372));
  NAND2_X1  g0423(.A1(new_n386), .A2(new_n393), .ZN(new_n624));
  INV_X1    g0424(.A(new_n345), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n443), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n624), .B1(new_n626), .B2(new_n437), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n397), .A2(new_n398), .ZN(new_n628));
  OR3_X1    g0428(.A1(new_n627), .A2(KEYINPUT88), .A3(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n304), .A2(new_n308), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT88), .B1(new_n627), .B2(new_n628), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n632), .A2(new_n313), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n534), .A2(new_n518), .B1(new_n530), .B2(new_n311), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT85), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n635), .B1(new_n525), .B2(new_n286), .ZN(new_n636));
  AOI211_X1 g0436(.A(KEYINPUT85), .B(new_n290), .C1(new_n524), .C2(new_n465), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n528), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n309), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  AND4_X1   g0440(.A1(new_n516), .A2(new_n536), .A3(new_n520), .A4(new_n537), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n638), .A2(G200), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n634), .A2(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n607), .A2(new_n270), .ZN(new_n644));
  INV_X1    g0444(.A(new_n599), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(new_n645), .A3(new_n610), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n612), .A2(new_n311), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n646), .A2(new_n598), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(KEYINPUT26), .B1(new_n643), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n646), .A2(new_n598), .A3(new_n647), .ZN(new_n650));
  XNOR2_X1  g0450(.A(KEYINPUT86), .B(KEYINPUT26), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n539), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n640), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT87), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n505), .A2(new_n584), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n544), .A2(new_n618), .A3(new_n643), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OAI211_X1 g0458(.A(KEYINPUT87), .B(new_n640), .C1(new_n649), .C2(new_n652), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n655), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n455), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n633), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT89), .ZN(G369));
  INV_X1    g0463(.A(G13), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n331), .A2(G1), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT91), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(new_n667), .A3(KEYINPUT27), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT27), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT91), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G213), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n665), .A2(KEYINPUT90), .A3(new_n669), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n233), .A2(new_n669), .A3(new_n271), .A4(G13), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT90), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n672), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n679), .A2(G343), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n564), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n584), .A2(new_n681), .A3(new_n621), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n584), .B2(new_n681), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT92), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT92), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n683), .A2(new_n686), .A3(G330), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n483), .A2(new_n680), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n544), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n505), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n479), .B1(new_n474), .B2(new_n270), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n501), .B1(new_n693), .B2(new_n482), .ZN(new_n694));
  INV_X1    g0494(.A(new_n680), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(new_n504), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n688), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n584), .A2(new_n680), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n697), .B1(new_n691), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(G399));
  NOR2_X1   g0502(.A1(new_n507), .A2(new_n508), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(G116), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(new_n705), .A3(new_n506), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT93), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n208), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n708), .A2(G1), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n237), .B2(new_n711), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n651), .B1(new_n539), .B2(new_n650), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT96), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n643), .A2(new_n648), .A3(KEYINPUT26), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT96), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n718), .B(new_n651), .C1(new_n539), .C2(new_n650), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n716), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n658), .A2(new_n640), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(KEYINPUT29), .A3(new_n695), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n660), .A2(new_n695), .ZN(new_n723));
  XNOR2_X1  g0523(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n582), .A2(new_n529), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n491), .A2(new_n499), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n726), .A2(new_n727), .A3(new_n612), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n500), .A2(new_n612), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(new_n311), .A3(new_n580), .A4(new_n638), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n728), .A2(KEYINPUT94), .A3(new_n729), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n730), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(KEYINPUT94), .B1(new_n728), .B2(new_n729), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n695), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n539), .B1(new_n694), .B2(new_n504), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n544), .A2(new_n618), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n584), .A2(new_n621), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n738), .A2(new_n739), .A3(new_n740), .A4(new_n695), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n737), .B1(new_n741), .B2(KEYINPUT31), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n730), .A2(new_n732), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n743), .B1(new_n729), .B2(new_n728), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n744), .A2(new_n745), .A3(new_n695), .ZN(new_n746));
  OAI21_X1  g0546(.A(G330), .B1(new_n742), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n725), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n714), .B1(new_n749), .B2(G1), .ZN(G364));
  NAND3_X1  g0550(.A1(new_n312), .A2(G190), .A3(new_n331), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n445), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n233), .A2(G190), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n312), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G200), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n752), .A2(G50), .B1(new_n755), .B2(G77), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n751), .A2(G200), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n756), .B1(new_n202), .B2(new_n758), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT97), .Z(new_n760));
  NAND2_X1  g0560(.A1(new_n753), .A2(new_n503), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n445), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n478), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n754), .A2(new_n445), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n503), .A2(G190), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n767), .A2(new_n229), .A3(new_n445), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n766), .A2(new_n203), .B1(new_n704), .B2(new_n769), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n760), .A2(new_n764), .A3(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT32), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n761), .A2(G200), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n772), .B1(new_n774), .B2(new_n349), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n773), .A2(KEYINPUT32), .A3(G159), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n319), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n331), .B1(G200), .B2(new_n767), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n771), .B(new_n777), .C1(new_n513), .C2(new_n779), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n755), .A2(G311), .ZN(new_n781));
  INV_X1    g0581(.A(G322), .ZN(new_n782));
  XOR2_X1   g0582(.A(KEYINPUT33), .B(G317), .Z(new_n783));
  OAI22_X1  g0583(.A1(new_n758), .A2(new_n782), .B1(new_n766), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT98), .ZN(new_n785));
  INV_X1    g0585(.A(new_n752), .ZN(new_n786));
  INV_X1    g0586(.A(G326), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G283), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n319), .B1(new_n763), .B2(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n788), .B(new_n790), .C1(G329), .C2(new_n773), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n778), .A2(G294), .B1(new_n768), .B2(G303), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n785), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n780), .B1(new_n781), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n234), .B1(G20), .B2(new_n309), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n331), .A2(new_n664), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n271), .B1(new_n797), .B2(G45), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n710), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G13), .A2(G33), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n683), .A2(new_n804), .ZN(new_n805));
  AND3_X1   g0605(.A1(new_n316), .A2(new_n318), .A3(KEYINPUT77), .ZN(new_n806));
  AOI21_X1  g0606(.A(KEYINPUT77), .B1(new_n316), .B2(new_n318), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n709), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n238), .A2(new_n496), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n809), .B(new_n810), .C1(new_n254), .C2(new_n496), .ZN(new_n811));
  INV_X1    g0611(.A(G355), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n281), .A2(new_n208), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n811), .B1(G116), .B2(new_n208), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n803), .A2(new_n795), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n796), .A2(new_n800), .A3(new_n805), .A4(new_n816), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT99), .Z(new_n818));
  NOR2_X1   g0618(.A1(new_n683), .A2(G330), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n688), .A2(new_n800), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G396));
  NAND2_X1  g0622(.A1(new_n680), .A2(new_n343), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n453), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n345), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT102), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n345), .A2(new_n680), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n625), .B1(new_n453), .B2(new_n823), .ZN(new_n830));
  OAI21_X1  g0630(.A(KEYINPUT102), .B1(new_n830), .B2(new_n827), .ZN(new_n831));
  AND3_X1   g0631(.A1(new_n829), .A2(KEYINPUT103), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(KEYINPUT103), .B1(new_n829), .B2(new_n831), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n829), .A2(new_n831), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  MUX2_X1   g0637(.A(new_n835), .B(new_n837), .S(new_n723), .Z(new_n838));
  INV_X1    g0638(.A(new_n747), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n800), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n838), .A2(new_n839), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n808), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n757), .A2(G143), .B1(new_n765), .B2(G150), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n752), .A2(G137), .ZN(new_n846));
  INV_X1    g0646(.A(new_n755), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n845), .B(new_n846), .C1(new_n349), .C2(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(KEYINPUT101), .B(KEYINPUT34), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n848), .B(new_n849), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n778), .A2(G58), .B1(new_n768), .B2(G50), .ZN(new_n851));
  INV_X1    g0651(.A(G132), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n850), .B(new_n851), .C1(new_n852), .C2(new_n774), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n844), .B(new_n853), .C1(G68), .C2(new_n762), .ZN(new_n854));
  AOI22_X1  g0654(.A1(G294), .A2(new_n757), .B1(new_n752), .B2(G303), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n549), .B2(new_n847), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G87), .A2(new_n762), .B1(new_n773), .B2(G311), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n281), .B1(new_n778), .B2(G97), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n857), .B(new_n858), .C1(new_n478), .C2(new_n769), .ZN(new_n859));
  XNOR2_X1  g0659(.A(KEYINPUT100), .B(G283), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n856), .B(new_n859), .C1(new_n765), .C2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n795), .B1(new_n854), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n841), .B1(new_n837), .B2(new_n801), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n795), .A2(new_n801), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n862), .B(new_n863), .C1(G77), .C2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n843), .A2(new_n866), .ZN(G384));
  NOR2_X1   g0667(.A1(new_n797), .A2(new_n271), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n436), .A2(new_n680), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n437), .A2(new_n443), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n418), .A2(new_n436), .A3(new_n680), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n826), .B1(new_n825), .B2(new_n828), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n830), .A2(KEYINPUT102), .A3(new_n827), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n730), .A2(new_n732), .A3(new_n733), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n680), .B1(new_n876), .B2(new_n735), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n541), .A2(new_n622), .A3(new_n680), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n877), .B1(new_n878), .B2(new_n745), .ZN(new_n879));
  OAI211_X1 g0679(.A(KEYINPUT31), .B(new_n680), .C1(new_n876), .C2(new_n735), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n875), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT105), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n319), .A2(new_n229), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n203), .B1(new_n883), .B2(KEYINPUT7), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n357), .B2(new_n808), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT16), .B1(new_n885), .B2(new_n353), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n348), .B1(new_n365), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n396), .B2(new_n679), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n391), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT37), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n396), .A2(new_n370), .ZN(new_n891));
  AOI211_X1 g0691(.A(KEYINPUT104), .B(new_n678), .C1(new_n390), .C2(new_n348), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT104), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n370), .B2(new_n679), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n391), .B(new_n891), .C1(new_n892), .C2(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n882), .B(new_n890), .C1(new_n895), .C2(KEYINPUT37), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n370), .A2(new_n679), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT104), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n370), .A2(new_n893), .A3(new_n679), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT37), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n891), .A2(new_n391), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n882), .B1(new_n904), .B2(new_n890), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n897), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n399), .A2(new_n679), .A3(new_n887), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT38), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n890), .B1(new_n895), .B2(KEYINPUT37), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT105), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n910), .A2(KEYINPUT38), .A3(new_n907), .A4(new_n896), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n881), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  XOR2_X1   g0713(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT40), .ZN(new_n916));
  INV_X1    g0716(.A(new_n901), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n399), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n895), .A2(KEYINPUT37), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n902), .B1(new_n901), .B2(new_n903), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT38), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n916), .B1(new_n911), .B2(new_n923), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n913), .A2(new_n915), .B1(new_n881), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n880), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n925), .B1(new_n742), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n927), .A2(new_n456), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n924), .A2(new_n881), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n829), .A2(new_n831), .B1(new_n870), .B2(new_n871), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n742), .B2(new_n926), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n910), .A2(new_n907), .A3(new_n896), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n922), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n931), .B1(new_n911), .B2(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(G330), .B(new_n929), .C1(new_n934), .C2(new_n914), .ZN(new_n935));
  INV_X1    g0735(.A(G330), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n879), .B2(new_n880), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n455), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n928), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  NOR3_X1   g0739(.A1(new_n397), .A2(new_n398), .A3(new_n679), .ZN(new_n940));
  INV_X1    g0740(.A(new_n872), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n660), .A2(new_n695), .A3(new_n836), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n941), .B1(new_n942), .B2(new_n828), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n933), .A2(new_n911), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n933), .A2(KEYINPUT39), .A3(new_n911), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n911), .A2(new_n923), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT39), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n437), .A2(new_n680), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n946), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n945), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n455), .B(new_n722), .C1(new_n723), .C2(new_n724), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n633), .A2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n952), .B(new_n954), .Z(new_n955));
  AOI21_X1  g0755(.A(new_n868), .B1(new_n939), .B2(new_n955), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT107), .Z(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n955), .B2(new_n939), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n705), .B1(new_n604), .B2(KEYINPUT35), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n959), .B(new_n235), .C1(KEYINPUT35), .C2(new_n604), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT36), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n238), .A2(G77), .A3(new_n351), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(G50), .B2(new_n203), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n963), .A2(G1), .A3(new_n664), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n958), .A2(new_n961), .A3(new_n964), .ZN(G367));
  INV_X1    g0765(.A(new_n699), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n680), .A2(new_n646), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n618), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n648), .B2(new_n680), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n966), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT108), .Z(new_n973));
  INV_X1    g0773(.A(new_n701), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n696), .A2(KEYINPUT42), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n974), .A2(new_n969), .A3(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n691), .A2(new_n696), .A3(new_n700), .ZN(new_n977));
  OAI21_X1  g0777(.A(KEYINPUT42), .B1(new_n977), .B2(new_n968), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n976), .B(new_n978), .C1(new_n650), .C2(new_n680), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT43), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n534), .A2(new_n537), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n680), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n983), .A2(new_n640), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(new_n643), .B2(new_n983), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n979), .B2(new_n980), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n981), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n981), .A2(new_n986), .ZN(new_n988));
  OR3_X1    g0788(.A1(new_n973), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n987), .A2(new_n988), .B1(KEYINPUT108), .B2(new_n972), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n710), .B(KEYINPUT41), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n692), .A2(new_n697), .B1(new_n584), .B2(new_n680), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT110), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n995), .A2(new_n687), .A3(new_n685), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n688), .A2(new_n994), .A3(new_n993), .ZN(new_n997));
  INV_X1    g0797(.A(new_n977), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n998), .B1(new_n996), .B2(new_n997), .ZN(new_n1001));
  NOR3_X1   g0801(.A1(new_n1000), .A2(new_n1001), .A3(new_n748), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n701), .A2(new_n971), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT45), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n701), .A2(new_n971), .A3(KEYINPUT45), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n974), .A2(new_n970), .ZN(new_n1008));
  XOR2_X1   g0808(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n974), .A2(new_n970), .A3(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1007), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT111), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1013), .A2(new_n1014), .A3(new_n699), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n966), .A2(KEYINPUT111), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1005), .A2(new_n1006), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n699), .A2(new_n1014), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .A4(new_n1012), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1002), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n992), .B1(new_n1021), .B2(new_n749), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n989), .B(new_n990), .C1(new_n1022), .C2(new_n799), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n757), .A2(G150), .B1(new_n762), .B2(G77), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n201), .B2(new_n847), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G58), .B2(new_n768), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n773), .A2(G137), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n778), .A2(G68), .ZN(new_n1028));
  INV_X1    g0828(.A(G143), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n281), .B1(new_n786), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G159), .B2(new_n765), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n762), .A2(G97), .ZN(new_n1033));
  INV_X1    g0833(.A(G303), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1033), .B1(new_n478), .B2(new_n779), .C1(new_n758), .C2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(G317), .B2(new_n773), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n752), .A2(G311), .B1(new_n765), .B2(G294), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT46), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n769), .B2(new_n549), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1038), .A2(new_n705), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n808), .B1(new_n768), .B2(new_n1040), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1036), .A2(new_n1037), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n860), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n847), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1032), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT47), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n795), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n985), .A2(new_n803), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n815), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n247), .B2(new_n809), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n208), .B2(new_n519), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1047), .A2(new_n800), .A3(new_n1048), .A4(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1023), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT112), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1023), .A2(KEYINPUT112), .A3(new_n1052), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(G387));
  OAI21_X1  g0857(.A(KEYINPUT114), .B1(new_n1002), .B2(new_n711), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n996), .A2(new_n997), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n977), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n749), .A2(new_n1060), .A3(new_n999), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT114), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1061), .A2(new_n1062), .A3(new_n710), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1058), .A2(new_n749), .A3(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G50), .A2(new_n757), .B1(new_n752), .B2(G159), .ZN(new_n1065));
  INV_X1    g0865(.A(G150), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1065), .B(new_n808), .C1(new_n1066), .C2(new_n774), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n265), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1067), .B1(new_n1068), .B2(new_n765), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n755), .A2(G68), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n778), .A2(new_n337), .B1(new_n768), .B2(G77), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1069), .A2(new_n1033), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n757), .A2(G317), .B1(new_n765), .B2(G311), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n1034), .B2(new_n847), .C1(new_n782), .C2(new_n786), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT48), .ZN(new_n1075));
  INV_X1    g0875(.A(G294), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1075), .B1(new_n1076), .B2(new_n769), .C1(new_n779), .C2(new_n1043), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT49), .Z(new_n1078));
  OAI221_X1 g0878(.A(new_n844), .B1(new_n774), .B2(new_n787), .C1(new_n549), .C2(new_n763), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1072), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n795), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n809), .B1(new_n243), .B2(new_n496), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n708), .B2(new_n813), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n707), .B1(G68), .B2(G77), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n328), .A2(new_n201), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT50), .Z(new_n1086));
  NAND3_X1  g0886(.A1(new_n1084), .A2(new_n496), .A3(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1083), .A2(new_n1087), .B1(new_n478), .B2(new_n709), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n800), .B1(new_n1088), .B2(new_n1049), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT113), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1081), .B(new_n1090), .C1(new_n698), .C2(new_n804), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n799), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1060), .A2(new_n999), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1064), .B(new_n1091), .C1(new_n1092), .C2(new_n1093), .ZN(G393));
  NAND3_X1  g0894(.A1(new_n1061), .A2(new_n1015), .A3(new_n1019), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1021), .A2(new_n1095), .A3(new_n710), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(KEYINPUT115), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT115), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1021), .A2(new_n1095), .A3(new_n1098), .A4(new_n710), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1020), .A2(new_n799), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n841), .B1(new_n970), .B2(new_n803), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n809), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n815), .B1(new_n513), .B2(new_n208), .C1(new_n1103), .C2(new_n251), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n795), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n762), .A2(G87), .B1(G77), .B2(new_n778), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n1029), .B2(new_n774), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n844), .B(new_n1107), .C1(new_n328), .C2(new_n755), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n225), .A2(new_n768), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(G150), .A2(new_n752), .B1(new_n757), .B2(G159), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1110), .A2(KEYINPUT51), .B1(G50), .B2(new_n765), .ZN(new_n1111));
  OR2_X1    g0911(.A1(new_n1110), .A2(KEYINPUT51), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1108), .A2(new_n1109), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G311), .A2(new_n757), .B1(new_n752), .B2(G317), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT52), .Z(new_n1115));
  OAI22_X1  g0915(.A1(new_n766), .A2(new_n1034), .B1(new_n769), .B2(new_n1043), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1116), .A2(new_n764), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n774), .A2(new_n782), .B1(new_n549), .B2(new_n779), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(G294), .B2(new_n755), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1115), .A2(new_n319), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1113), .A2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1102), .B(new_n1104), .C1(new_n1105), .C2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1100), .A2(new_n1101), .A3(new_n1122), .ZN(G390));
  NAND2_X1  g0923(.A1(new_n937), .A2(new_n930), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n942), .A2(new_n828), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n872), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n950), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1127), .A2(new_n1128), .B1(new_n946), .B2(new_n949), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n947), .A2(new_n1128), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n721), .A2(new_n695), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n828), .B1(new_n1131), .B2(new_n837), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1130), .B1(new_n872), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1125), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n872), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1135), .A2(new_n1128), .A3(new_n947), .ZN(new_n1136));
  OAI211_X1 g0936(.A(G330), .B(new_n930), .C1(new_n742), .C2(new_n746), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n946), .A2(new_n949), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n943), .A2(new_n950), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1136), .B(new_n1137), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1134), .A2(new_n1140), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n633), .A2(new_n953), .A3(new_n938), .ZN(new_n1142));
  OAI21_X1  g0942(.A(G330), .B1(new_n742), .B2(new_n926), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n941), .B1(new_n1143), .B2(new_n834), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1132), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1144), .A2(new_n1145), .A3(new_n1137), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  OAI211_X1 g0947(.A(G330), .B(new_n836), .C1(new_n742), .C2(new_n746), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n941), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1124), .A2(new_n1149), .B1(new_n828), .B2(new_n942), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1142), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1141), .A2(KEYINPUT116), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n633), .A2(new_n953), .A3(new_n938), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1124), .A2(new_n1149), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n1126), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1153), .B1(new_n1155), .B2(new_n1146), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT116), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1140), .B(new_n1134), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1152), .A2(new_n1158), .A3(new_n710), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n946), .A2(new_n949), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n841), .B1(new_n1160), .B2(new_n801), .ZN(new_n1161));
  INV_X1    g0961(.A(G125), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n281), .B1(new_n774), .B2(new_n1162), .C1(new_n201), .C2(new_n763), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT117), .Z(new_n1164));
  XOR2_X1   g0964(.A(KEYINPUT54), .B(G143), .Z(new_n1165));
  AOI22_X1  g0965(.A1(G137), .A2(new_n765), .B1(new_n755), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(G128), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1166), .B1(new_n1167), .B2(new_n786), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1164), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n768), .A2(G150), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n1170), .B(KEYINPUT53), .Z(new_n1171));
  OAI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(new_n349), .C2(new_n779), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G132), .B2(new_n757), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n705), .A2(new_n758), .B1(new_n786), .B2(new_n789), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G294), .B2(new_n773), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n478), .B2(new_n766), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n847), .A2(new_n513), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n319), .B1(new_n779), .B2(new_n219), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n763), .A2(new_n203), .B1(new_n214), .B2(new_n769), .ZN(new_n1179));
  NOR4_X1   g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n795), .B1(new_n1173), .B2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1161), .B(new_n1181), .C1(new_n1068), .C2(new_n865), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT118), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1182), .B(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1134), .A2(new_n799), .A3(new_n1140), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1159), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(G378));
  NAND2_X1  g0987(.A1(new_n1155), .A2(new_n1146), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1134), .A2(new_n1188), .A3(new_n1140), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1142), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n935), .A2(new_n951), .A3(new_n945), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n952), .A2(new_n925), .A3(G330), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  XOR2_X1   g0993(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n304), .A2(new_n308), .A3(new_n313), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT55), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1196), .B(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n678), .B1(new_n276), .B2(new_n274), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1195), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1203), .A2(new_n1194), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1202), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1193), .A2(new_n1206), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1202), .A2(new_n1205), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1208), .A2(new_n1192), .A3(new_n1191), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1190), .A2(new_n1207), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT57), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1190), .A2(new_n1207), .A3(KEYINPUT57), .A4(new_n1209), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(new_n710), .A3(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1207), .A2(new_n799), .A3(new_n1209), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1208), .A2(new_n802), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n766), .A2(new_n513), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n757), .A2(G107), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n773), .A2(G283), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n762), .A2(G58), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .A4(new_n1028), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n844), .B(new_n570), .C1(new_n219), .C2(new_n769), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1222), .A2(KEYINPUT119), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1217), .B(new_n1224), .C1(KEYINPUT119), .C2(new_n1222), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n705), .B2(new_n786), .C1(new_n519), .C2(new_n847), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT58), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n570), .B1(new_n844), .B2(new_n256), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1226), .A2(new_n1227), .B1(new_n201), .B2(new_n1228), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT120), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(G132), .A2(new_n765), .B1(new_n755), .B2(G137), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n1167), .B2(new_n758), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n768), .A2(new_n1165), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT121), .Z(new_n1234));
  OAI22_X1  g1034(.A1(new_n786), .A2(new_n1162), .B1(new_n1066), .B2(new_n779), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1232), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT59), .ZN(new_n1237));
  AOI21_X1  g1037(.A(G33), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(G41), .B1(new_n773), .B2(G124), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1238), .B(new_n1239), .C1(new_n349), .C2(new_n763), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n1226), .A2(new_n1227), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n795), .B1(new_n1230), .B2(new_n1242), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1243), .B(new_n800), .C1(G50), .C2(new_n865), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1216), .A2(new_n1244), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1215), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1214), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(KEYINPUT123), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1215), .A2(new_n1245), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n711), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1249), .B1(new_n1250), .B2(new_n1213), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT123), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1248), .A2(new_n1253), .ZN(G375));
  NAND3_X1  g1054(.A1(new_n1155), .A2(new_n1153), .A3(new_n1146), .ZN(new_n1255));
  XOR2_X1   g1055(.A(new_n991), .B(KEYINPUT124), .Z(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1151), .A2(new_n1255), .A3(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n847), .A2(new_n478), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n789), .A2(new_n758), .B1(new_n786), .B2(new_n1076), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1259), .B(new_n1260), .C1(G303), .C2(new_n773), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n765), .A2(new_n548), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n281), .B1(new_n778), .B2(new_n337), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n762), .A2(G77), .B1(G97), .B2(new_n768), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .A4(new_n1264), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1220), .B1(new_n774), .B2(new_n1167), .C1(new_n786), .C2(new_n852), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(G137), .B2(new_n757), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n755), .A2(G150), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n765), .A2(new_n1165), .B1(G50), .B2(new_n778), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1267), .A2(new_n808), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n769), .A2(new_n349), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1265), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n795), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1273), .B(new_n800), .C1(new_n802), .C2(new_n872), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(new_n203), .B2(new_n864), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(new_n1188), .B2(new_n799), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1258), .A2(new_n1276), .ZN(G381));
  NAND3_X1  g1077(.A1(new_n1248), .A2(new_n1186), .A3(new_n1253), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1278), .A2(G381), .ZN(new_n1279));
  INV_X1    g1079(.A(G384), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1100), .A2(new_n1101), .A3(new_n1122), .ZN(new_n1281));
  NOR3_X1   g1081(.A1(G387), .A2(G396), .A3(G393), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .A4(new_n1282), .ZN(G407));
  OAI211_X1 g1083(.A(G407), .B(G213), .C1(G343), .C2(new_n1278), .ZN(G409));
  AND3_X1   g1084(.A1(new_n1023), .A2(KEYINPUT112), .A3(new_n1052), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT112), .B1(new_n1023), .B2(new_n1052), .ZN(new_n1286));
  OAI211_X1 g1086(.A(KEYINPUT126), .B(new_n1281), .C1(new_n1285), .C2(new_n1286), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(G393), .B(G396), .ZN(new_n1288));
  AOI21_X1  g1088(.A(G390), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT126), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1053), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1290), .B1(new_n1291), .B2(G390), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1287), .B(new_n1288), .C1(new_n1289), .C2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1288), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1281), .A2(new_n1053), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1291), .A2(G390), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1294), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1293), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n672), .A2(G343), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1300), .B1(new_n1247), .B2(G378), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT125), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT60), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1151), .B(new_n710), .C1(new_n1255), .C2(new_n1303), .ZN(new_n1304));
  AND2_X1   g1104(.A1(new_n1255), .A2(new_n1303), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1276), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  OR2_X1    g1106(.A1(new_n1306), .A2(new_n1280), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1280), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1190), .A2(new_n1207), .A3(new_n1209), .A4(new_n1257), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1186), .A2(new_n1246), .A3(new_n1311), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1301), .A2(new_n1302), .A3(new_n1310), .A4(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1300), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1314), .B(new_n1312), .C1(new_n1251), .C2(new_n1186), .ZN(new_n1315));
  OAI21_X1  g1115(.A(KEYINPUT125), .B1(new_n1315), .B2(new_n1309), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT62), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1313), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1300), .A2(G2897), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1307), .A2(new_n1308), .A3(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1319), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT61), .B1(new_n1322), .B2(new_n1315), .ZN(new_n1323));
  OAI21_X1  g1123(.A(KEYINPUT62), .B1(new_n1315), .B2(new_n1309), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1299), .B1(new_n1318), .B2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1313), .A2(new_n1316), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT63), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1301), .A2(KEYINPUT63), .A3(new_n1310), .A4(new_n1312), .ZN(new_n1330));
  AND2_X1   g1130(.A1(new_n1323), .A2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1329), .A2(new_n1298), .A3(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1326), .A2(new_n1332), .ZN(G405));
  NAND2_X1  g1133(.A1(new_n1298), .A2(KEYINPUT127), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT127), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1293), .A2(new_n1297), .A3(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1247), .A2(G378), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1278), .A2(new_n1310), .A3(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1310), .B1(new_n1278), .B2(new_n1337), .ZN(new_n1340));
  OAI211_X1 g1140(.A(new_n1334), .B(new_n1336), .C1(new_n1339), .C2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1340), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1342), .A2(KEYINPUT127), .A3(new_n1298), .A4(new_n1338), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1341), .A2(new_n1343), .ZN(G402));
endmodule


