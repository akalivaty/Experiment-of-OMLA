//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 1 1 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n791, new_n792, new_n793,
    new_n794, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G8gat), .ZN(new_n206));
  XOR2_X1   g005(.A(G57gat), .B(G64gat), .Z(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(KEYINPUT96), .B2(KEYINPUT9), .ZN(new_n208));
  NOR2_X1   g007(.A1(G71gat), .A2(G78gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G71gat), .A2(G78gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n209), .B1(KEYINPUT96), .B2(new_n210), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n208), .B(new_n211), .C1(KEYINPUT96), .C2(new_n210), .ZN(new_n212));
  INV_X1    g011(.A(G64gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G57gat), .ZN(new_n214));
  XOR2_X1   g013(.A(KEYINPUT97), .B(G57gat), .Z(new_n215));
  OAI21_X1  g014(.A(new_n214), .B1(new_n215), .B2(new_n213), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n209), .A2(KEYINPUT9), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(new_n210), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n212), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n206), .B1(new_n221), .B2(KEYINPUT21), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(KEYINPUT101), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n221), .A2(KEYINPUT21), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n223), .B(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G231gat), .A2(G233gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G183gat), .B(G211gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g031(.A(G127gat), .B(G155gat), .Z(new_n233));
  XNOR2_X1  g032(.A(new_n233), .B(KEYINPUT20), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n232), .B(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n227), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n227), .A2(new_n235), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT102), .ZN(new_n239));
  XOR2_X1   g038(.A(KEYINPUT92), .B(G29gat), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G36gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(G43gat), .A2(G50gat), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(G43gat), .A2(G50gat), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT15), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT14), .ZN(new_n247));
  INV_X1    g046(.A(G29gat), .ZN(new_n248));
  INV_X1    g047(.A(G36gat), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n247), .A2(new_n248), .A3(new_n249), .A4(KEYINPUT94), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT94), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n243), .A2(KEYINPUT15), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT93), .B(G50gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n255), .B1(new_n256), .B2(G43gat), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n246), .A2(new_n250), .A3(new_n254), .A4(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT91), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n251), .A2(new_n259), .A3(new_n253), .ZN(new_n260));
  OAI211_X1 g059(.A(KEYINPUT91), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n241), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n245), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n239), .B1(new_n265), .B2(KEYINPUT17), .ZN(new_n266));
  NAND2_X1  g065(.A1(G85gat), .A2(G92gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT7), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT8), .ZN(new_n269));
  AND2_X1   g068(.A1(G99gat), .A2(G106gat), .ZN(new_n270));
  OAI221_X1 g069(.A(new_n268), .B1(new_n269), .B2(new_n270), .C1(G85gat), .C2(G92gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(G99gat), .A2(G106gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n271), .B(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT17), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n275), .B1(new_n274), .B2(KEYINPUT102), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n266), .A2(new_n274), .B1(new_n276), .B2(new_n265), .ZN(new_n277));
  NAND3_X1  g076(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT104), .ZN(new_n280));
  XOR2_X1   g079(.A(G190gat), .B(G218gat), .Z(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT103), .ZN(new_n282));
  OAI22_X1  g081(.A1(new_n277), .A2(new_n279), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n280), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G134gat), .B(G162gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  OR2_X1    g088(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n283), .A2(new_n289), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n238), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G15gat), .B(G43gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(G71gat), .B(G99gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT27), .B(G183gat), .ZN(new_n298));
  INV_X1    g097(.A(G190gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT28), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(G169gat), .A2(G176gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  XOR2_X1   g105(.A(new_n306), .B(KEYINPUT26), .Z(new_n307));
  OAI211_X1 g106(.A(new_n302), .B(new_n303), .C1(new_n305), .C2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT24), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n309), .B1(new_n310), .B2(new_n303), .ZN(new_n311));
  NAND3_X1  g110(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n306), .A2(KEYINPUT23), .B1(new_n304), .B2(KEYINPUT65), .ZN(new_n314));
  OR2_X1    g113(.A1(new_n304), .A2(KEYINPUT65), .ZN(new_n315));
  OR2_X1    g114(.A1(new_n306), .A2(KEYINPUT23), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n313), .A2(new_n314), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  OR2_X1    g116(.A1(new_n312), .A2(KEYINPUT64), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(KEYINPUT64), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(new_n311), .A3(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n305), .A2(KEYINPUT25), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT23), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n316), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n317), .A2(KEYINPUT25), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n308), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G113gat), .B(G120gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT67), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT67), .ZN(new_n328));
  INV_X1    g127(.A(G113gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n329), .A2(G120gat), .ZN(new_n330));
  INV_X1    g129(.A(G120gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n331), .A2(G113gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n328), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G134gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(G127gat), .ZN(new_n335));
  INV_X1    g134(.A(G127gat), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT1), .B1(new_n336), .B2(G134gat), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n327), .A2(new_n333), .A3(new_n335), .A4(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n335), .A2(KEYINPUT66), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT66), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n340), .A2(new_n334), .A3(G127gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n336), .A2(G134gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT1), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(new_n330), .B2(new_n332), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n338), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n325), .A2(KEYINPUT68), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G227gat), .ZN(new_n349));
  INV_X1    g148(.A(G233gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n308), .A2(new_n324), .ZN(new_n352));
  OR2_X1    g151(.A1(new_n347), .A2(KEYINPUT68), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n347), .A2(KEYINPUT68), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n348), .A2(new_n351), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT33), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n297), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(KEYINPUT32), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n356), .B(KEYINPUT32), .C1(new_n357), .C2(new_n297), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n351), .B1(new_n348), .B2(new_n355), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT34), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI211_X1 g164(.A(KEYINPUT34), .B(new_n351), .C1(new_n348), .C2(new_n355), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT70), .B1(new_n362), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT70), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n367), .A2(new_n360), .A3(new_n370), .A4(new_n361), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT71), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n367), .B1(new_n361), .B2(new_n360), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n369), .A2(KEYINPUT71), .A3(new_n371), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n374), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G228gat), .A2(G233gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(G211gat), .B(G218gat), .Z(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT72), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n383));
  OR2_X1    g182(.A1(G197gat), .A2(G204gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(G197gat), .A2(G204gat), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n382), .B(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT73), .B(KEYINPUT29), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT87), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT3), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(new_n391), .B2(new_n390), .ZN(new_n393));
  INV_X1    g192(.A(G155gat), .ZN(new_n394));
  INV_X1    g193(.A(G162gat), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT2), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(G141gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n397), .A2(G148gat), .ZN(new_n398));
  INV_X1    g197(.A(G148gat), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n399), .A2(G141gat), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n396), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT76), .B1(new_n398), .B2(new_n400), .ZN(new_n402));
  AND2_X1   g201(.A1(G155gat), .A2(G162gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(G155gat), .A2(G162gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n401), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  XOR2_X1   g206(.A(G141gat), .B(G148gat), .Z(new_n408));
  OAI211_X1 g207(.A(new_n408), .B(new_n396), .C1(KEYINPUT76), .C2(new_n405), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n387), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n407), .A2(new_n409), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT3), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n412), .B1(new_n416), .B2(new_n388), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n380), .B1(new_n411), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G22gat), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n414), .B1(new_n412), .B2(KEYINPUT29), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n410), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n422), .A2(new_n380), .A3(new_n417), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n419), .A2(KEYINPUT88), .A3(new_n420), .A4(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G78gat), .B(G106gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT31), .B(G50gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(KEYINPUT86), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n423), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n418), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n420), .ZN(new_n432));
  OAI21_X1  g231(.A(G22gat), .B1(new_n418), .B2(new_n430), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT88), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n427), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n436), .B1(new_n431), .B2(new_n420), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n429), .A2(new_n435), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n378), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT78), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n440), .B1(new_n410), .B2(new_n347), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n337), .A2(new_n335), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n442), .B1(KEYINPUT67), .B2(new_n326), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n443), .A2(new_n333), .B1(new_n345), .B2(new_n343), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n444), .A2(KEYINPUT78), .A3(new_n413), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(KEYINPUT4), .A3(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n447));
  NAND2_X1  g246(.A1(G225gat), .A2(G233gat), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n410), .A2(KEYINPUT3), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n451), .A2(new_n347), .A3(new_n415), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n452), .A2(KEYINPUT4), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n410), .A2(new_n347), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n446), .B(new_n450), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT4), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n441), .A2(new_n457), .A3(new_n445), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT4), .B1(new_n410), .B2(new_n347), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT77), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT77), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n461), .B(KEYINPUT4), .C1(new_n410), .C2(new_n347), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n458), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n452), .A2(new_n448), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n444), .A2(new_n413), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n466), .B1(new_n441), .B2(new_n445), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT79), .B1(new_n467), .B2(new_n448), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n410), .A2(new_n347), .ZN(new_n469));
  AND4_X1   g268(.A1(KEYINPUT78), .A2(new_n413), .A3(new_n346), .A4(new_n338), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT78), .B1(new_n444), .B2(new_n413), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT79), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n473), .A3(new_n449), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n465), .A2(new_n447), .A3(new_n468), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT81), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n468), .A2(new_n474), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT81), .ZN(new_n478));
  INV_X1    g277(.A(new_n447), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n479), .B1(new_n463), .B2(new_n464), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n477), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n456), .B1(new_n476), .B2(new_n481), .ZN(new_n482));
  XOR2_X1   g281(.A(G57gat), .B(G85gat), .Z(new_n483));
  XNOR2_X1  g282(.A(G1gat), .B(G29gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n486));
  XOR2_X1   g285(.A(new_n485), .B(new_n486), .Z(new_n487));
  NOR2_X1   g286(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT6), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n475), .A2(KEYINPUT81), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n478), .B1(new_n477), .B2(new_n480), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n487), .B(new_n455), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n489), .B1(new_n488), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g294(.A1(G226gat), .A2(G233gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n352), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n388), .B1(new_n308), .B2(new_n324), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n497), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT74), .B1(new_n499), .B2(new_n412), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n325), .A2(KEYINPUT29), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n497), .B(new_n387), .C1(new_n501), .C2(new_n496), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n499), .A2(new_n412), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n500), .B1(new_n504), .B2(KEYINPUT74), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G8gat), .B(G36gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(G64gat), .B(G92gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n509), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n505), .A2(KEYINPUT30), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT75), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n505), .A2(new_n511), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT30), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI211_X1 g315(.A(KEYINPUT75), .B(KEYINPUT30), .C1(new_n505), .C2(new_n511), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n510), .B(new_n512), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n518), .A2(KEYINPUT35), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n439), .A2(new_n495), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n518), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT84), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n455), .B1(new_n490), .B2(new_n491), .ZN(new_n524));
  INV_X1    g323(.A(new_n487), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT83), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n526), .A2(new_n494), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n524), .A2(KEYINPUT83), .A3(new_n525), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n523), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT83), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(new_n482), .B2(new_n487), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT6), .B1(new_n482), .B2(new_n487), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n528), .A2(new_n531), .A3(new_n532), .A4(new_n523), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n489), .ZN(new_n534));
  OAI211_X1 g333(.A(KEYINPUT85), .B(new_n522), .C1(new_n529), .C2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n528), .A2(new_n531), .A3(new_n532), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT84), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n538), .A2(new_n489), .A3(new_n533), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT85), .B1(new_n539), .B2(new_n522), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n429), .A2(new_n435), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n437), .A2(new_n433), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n375), .B(KEYINPUT69), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n543), .A2(new_n372), .A3(new_n544), .ZN(new_n545));
  NOR3_X1   g344(.A1(new_n536), .A2(new_n540), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT35), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n521), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n446), .B1(new_n453), .B2(new_n454), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n549), .A2(new_n449), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT39), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n525), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT39), .B1(new_n472), .B2(new_n449), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n552), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT40), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n554), .A2(new_n555), .ZN(new_n557));
  NOR3_X1   g356(.A1(new_n556), .A2(new_n557), .A3(new_n488), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(new_n518), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT37), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n511), .B1(new_n505), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n497), .B1(new_n501), .B2(new_n496), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n562), .A2(KEYINPUT89), .A3(new_n412), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n563), .B1(new_n499), .B2(new_n412), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT89), .B1(new_n562), .B2(new_n412), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT37), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT38), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n561), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n506), .A2(KEYINPUT37), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n569), .A2(new_n561), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n514), .B(new_n568), .C1(new_n570), .C2(new_n567), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n559), .B(new_n543), .C1(new_n495), .C2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n544), .A2(KEYINPUT36), .A3(new_n372), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n369), .A2(KEYINPUT71), .A3(new_n371), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT71), .B1(new_n369), .B2(new_n371), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n574), .A2(new_n575), .A3(new_n375), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n573), .B1(new_n576), .B2(KEYINPUT36), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n536), .A2(new_n540), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n572), .B(new_n577), .C1(new_n578), .C2(new_n543), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n294), .B1(new_n548), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n206), .A2(KEYINPUT17), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n581), .B(new_n265), .Z(new_n582));
  NAND2_X1  g381(.A1(G229gat), .A2(G233gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT18), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT95), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n265), .B(new_n206), .Z(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n583), .B(KEYINPUT13), .ZN(new_n590));
  OAI22_X1  g389(.A1(new_n584), .A2(new_n585), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G113gat), .B(G141gat), .ZN(new_n592));
  INV_X1    g391(.A(G197gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT11), .B(G169gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT90), .B(KEYINPUT12), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n591), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n587), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n586), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n598), .B1(new_n601), .B2(new_n591), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G230gat), .A2(G233gat), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n274), .A2(new_n220), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT105), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n274), .A2(new_n220), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n274), .A2(KEYINPUT105), .A3(new_n220), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT10), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n606), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n605), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n609), .A2(new_n610), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n614), .B1(new_n605), .B2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G120gat), .B(G148gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n604), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n580), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n539), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n518), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT106), .B(KEYINPUT16), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G8gat), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n629), .A2(KEYINPUT42), .A3(new_n631), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n629), .A2(new_n631), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT42), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n634), .B1(new_n629), .B2(G8gat), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n632), .B1(new_n633), .B2(new_n635), .ZN(G1325gat));
  INV_X1    g435(.A(G15gat), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n624), .A2(new_n637), .A3(new_n577), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n625), .A2(new_n576), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n638), .B1(new_n637), .B2(new_n639), .ZN(G1326gat));
  NOR2_X1   g439(.A1(new_n624), .A2(new_n543), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT43), .B(G22gat), .Z(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(G1327gat));
  INV_X1    g442(.A(new_n623), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(new_n238), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n522), .B1(new_n529), .B2(new_n534), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT85), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n544), .A2(new_n372), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n438), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n648), .A2(new_n535), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n520), .B1(new_n651), .B2(KEYINPUT35), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n572), .A2(new_n577), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n648), .A2(new_n535), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n653), .B1(new_n654), .B2(new_n438), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n292), .B(new_n645), .C1(new_n652), .C2(new_n655), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n656), .A2(new_n539), .A3(new_n240), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n657), .B(KEYINPUT45), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n292), .B(KEYINPUT107), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n659), .B1(new_n652), .B2(new_n655), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n238), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI211_X1 g461(.A(KEYINPUT44), .B(new_n292), .C1(new_n652), .C2(new_n655), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n662), .A2(new_n623), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n240), .B1(new_n664), .B2(new_n539), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n658), .A2(new_n665), .ZN(G1328gat));
  NOR3_X1   g465(.A1(new_n656), .A2(G36gat), .A3(new_n522), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT46), .ZN(new_n668));
  OAI21_X1  g467(.A(G36gat), .B1(new_n664), .B2(new_n522), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(G1329gat));
  OAI21_X1  g469(.A(G43gat), .B1(new_n664), .B2(new_n577), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n378), .A2(G43gat), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  OR3_X1    g472(.A1(new_n656), .A2(KEYINPUT109), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT109), .B1(new_n656), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT47), .B1(new_n676), .B2(KEYINPUT108), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n671), .B(new_n676), .C1(KEYINPUT108), .C2(KEYINPUT47), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(G1330gat));
  OR2_X1    g480(.A1(new_n656), .A2(KEYINPUT110), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n543), .B1(new_n656), .B2(KEYINPUT110), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n256), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT48), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n438), .A2(new_n256), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n685), .B(new_n686), .C1(new_n664), .C2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n664), .A2(new_n687), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT48), .B1(new_n689), .B2(new_n684), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(G1331gat));
  INV_X1    g490(.A(new_n622), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n603), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n580), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n626), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(new_n215), .ZN(G1332gat));
  AOI21_X1  g496(.A(new_n522), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT111), .B(KEYINPUT112), .ZN(new_n700));
  NOR2_X1   g499(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n699), .B(new_n702), .ZN(G1333gat));
  INV_X1    g502(.A(new_n577), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n695), .A2(G71gat), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(G71gat), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(new_n694), .B2(new_n378), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g508(.A1(new_n695), .A2(new_n438), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g510(.A1(new_n662), .A2(new_n663), .ZN(new_n712));
  INV_X1    g511(.A(new_n693), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n712), .A2(new_n539), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(G85gat), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n548), .A2(new_n579), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT51), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n238), .A2(new_n603), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n716), .A2(new_n717), .A3(new_n292), .A4(new_n718), .ZN(new_n719));
  OAI211_X1 g518(.A(new_n292), .B(new_n718), .C1(new_n652), .C2(new_n655), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT51), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n626), .A2(new_n715), .A3(new_n622), .ZN(new_n723));
  OAI22_X1  g522(.A1(new_n714), .A2(new_n715), .B1(new_n722), .B2(new_n723), .ZN(G1336gat));
  INV_X1    g523(.A(KEYINPUT113), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n719), .A2(new_n721), .B1(new_n725), .B2(new_n720), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n720), .A2(new_n725), .A3(new_n717), .ZN(new_n727));
  OR3_X1    g526(.A1(new_n522), .A2(G92gat), .A3(new_n692), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n662), .A2(new_n518), .A3(new_n663), .A4(new_n693), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n730), .A2(G92gat), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT52), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(G92gat), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT52), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n733), .B(new_n734), .C1(new_n722), .C2(new_n728), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(G1337gat));
  NOR3_X1   g535(.A1(new_n712), .A2(new_n577), .A3(new_n713), .ZN(new_n737));
  INV_X1    g536(.A(G99gat), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n576), .A2(new_n738), .A3(new_n622), .ZN(new_n739));
  OAI22_X1  g538(.A1(new_n737), .A2(new_n738), .B1(new_n722), .B2(new_n739), .ZN(G1338gat));
  OR3_X1    g539(.A1(new_n543), .A2(new_n692), .A3(G106gat), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n726), .A2(new_n727), .A3(new_n741), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n662), .A2(new_n438), .A3(new_n663), .A4(new_n693), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n743), .A2(G106gat), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT53), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(G106gat), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT53), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n746), .B(new_n747), .C1(new_n722), .C2(new_n741), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(G1339gat));
  INV_X1    g548(.A(new_n238), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT54), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n751), .B(new_n605), .C1(new_n611), .C2(new_n613), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n752), .A2(KEYINPUT114), .A3(new_n619), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT114), .B1(new_n752), .B2(new_n619), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n611), .A2(new_n605), .A3(new_n613), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n614), .A2(KEYINPUT54), .ZN(new_n756));
  OAI22_X1  g555(.A1(new_n753), .A2(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n620), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI211_X1 g560(.A(KEYINPUT115), .B(new_n620), .C1(new_n757), .C2(new_n758), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n757), .A2(new_n758), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n761), .A2(new_n603), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n582), .A2(new_n583), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n765), .A2(KEYINPUT116), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(KEYINPUT116), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n589), .A2(new_n590), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  AOI22_X1  g568(.A1(new_n596), .A2(new_n769), .B1(new_n587), .B2(new_n599), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n622), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n659), .B1(new_n764), .B2(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n761), .A2(new_n770), .A3(new_n762), .A4(new_n763), .ZN(new_n773));
  INV_X1    g572(.A(new_n659), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n750), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n604), .A2(new_n692), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n294), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n539), .A2(new_n518), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n782), .A2(new_n650), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n783), .A2(new_n329), .A3(new_n603), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n439), .ZN(new_n785));
  OAI21_X1  g584(.A(G113gat), .B1(new_n785), .B2(new_n604), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(G1340gat));
  NAND3_X1  g586(.A1(new_n783), .A2(new_n331), .A3(new_n622), .ZN(new_n788));
  OAI21_X1  g587(.A(G120gat), .B1(new_n785), .B2(new_n692), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(G1341gat));
  NOR3_X1   g589(.A1(new_n785), .A2(new_n336), .A3(new_n750), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n783), .A2(new_n238), .ZN(new_n792));
  OR2_X1    g591(.A1(new_n792), .A2(KEYINPUT117), .ZN(new_n793));
  AOI21_X1  g592(.A(G127gat), .B1(new_n792), .B2(KEYINPUT117), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n791), .B1(new_n793), .B2(new_n794), .ZN(G1342gat));
  NAND3_X1  g594(.A1(new_n783), .A2(new_n334), .A3(new_n292), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n796), .A2(KEYINPUT56), .ZN(new_n797));
  OAI21_X1  g596(.A(G134gat), .B1(new_n785), .B2(new_n293), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(KEYINPUT56), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(G1343gat));
  OR2_X1    g599(.A1(new_n773), .A2(new_n774), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n763), .A2(new_n603), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n771), .B1(new_n802), .B2(new_n759), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n293), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n238), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  OAI211_X1 g604(.A(KEYINPUT57), .B(new_n438), .C1(new_n805), .C2(new_n778), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n543), .B1(new_n776), .B2(new_n779), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n806), .B1(new_n807), .B2(KEYINPUT57), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n577), .A2(new_n781), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT118), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(G141gat), .B1(new_n811), .B2(new_n604), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n704), .A2(new_n543), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT119), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n782), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n603), .A2(new_n397), .ZN(new_n816));
  XOR2_X1   g615(.A(new_n816), .B(KEYINPUT120), .Z(new_n817));
  INV_X1    g616(.A(KEYINPUT121), .ZN(new_n818));
  AOI22_X1  g617(.A1(new_n815), .A2(new_n817), .B1(new_n818), .B2(KEYINPUT58), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n818), .A2(KEYINPUT58), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n812), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n820), .B1(new_n812), .B2(new_n819), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(G1344gat));
  NAND3_X1  g622(.A1(new_n815), .A2(new_n399), .A3(new_n622), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n811), .A2(new_n692), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n825), .A2(KEYINPUT59), .A3(new_n399), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n438), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n773), .A2(new_n293), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n238), .B1(new_n830), .B2(new_n804), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n778), .B(KEYINPUT123), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n829), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n833), .B1(new_n807), .B2(new_n827), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n810), .A2(new_n622), .ZN(new_n835));
  OAI21_X1  g634(.A(G148gat), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g635(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n824), .B1(new_n826), .B2(new_n838), .ZN(G1345gat));
  NOR3_X1   g638(.A1(new_n811), .A2(new_n394), .A3(new_n750), .ZN(new_n840));
  AOI21_X1  g639(.A(G155gat), .B1(new_n815), .B2(new_n238), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(G1346gat));
  OAI21_X1  g641(.A(G162gat), .B1(new_n811), .B2(new_n774), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n815), .A2(new_n395), .A3(new_n292), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT124), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT124), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n843), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(G1347gat));
  NAND2_X1  g648(.A1(new_n780), .A2(new_n539), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT125), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n522), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n780), .A2(KEYINPUT125), .A3(new_n539), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n650), .A3(new_n853), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n854), .A2(G169gat), .A3(new_n604), .ZN(new_n855));
  INV_X1    g654(.A(G169gat), .ZN(new_n856));
  INV_X1    g655(.A(new_n439), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n850), .A2(new_n522), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n856), .B1(new_n858), .B2(new_n603), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n855), .A2(new_n859), .ZN(G1348gat));
  OR2_X1    g659(.A1(new_n854), .A2(new_n692), .ZN(new_n861));
  INV_X1    g660(.A(G176gat), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n692), .A2(new_n862), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n861), .A2(new_n862), .B1(new_n858), .B2(new_n863), .ZN(G1349gat));
  NAND2_X1  g663(.A1(new_n858), .A2(new_n238), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(G183gat), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n238), .A2(new_n298), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n854), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT60), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT60), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n866), .B(new_n870), .C1(new_n854), .C2(new_n867), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(G1350gat));
  NAND2_X1  g671(.A1(new_n858), .A2(new_n292), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(G190gat), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n874), .A2(KEYINPUT61), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n874), .A2(KEYINPUT61), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n659), .A2(new_n299), .ZN(new_n877));
  OAI22_X1  g676(.A1(new_n875), .A2(new_n876), .B1(new_n854), .B2(new_n877), .ZN(G1351gat));
  AND3_X1   g677(.A1(new_n852), .A2(new_n813), .A3(new_n853), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n593), .A3(new_n603), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n577), .A2(new_n539), .A3(new_n518), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n834), .A2(KEYINPUT126), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT126), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n833), .B(new_n883), .C1(new_n807), .C2(new_n827), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n881), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(new_n603), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n880), .B1(new_n886), .B2(new_n593), .ZN(G1352gat));
  NOR2_X1   g686(.A1(new_n692), .A2(G204gat), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n852), .A2(new_n813), .A3(new_n853), .A4(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n889), .B(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n882), .A2(new_n884), .ZN(new_n892));
  INV_X1    g691(.A(new_n881), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n892), .A2(KEYINPUT127), .A3(new_n622), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(G204gat), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT127), .B1(new_n885), .B2(new_n622), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n891), .B1(new_n895), .B2(new_n896), .ZN(G1353gat));
  INV_X1    g696(.A(G211gat), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n879), .A2(new_n898), .A3(new_n238), .ZN(new_n899));
  OR3_X1    g698(.A1(new_n834), .A2(new_n750), .A3(new_n881), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n900), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT63), .B1(new_n900), .B2(G211gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(G1354gat));
  AOI21_X1  g702(.A(G218gat), .B1(new_n879), .B2(new_n659), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n292), .A2(G218gat), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n885), .B2(new_n905), .ZN(G1355gat));
endmodule


