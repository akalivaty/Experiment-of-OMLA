//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n556, new_n558, new_n559, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1154;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  XNOR2_X1  g032(.A(G325), .B(KEYINPUT66), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(new_n455), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  AND3_X1   g037(.A1(KEYINPUT68), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(KEYINPUT3), .B1(KEYINPUT68), .B2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT67), .B(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(G137), .A3(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n476), .A2(G125), .ZN(new_n477));
  AND2_X1   g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  OAI221_X1 g056(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n467), .C2(G112), .ZN(new_n482));
  OR2_X1    g057(.A1(new_n482), .A2(KEYINPUT69), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(KEYINPUT69), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n465), .A2(G2105), .ZN(new_n485));
  AOI22_X1  g060(.A1(new_n483), .A2(new_n484), .B1(G136), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(G124), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n465), .A2(new_n467), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n486), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  OAI22_X1  g066(.A1(new_n463), .A2(new_n464), .B1(new_n473), .B2(new_n474), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT4), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n496));
  AND2_X1   g071(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n497));
  NOR2_X1   g072(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n495), .B1(new_n499), .B2(new_n475), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n467), .A2(new_n476), .A3(KEYINPUT70), .A4(new_n496), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n494), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(G126), .B1(new_n463), .B2(new_n464), .ZN(new_n503));
  NAND2_X1  g078(.A1(G114), .A2(G2104), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G2105), .B1(G102), .B2(new_n470), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n502), .A2(KEYINPUT71), .A3(new_n506), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(G164));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G62), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n512), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  XOR2_X1   g095(.A(new_n520), .B(KEYINPUT72), .Z(new_n521));
  INV_X1    g096(.A(new_n517), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT6), .B(G651), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n524), .A2(G88), .B1(G50), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n521), .A2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NAND3_X1  g104(.A1(new_n522), .A2(G63), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT73), .B(G51), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n525), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT74), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n524), .A2(G89), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  AOI22_X1  g113(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G651), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n522), .A2(new_n523), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  INV_X1    g118(.A(G52), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n542), .A2(new_n543), .B1(new_n525), .B2(new_n544), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n541), .A2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  AOI22_X1  g122(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n540), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(KEYINPUT75), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n524), .A2(G81), .B1(G43), .B2(new_n526), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n549), .A2(KEYINPUT75), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OR3_X1    g136(.A1(new_n525), .A2(KEYINPUT9), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT9), .B1(new_n525), .B2(new_n561), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT76), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n522), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G91), .ZN(new_n567));
  OAI22_X1  g142(.A1(new_n566), .A2(new_n540), .B1(new_n542), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT76), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n562), .A2(new_n570), .A3(new_n563), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n565), .A2(new_n569), .A3(new_n571), .ZN(G299));
  NAND2_X1  g147(.A1(new_n524), .A2(G87), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n526), .A2(G49), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  INV_X1    g151(.A(KEYINPUT77), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n522), .A2(new_n577), .A3(G61), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT77), .B1(new_n517), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G651), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n524), .A2(G86), .B1(G48), .B2(new_n526), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G305));
  AOI22_X1  g160(.A1(new_n524), .A2(G85), .B1(G47), .B2(new_n526), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n540), .B2(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n524), .A2(G92), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT10), .ZN(new_n591));
  XNOR2_X1  g166(.A(KEYINPUT78), .B(G66), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n522), .A2(new_n592), .B1(G79), .B2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G54), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n593), .A2(new_n540), .B1(new_n594), .B2(new_n525), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n589), .B1(new_n596), .B2(G868), .ZN(G284));
  OAI21_X1  g172(.A(new_n589), .B1(new_n596), .B2(G868), .ZN(G321));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(G299), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(G168), .B2(new_n599), .ZN(G297));
  OAI21_X1  g176(.A(new_n600), .B1(G168), .B2(new_n599), .ZN(G280));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n596), .B1(new_n603), .B2(G860), .ZN(G148));
  INV_X1    g179(.A(new_n596), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(G559), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n606), .A2(new_n599), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n608), .B(KEYINPUT79), .C1(G868), .C2(new_n554), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(KEYINPUT79), .B2(new_n608), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT80), .Z(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n488), .A2(G123), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n485), .A2(G135), .ZN(new_n614));
  OAI221_X1 g189(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n467), .C2(G111), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(G2096), .Z(new_n617));
  NAND2_X1  g192(.A1(new_n476), .A2(new_n470), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(KEYINPUT13), .B(G2100), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n617), .A2(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(G2451), .B(G2454), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2427), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT15), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n628), .A2(G2435), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(G2435), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(KEYINPUT14), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G2443), .B(G2446), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n633), .A2(new_n637), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n625), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n642), .A2(new_n624), .A3(new_n638), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n641), .A2(new_n643), .A3(G14), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT83), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT83), .ZN(new_n646));
  NAND4_X1  g221(.A1(new_n641), .A2(new_n643), .A3(new_n646), .A4(G14), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(G401));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2067), .B(G2678), .Z(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(new_n654), .A3(KEYINPUT17), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT18), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n653), .B2(KEYINPUT18), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2096), .B(G2100), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT84), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n660), .B(new_n662), .ZN(G227));
  XNOR2_X1  g238(.A(G1961), .B(G1966), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT85), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  AND2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n665), .A2(new_n666), .ZN(new_n672));
  AOI22_X1  g247(.A1(new_n670), .A2(new_n671), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  OR3_X1    g248(.A1(new_n667), .A2(new_n672), .A3(new_n669), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n673), .B(new_n674), .C1(new_n671), .C2(new_n670), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  INV_X1    g253(.A(G1981), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n677), .B(new_n681), .ZN(G229));
  NAND2_X1  g257(.A1(G299), .A2(G16), .ZN(new_n683));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n684), .A2(KEYINPUT23), .A3(G20), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT23), .ZN(new_n686));
  INV_X1    g261(.A(G20), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n687), .B2(G16), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n683), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G1956), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT86), .B(G29), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G35), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G162), .B2(new_n693), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT29), .Z(new_n696));
  INV_X1    g271(.A(G2090), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n691), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT96), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  AND2_X1   g276(.A1(KEYINPUT30), .A2(G28), .ZN(new_n702));
  NOR2_X1   g277(.A1(KEYINPUT30), .A2(G28), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT31), .B(G11), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n704), .B(new_n705), .C1(new_n616), .C2(new_n693), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT95), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT24), .B(G34), .Z(new_n708));
  OAI21_X1  g283(.A(KEYINPUT93), .B1(new_n708), .B2(new_n692), .ZN(new_n709));
  OR3_X1    g284(.A1(new_n708), .A2(KEYINPUT93), .A3(new_n692), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n709), .B(new_n710), .C1(new_n480), .C2(new_n701), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT94), .Z(new_n712));
  AOI21_X1  g287(.A(new_n707), .B1(new_n712), .B2(G2084), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n684), .A2(G5), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G171), .B2(new_n684), .ZN(new_n715));
  INV_X1    g290(.A(G1961), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n692), .A2(G27), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G164), .B2(new_n692), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G2078), .ZN(new_n720));
  NOR2_X1   g295(.A1(G29), .A2(G32), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n485), .A2(G141), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n470), .A2(G105), .ZN(new_n723));
  NAND3_X1  g298(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT26), .Z(new_n725));
  NAND3_X1  g300(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n488), .A2(G129), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n721), .B1(new_n728), .B2(G29), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT27), .B(G1996), .Z(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n720), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n700), .A2(new_n713), .A3(new_n717), .A4(new_n732), .ZN(new_n733));
  OR2_X1    g308(.A1(G29), .A2(G33), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT91), .Z(new_n736));
  AOI22_X1  g311(.A1(new_n736), .A2(new_n475), .B1(G139), .B2(new_n485), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT90), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT25), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n734), .B1(new_n741), .B2(new_n701), .ZN(new_n742));
  INV_X1    g317(.A(G2072), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT92), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n485), .A2(G140), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT89), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  OAI221_X1 g323(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n467), .C2(G116), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n488), .A2(G128), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G29), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n693), .A2(KEYINPUT28), .A3(G26), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(KEYINPUT28), .B1(new_n693), .B2(G26), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(G2067), .Z(new_n757));
  NOR2_X1   g332(.A1(G16), .A2(G21), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G168), .B2(G16), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n759), .A2(G1966), .ZN(new_n760));
  NOR4_X1   g335(.A1(new_n733), .A2(new_n745), .A3(new_n757), .A4(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n692), .A2(G25), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n485), .A2(G131), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT87), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  OAI221_X1 g340(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n467), .C2(G107), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n488), .A2(G119), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT88), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n762), .B1(new_n769), .B2(new_n692), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT35), .B(G1991), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  MUX2_X1   g347(.A(G24), .B(G290), .S(G16), .Z(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(G1986), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n684), .A2(G6), .ZN(new_n775));
  INV_X1    g350(.A(G305), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(new_n684), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT32), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(new_n679), .ZN(new_n779));
  NAND2_X1  g354(.A1(G166), .A2(G16), .ZN(new_n780));
  OR2_X1    g355(.A1(G16), .A2(G22), .ZN(new_n781));
  AND3_X1   g356(.A1(new_n780), .A2(G1971), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(G1971), .B1(new_n780), .B2(new_n781), .ZN(new_n783));
  NOR2_X1   g358(.A1(G16), .A2(G23), .ZN(new_n784));
  INV_X1    g359(.A(G288), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(G16), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT33), .B(G1976), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n782), .A2(new_n783), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n779), .A2(KEYINPUT34), .A3(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(KEYINPUT34), .B1(new_n779), .B2(new_n789), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n772), .B(new_n774), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT36), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n729), .A2(new_n730), .ZN(new_n795));
  INV_X1    g370(.A(G1341), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n554), .A2(G16), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G16), .B2(G19), .ZN(new_n798));
  OAI221_X1 g373(.A(new_n795), .B1(new_n759), .B2(G1966), .C1(new_n796), .C2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n796), .ZN(new_n801));
  INV_X1    g376(.A(G1348), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n596), .A2(new_n684), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G4), .B2(new_n684), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n801), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n802), .B2(new_n804), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n761), .A2(new_n794), .A3(new_n800), .A4(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n742), .A2(new_n743), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n712), .A2(G2084), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n696), .A2(new_n697), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  NOR4_X1   g387(.A1(new_n807), .A2(new_n809), .A3(new_n810), .A4(new_n812), .ZN(G311));
  INV_X1    g388(.A(new_n807), .ZN(new_n814));
  INV_X1    g389(.A(new_n810), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n814), .A2(new_n808), .A3(new_n815), .A4(new_n811), .ZN(G150));
  AOI22_X1  g391(.A1(new_n524), .A2(G93), .B1(G55), .B2(new_n526), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n540), .B2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT97), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(G860), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT37), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n821), .A2(new_n553), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n554), .A2(new_n819), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n596), .A2(G559), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n824), .B1(new_n831), .B2(G860), .ZN(G145));
  INV_X1    g407(.A(G37), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n741), .B(new_n728), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n751), .B(new_n507), .Z(new_n835));
  OR2_X1    g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n488), .A2(G130), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n485), .A2(G142), .ZN(new_n839));
  OAI221_X1 g414(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n467), .C2(G118), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n620), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(new_n768), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n768), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT98), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n836), .B(new_n837), .C1(new_n847), .C2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n480), .B(new_n616), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n490), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n834), .A2(new_n835), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n834), .A2(new_n835), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n850), .B(new_n853), .C1(new_n856), .C2(new_n845), .ZN(new_n857));
  INV_X1    g432(.A(new_n847), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n858), .B(new_n848), .C1(new_n854), .C2(new_n855), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n850), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(KEYINPUT99), .B1(new_n860), .B2(new_n852), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n862));
  AOI211_X1 g437(.A(new_n862), .B(new_n853), .C1(new_n850), .C2(new_n859), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n833), .B(new_n857), .C1(new_n861), .C2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g440(.A(G305), .B(G288), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G290), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(G166), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT101), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(KEYINPUT42), .Z(new_n870));
  AND2_X1   g445(.A1(new_n825), .A2(new_n826), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n606), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n596), .B(G299), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n873), .A2(KEYINPUT41), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT100), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n596), .A2(G299), .A3(new_n875), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n876), .B(KEYINPUT41), .C1(new_n873), .C2(new_n875), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n872), .A2(new_n874), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n876), .B1(new_n873), .B2(new_n875), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n879), .B2(new_n872), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n870), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT102), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n870), .A2(new_n880), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n883), .A2(new_n599), .ZN(new_n884));
  AOI22_X1  g459(.A1(new_n882), .A2(new_n884), .B1(new_n599), .B2(new_n821), .ZN(G295));
  AOI22_X1  g460(.A1(new_n882), .A2(new_n884), .B1(new_n599), .B2(new_n821), .ZN(G331));
  INV_X1    g461(.A(new_n868), .ZN(new_n887));
  XNOR2_X1  g462(.A(G286), .B(G301), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n871), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(G286), .B(G171), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n827), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n879), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI22_X1  g469(.A1(new_n874), .A2(new_n877), .B1(new_n889), .B2(new_n891), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n887), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n896), .A2(new_n833), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT41), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n898), .B1(new_n889), .B2(new_n891), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n873), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n900), .B(new_n868), .C1(new_n893), .C2(new_n899), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n897), .A2(KEYINPUT43), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n877), .A2(new_n874), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n892), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n904), .B(new_n868), .C1(new_n893), .C2(new_n892), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n905), .A2(new_n896), .A3(new_n833), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT44), .B1(new_n902), .B2(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n897), .A2(KEYINPUT103), .A3(new_n907), .A4(new_n901), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT103), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n911), .B1(new_n906), .B2(KEYINPUT43), .ZN(new_n912));
  AND4_X1   g487(.A1(new_n907), .A2(new_n901), .A3(new_n833), .A4(new_n896), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n909), .B1(new_n915), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g491(.A(G1384), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT45), .B1(new_n507), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n472), .A2(G40), .A3(new_n479), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n751), .B(G2067), .ZN(new_n922));
  INV_X1    g497(.A(G1996), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n728), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n921), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT106), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n926), .A2(new_n771), .A3(new_n769), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n751), .A2(G2067), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n921), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  XOR2_X1   g504(.A(new_n768), .B(new_n771), .Z(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n921), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n926), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(G290), .A2(G1986), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n921), .A2(new_n933), .ZN(new_n934));
  XOR2_X1   g509(.A(new_n934), .B(KEYINPUT126), .Z(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT48), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n929), .B1(new_n932), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n728), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n921), .B1(new_n922), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT46), .ZN(new_n940));
  INV_X1    g515(.A(new_n921), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n940), .B1(new_n941), .B2(G1996), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n921), .A2(KEYINPUT46), .A3(new_n923), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n939), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  XOR2_X1   g519(.A(new_n944), .B(KEYINPUT125), .Z(new_n945));
  XNOR2_X1  g520(.A(new_n945), .B(KEYINPUT47), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n937), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G8), .ZN(new_n948));
  NOR2_X1   g523(.A1(G168), .A2(new_n948), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n502), .A2(KEYINPUT71), .A3(new_n506), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT71), .B1(new_n502), .B2(new_n506), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n950), .A2(new_n951), .A3(G1384), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT50), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT107), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G2084), .ZN(new_n955));
  AOI21_X1  g530(.A(G1384), .B1(new_n502), .B2(new_n506), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n920), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n509), .A2(new_n917), .A3(new_n510), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n959), .A3(KEYINPUT50), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n954), .A2(new_n955), .A3(new_n957), .A4(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT121), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT111), .B1(new_n918), .B2(new_n920), .ZN(new_n963));
  AND4_X1   g538(.A1(G40), .A2(new_n479), .A3(new_n471), .A4(new_n468), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n964), .B(new_n965), .C1(new_n956), .C2(KEYINPUT45), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n509), .A2(KEYINPUT45), .A3(new_n917), .A4(new_n510), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n963), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1966), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n961), .A2(new_n962), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n962), .B1(new_n961), .B2(new_n970), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n949), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT122), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g550(.A(KEYINPUT122), .B(new_n949), .C1(new_n971), .C2(new_n972), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n961), .A2(new_n970), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(G8), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n949), .A2(KEYINPUT51), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n971), .A2(new_n972), .A3(G286), .ZN(new_n982));
  NAND2_X1  g557(.A1(KEYINPUT51), .A2(G8), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n977), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n954), .A2(new_n957), .A3(new_n960), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n958), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G2078), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n920), .B1(KEYINPUT45), .B2(new_n956), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  AOI22_X1  g568(.A1(new_n987), .A2(new_n716), .B1(new_n988), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n988), .A2(G2078), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n963), .A2(new_n966), .A3(new_n967), .A4(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(G301), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n986), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n917), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n964), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n1000), .B1(new_n989), .B2(new_n958), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1001), .A2(G1971), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n507), .A2(new_n917), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n920), .B1(new_n1003), .B2(KEYINPUT50), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n509), .A2(new_n953), .A3(new_n917), .A4(new_n510), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(KEYINPUT108), .B(G2090), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(G8), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(G303), .A2(G8), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(KEYINPUT109), .A2(KEYINPUT55), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1009), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1007), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n954), .A2(new_n1017), .A3(new_n957), .A4(new_n960), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n990), .A2(new_n992), .ZN(new_n1019));
  INV_X1    g594(.A(G1971), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n948), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  MUX2_X1   g597(.A(new_n1012), .B(new_n1014), .S(new_n1010), .Z(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(KEYINPUT110), .A2(KEYINPUT49), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G305), .A2(G1981), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(KEYINPUT110), .B2(KEYINPUT49), .ZN(new_n1027));
  NOR2_X1   g602(.A1(G305), .A2(G1981), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1003), .A2(new_n920), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1030), .A2(new_n948), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1028), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1032), .A2(KEYINPUT110), .A3(KEYINPUT49), .A4(new_n1026), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1029), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1031), .ZN(new_n1035));
  INV_X1    g610(.A(G1976), .ZN(new_n1036));
  NOR2_X1   g611(.A1(G288), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT52), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT52), .B1(G288), .B2(new_n1036), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1031), .B(new_n1039), .C1(new_n1036), .C2(G288), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1034), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1016), .A2(new_n1024), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1042), .B1(new_n985), .B2(KEYINPUT62), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n998), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT56), .B(G2072), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1001), .A2(new_n1046), .B1(new_n1006), .B2(new_n690), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n568), .A2(KEYINPUT113), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n564), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n568), .A2(KEYINPUT113), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n565), .A2(KEYINPUT57), .A3(new_n569), .A4(new_n571), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1045), .B1(new_n1047), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1006), .A2(new_n690), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n990), .A2(new_n992), .A3(new_n1046), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n1057), .A3(new_n1054), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT114), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1054), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(KEYINPUT118), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1056), .A2(new_n1057), .A3(new_n1054), .A4(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1055), .A2(new_n1059), .A3(new_n1062), .A4(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT117), .B(KEYINPUT61), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n923), .B(new_n992), .C1(new_n952), .C2(KEYINPUT45), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT58), .B(G1341), .Z(new_n1069));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n964), .A2(new_n956), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1070), .B1(new_n964), .B2(new_n956), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1069), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1068), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1068), .A2(KEYINPUT116), .A3(new_n1073), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(new_n554), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT59), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1076), .A2(new_n1077), .A3(new_n1080), .A4(new_n554), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1083), .A2(KEYINPUT61), .A3(new_n1058), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1067), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT119), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1071), .A2(new_n1072), .A3(G2067), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1088), .B1(new_n987), .B2(new_n802), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1089), .A2(KEYINPUT120), .A3(KEYINPUT60), .ZN(new_n1090));
  AOI211_X1 g665(.A(KEYINPUT120), .B(new_n596), .C1(new_n1089), .C2(KEYINPUT60), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n987), .A2(new_n802), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1088), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1092), .A2(KEYINPUT60), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n605), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1090), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1089), .A2(KEYINPUT60), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1067), .A2(new_n1082), .A3(KEYINPUT119), .A4(new_n1084), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1087), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1083), .B1(new_n1089), .B2(new_n605), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1102), .A2(new_n1059), .A3(new_n1064), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n987), .A2(new_n716), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n993), .A2(new_n988), .ZN(new_n1107));
  XOR2_X1   g682(.A(new_n472), .B(KEYINPUT123), .Z(new_n1108));
  AND3_X1   g683(.A1(new_n1108), .A2(G40), .A3(new_n999), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1109), .A2(new_n479), .A3(new_n919), .A4(new_n995), .ZN(new_n1110));
  AND4_X1   g685(.A1(G301), .A2(new_n1106), .A3(new_n1107), .A4(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1105), .B1(new_n1111), .B2(new_n997), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n994), .A2(G301), .A3(new_n996), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1106), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1113), .B(KEYINPUT54), .C1(new_n1114), .C2(G301), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1112), .A2(new_n1042), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n985), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1104), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT124), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1041), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT112), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT63), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1124), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n979), .A2(G286), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1123), .A2(new_n1125), .A3(new_n1024), .A4(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1042), .A2(new_n1126), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1124), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1034), .A2(new_n1036), .A3(new_n785), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1035), .B1(new_n1131), .B2(new_n1032), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1024), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1132), .B1(new_n1133), .B2(new_n1041), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1130), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1119), .A2(new_n1120), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1117), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1130), .A2(new_n1134), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT124), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1044), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(G290), .A2(G1986), .ZN(new_n1141));
  OR3_X1    g716(.A1(new_n1141), .A2(new_n933), .A3(KEYINPUT104), .ZN(new_n1142));
  NAND3_X1  g717(.A1(G290), .A2(KEYINPUT104), .A3(G1986), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1142), .A2(new_n921), .A3(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT105), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n926), .A2(new_n1145), .A3(new_n931), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n947), .B1(new_n1140), .B2(new_n1146), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g722(.A(G227), .ZN(new_n1149));
  AND3_X1   g723(.A1(new_n864), .A2(new_n648), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g724(.A(G229), .ZN(new_n1151));
  NAND4_X1  g725(.A1(new_n1150), .A2(new_n914), .A3(G319), .A4(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g726(.A(new_n1152), .B(KEYINPUT127), .ZN(G308));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n1154));
  XNOR2_X1  g728(.A(new_n1152), .B(new_n1154), .ZN(G225));
endmodule


