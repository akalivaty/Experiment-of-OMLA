//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 1 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G116), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G119), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT68), .B(G116), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  OAI211_X1 g006(.A(KEYINPUT5), .B(new_n190), .C1(new_n191), .C2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT85), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n188), .A2(KEYINPUT68), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT68), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G116), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G119), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT85), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n199), .A2(new_n200), .A3(KEYINPUT5), .A4(new_n190), .ZN(new_n201));
  INV_X1    g015(.A(G113), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT5), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n202), .B1(new_n189), .B2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n194), .A2(new_n201), .A3(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n192), .B1(new_n195), .B2(new_n197), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT2), .B(G113), .ZN(new_n207));
  OR3_X1    g021(.A1(new_n206), .A2(new_n207), .A3(new_n189), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  OR2_X1    g023(.A1(KEYINPUT77), .A2(G104), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT77), .A2(G104), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n213), .A3(G104), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT3), .A2(G107), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NOR3_X1   g031(.A1(new_n214), .A2(new_n217), .A3(G101), .ZN(new_n218));
  INV_X1    g032(.A(G101), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n210), .A2(new_n213), .A3(new_n211), .ZN(new_n220));
  INV_X1    g034(.A(G104), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G107), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n219), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n209), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G110), .B(G122), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n226), .B(KEYINPUT8), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n193), .A2(new_n204), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n208), .A2(new_n228), .ZN(new_n229));
  OR2_X1    g043(.A1(new_n229), .A2(new_n224), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n225), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT86), .ZN(new_n232));
  OAI21_X1  g046(.A(G101), .B1(new_n214), .B2(new_n217), .ZN(new_n233));
  AND2_X1   g047(.A1(KEYINPUT77), .A2(G104), .ZN(new_n234));
  NOR2_X1   g048(.A1(KEYINPUT77), .A2(G104), .ZN(new_n235));
  OAI22_X1  g049(.A1(new_n234), .A2(new_n235), .B1(KEYINPUT3), .B2(G107), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n236), .A2(new_n219), .A3(new_n215), .A4(new_n216), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n233), .A2(new_n237), .A3(KEYINPUT4), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT78), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n233), .A2(new_n237), .A3(KEYINPUT78), .A4(KEYINPUT4), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n243), .B(G101), .C1(new_n214), .C2(new_n217), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n190), .B1(new_n191), .B2(new_n192), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n207), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n247), .B(new_n207), .C1(new_n206), .C2(new_n189), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n245), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n242), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT80), .B1(new_n218), .B2(new_n223), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n220), .A2(new_n222), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G101), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT80), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(new_n256), .A3(new_n237), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(new_n208), .A3(new_n228), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n252), .A2(new_n226), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G146), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(G143), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT64), .B(G143), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n262), .B1(new_n263), .B2(new_n261), .ZN(new_n264));
  INV_X1    g078(.A(G128), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n261), .A2(G143), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(KEYINPUT1), .ZN(new_n267));
  OR2_X1    g081(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n266), .ZN(new_n269));
  INV_X1    g083(.A(G143), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT64), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT64), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G143), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n269), .B1(new_n274), .B2(G146), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT1), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n276), .A3(G128), .ZN(new_n277));
  AOI21_X1  g091(.A(G125), .B1(new_n268), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  AND2_X1   g093(.A1(KEYINPUT0), .A2(G128), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n266), .B(new_n280), .C1(new_n263), .C2(new_n261), .ZN(new_n281));
  NOR2_X1   g095(.A1(KEYINPUT0), .A2(G128), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n281), .B1(new_n264), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G125), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G953), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G224), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT7), .ZN(new_n291));
  OR2_X1    g105(.A1(new_n291), .A2(KEYINPUT87), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(KEYINPUT87), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n279), .A2(new_n288), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  OAI211_X1 g108(.A(KEYINPUT87), .B(new_n291), .C1(new_n278), .C2(new_n287), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT86), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n225), .A2(new_n230), .A3(new_n297), .A4(new_n227), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n232), .A2(new_n260), .A3(new_n296), .A4(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G902), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT88), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n299), .A2(KEYINPUT88), .A3(new_n300), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G210), .B1(G237), .B2(G902), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n279), .A2(new_n288), .ZN(new_n307));
  XOR2_X1   g121(.A(new_n290), .B(KEYINPUT84), .Z(new_n308));
  XNOR2_X1  g122(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n250), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n244), .B1(new_n311), .B2(new_n248), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(new_n240), .B2(new_n241), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n229), .B1(new_n253), .B2(new_n257), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT83), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n226), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT83), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n252), .A2(new_n317), .A3(new_n259), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT6), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n320), .B1(new_n319), .B2(new_n260), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n310), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n305), .A2(new_n306), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n306), .B1(new_n305), .B2(new_n324), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n187), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT89), .ZN(new_n328));
  INV_X1    g142(.A(new_n187), .ZN(new_n329));
  INV_X1    g143(.A(new_n306), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n299), .A2(KEYINPUT88), .A3(new_n300), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT88), .B1(new_n299), .B2(new_n300), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n319), .A2(new_n260), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT6), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n309), .B1(new_n335), .B2(new_n321), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n330), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n305), .A2(new_n306), .A3(new_n324), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n329), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT89), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n328), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G217), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n343), .B1(G234), .B2(new_n300), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT72), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(new_n192), .B2(G128), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n192), .A2(G128), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n265), .A2(KEYINPUT23), .A3(G119), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(G119), .B(G128), .ZN(new_n351));
  AND2_X1   g165(.A1(KEYINPUT24), .A2(G110), .ZN(new_n352));
  NOR2_X1   g166(.A1(KEYINPUT24), .A2(G110), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n350), .A2(G110), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  AND2_X1   g169(.A1(G125), .A2(G140), .ZN(new_n356));
  NOR2_X1   g170(.A1(G125), .A2(G140), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT16), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OR3_X1    g172(.A1(new_n286), .A2(KEYINPUT16), .A3(G140), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n358), .A2(G146), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(G146), .B1(new_n358), .B2(new_n359), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n355), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n265), .A2(G119), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n192), .A2(G128), .ZN(new_n364));
  OAI22_X1  g178(.A1(new_n363), .A2(new_n364), .B1(new_n353), .B2(new_n352), .ZN(new_n365));
  INV_X1    g179(.A(G110), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n347), .A2(new_n349), .A3(new_n366), .A4(new_n348), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n358), .A2(new_n359), .A3(G146), .ZN(new_n369));
  OR2_X1    g183(.A1(new_n356), .A2(new_n357), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n261), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n362), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT71), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT71), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n362), .A2(new_n375), .A3(new_n372), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT22), .B(G137), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n289), .A2(G221), .A3(G234), .ZN(new_n379));
  XOR2_X1   g193(.A(new_n378), .B(new_n379), .Z(new_n380));
  AOI21_X1  g194(.A(new_n345), .B1(new_n377), .B2(new_n380), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n362), .A2(new_n375), .A3(new_n372), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n375), .B1(new_n362), .B2(new_n372), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n345), .B(new_n380), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT73), .ZN(new_n387));
  OR2_X1    g201(.A1(new_n373), .A2(new_n380), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n386), .A2(new_n387), .A3(new_n300), .A4(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n380), .B1(new_n382), .B2(new_n383), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT72), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n391), .A2(new_n300), .A3(new_n388), .A4(new_n384), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT73), .ZN(new_n393));
  XOR2_X1   g207(.A(KEYINPUT74), .B(KEYINPUT25), .Z(new_n394));
  AND3_X1   g208(.A1(new_n389), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n391), .A2(new_n388), .A3(new_n384), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n396), .A2(KEYINPUT75), .A3(KEYINPUT25), .A4(new_n300), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT75), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT25), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n398), .B1(new_n392), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n344), .B1(new_n395), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n344), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n396), .A2(new_n300), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n271), .A2(new_n273), .A3(new_n261), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(G143), .B2(new_n261), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n407), .A2(new_n283), .B1(new_n275), .B2(new_n280), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT65), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT11), .ZN(new_n410));
  INV_X1    g224(.A(G134), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n410), .B1(new_n411), .B2(G137), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(G137), .ZN(new_n413));
  INV_X1    g227(.A(G137), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(KEYINPUT11), .A3(G134), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(G131), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n408), .A2(new_n409), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G131), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n416), .B(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT65), .B1(new_n420), .B2(new_n285), .ZN(new_n421));
  INV_X1    g235(.A(new_n416), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n414), .A2(G134), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n413), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G131), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n422), .A2(new_n419), .B1(new_n425), .B2(KEYINPUT66), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n425), .A2(KEYINPUT66), .ZN(new_n427));
  OAI211_X1 g241(.A(G128), .B(new_n266), .C1(new_n263), .C2(new_n261), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n428), .A2(KEYINPUT1), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n264), .A2(new_n267), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n426), .B(new_n427), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n418), .A2(new_n421), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT30), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n249), .A2(new_n250), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n408), .A2(new_n417), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n431), .A2(new_n436), .A3(KEYINPUT30), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n431), .A2(new_n436), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(new_n435), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G237), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(new_n289), .A3(G210), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(new_n219), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n445));
  XOR2_X1   g259(.A(new_n444), .B(new_n445), .Z(new_n446));
  NAND4_X1  g260(.A1(new_n438), .A2(KEYINPUT69), .A3(new_n441), .A4(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT31), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n447), .A2(new_n448), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT28), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n440), .B(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n432), .A2(new_n435), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI22_X1  g268(.A1(new_n449), .A2(new_n450), .B1(new_n454), .B2(new_n446), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT32), .ZN(new_n456));
  NOR2_X1   g270(.A1(G472), .A2(G902), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n446), .B1(new_n452), .B2(new_n453), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n431), .A2(new_n436), .A3(KEYINPUT30), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n460), .B1(new_n433), .B2(new_n432), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n440), .B1(new_n461), .B2(new_n435), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n462), .A2(KEYINPUT69), .A3(KEYINPUT31), .A4(new_n446), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n447), .A2(new_n448), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n459), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n457), .ZN(new_n466));
  OAI21_X1  g280(.A(KEYINPUT32), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n458), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT70), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n469), .B1(new_n462), .B2(new_n446), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT29), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n438), .A2(new_n441), .ZN(new_n472));
  INV_X1    g286(.A(new_n446), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(KEYINPUT70), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n452), .A2(new_n453), .A3(new_n446), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n470), .A2(new_n471), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n439), .A2(new_n435), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n452), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n473), .A2(new_n471), .ZN(new_n479));
  AOI21_X1  g293(.A(G902), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G472), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n405), .B1(new_n468), .B2(new_n482), .ZN(new_n483));
  XOR2_X1   g297(.A(KEYINPUT81), .B(G469), .Z(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n268), .A2(new_n277), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n486), .A2(new_n224), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n265), .B1(new_n406), .B2(KEYINPUT1), .ZN(new_n488));
  OAI22_X1  g302(.A1(new_n488), .A2(new_n275), .B1(new_n428), .B2(KEYINPUT1), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n224), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT79), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n489), .A2(new_n224), .A3(KEYINPUT79), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n487), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT12), .B1(new_n494), .B2(new_n420), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT10), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n489), .A2(new_n224), .A3(KEYINPUT79), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT79), .B1(new_n489), .B2(new_n224), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n242), .A2(new_n408), .A3(new_n244), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n253), .A2(new_n257), .B1(new_n268), .B2(new_n277), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT10), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n499), .A2(new_n420), .A3(new_n500), .A4(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT12), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n497), .A2(new_n498), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n504), .B(new_n417), .C1(new_n505), .C2(new_n487), .ZN(new_n506));
  XNOR2_X1  g320(.A(G110), .B(G140), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n289), .A2(G227), .ZN(new_n508));
  XOR2_X1   g322(.A(new_n507), .B(new_n508), .Z(new_n509));
  AND4_X1   g323(.A1(new_n495), .A2(new_n503), .A3(new_n506), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n500), .A2(new_n502), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT10), .B1(new_n492), .B2(new_n493), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n417), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n509), .B1(new_n513), .B2(new_n503), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n300), .B(new_n485), .C1(new_n510), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT82), .ZN(new_n516));
  INV_X1    g330(.A(new_n509), .ZN(new_n517));
  INV_X1    g331(.A(new_n503), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n285), .B1(new_n240), .B2(new_n241), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n519), .A2(new_n244), .B1(new_n501), .B2(KEYINPUT10), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n420), .B1(new_n520), .B2(new_n499), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n517), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n495), .A2(new_n503), .A3(new_n506), .A4(new_n509), .ZN(new_n523));
  AOI21_X1  g337(.A(G902), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT82), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n485), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n495), .A2(new_n503), .A3(new_n506), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n517), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n513), .A2(new_n503), .A3(new_n509), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n300), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n516), .A2(new_n526), .B1(G469), .B2(new_n531), .ZN(new_n532));
  XOR2_X1   g346(.A(KEYINPUT9), .B(G234), .Z(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(KEYINPUT76), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n300), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(G221), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT20), .ZN(new_n539));
  XNOR2_X1  g353(.A(G113), .B(G122), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(new_n221), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n442), .A2(new_n289), .A3(G214), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n263), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(G143), .B2(new_n543), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(G131), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n370), .B(KEYINPUT19), .ZN(new_n547));
  AOI211_X1 g361(.A(new_n360), .B(new_n546), .C1(new_n261), .C2(new_n547), .ZN(new_n548));
  OR2_X1    g362(.A1(new_n545), .A2(new_n419), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT18), .ZN(new_n550));
  OR2_X1    g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n545), .B1(new_n550), .B2(new_n419), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n370), .B(new_n261), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n542), .B1(new_n548), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n360), .A2(new_n361), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT17), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n556), .B1(new_n549), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT90), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n546), .A2(new_n557), .ZN(new_n561));
  OAI211_X1 g375(.A(KEYINPUT90), .B(new_n556), .C1(new_n549), .C2(new_n557), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n541), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(G475), .B1(new_n555), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n539), .B1(new_n566), .B2(new_n300), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n539), .A3(new_n300), .ZN(new_n569));
  INV_X1    g383(.A(new_n565), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n541), .B1(new_n563), .B2(new_n564), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n300), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT91), .B(G475), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n568), .A2(new_n569), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n289), .A2(G952), .ZN(new_n575));
  NAND2_X1  g389(.A1(G234), .A2(G237), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  XOR2_X1   g392(.A(KEYINPUT21), .B(G898), .Z(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n576), .A2(G902), .A3(G953), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n578), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(G122), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(G116), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n586), .B1(new_n191), .B2(new_n585), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G107), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT13), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n274), .A2(new_n589), .A3(G128), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n265), .A2(G143), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n591), .B1(new_n263), .B2(new_n265), .ZN(new_n592));
  OAI211_X1 g406(.A(G134), .B(new_n590), .C1(new_n592), .C2(new_n589), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n588), .B(new_n593), .C1(G134), .C2(new_n592), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n592), .B(G134), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n198), .A2(KEYINPUT14), .A3(G122), .ZN(new_n596));
  OAI211_X1 g410(.A(G107), .B(new_n596), .C1(new_n587), .C2(KEYINPUT14), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n595), .B(new_n597), .C1(G107), .C2(new_n587), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n534), .A2(G217), .A3(new_n289), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n594), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n600), .B1(new_n594), .B2(new_n598), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(G902), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT15), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(G478), .ZN(new_n606));
  OR2_X1    g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n604), .A2(new_n606), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n574), .A2(new_n584), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n342), .A2(new_n483), .A3(new_n538), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  OAI21_X1  g426(.A(G472), .B1(new_n465), .B2(G902), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n455), .A2(new_n457), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n613), .A2(new_n402), .A3(new_n614), .A4(new_n404), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n615), .A2(new_n537), .A3(new_n532), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n572), .A2(new_n573), .ZN(new_n617));
  INV_X1    g431(.A(new_n569), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n617), .B1(new_n618), .B2(new_n567), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n604), .A2(G478), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT92), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n603), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g438(.A1(KEYINPUT92), .A2(KEYINPUT33), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n624), .B(new_n625), .C1(new_n601), .C2(new_n602), .ZN(new_n626));
  AOI21_X1  g440(.A(G902), .B1(new_n623), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n620), .B1(new_n627), .B2(G478), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n619), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n327), .A2(new_n583), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n616), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT34), .B(G104), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  NAND2_X1  g449(.A1(new_n607), .A2(new_n608), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n636), .B(new_n617), .C1(new_n618), .C2(new_n567), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n616), .A2(new_n632), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT35), .B(G107), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G9));
  NAND2_X1  g455(.A1(new_n337), .A2(new_n338), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n340), .B1(new_n642), .B2(new_n187), .ZN(new_n643));
  AOI211_X1 g457(.A(KEYINPUT89), .B(new_n329), .C1(new_n337), .C2(new_n338), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n538), .B(new_n610), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT94), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT93), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n380), .A2(KEYINPUT36), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n377), .B(new_n648), .Z(new_n649));
  NOR3_X1   g463(.A1(new_n649), .A2(G902), .A3(new_n344), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n389), .A2(new_n393), .A3(new_n394), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n651), .A2(new_n400), .A3(new_n397), .ZN(new_n652));
  AOI211_X1 g466(.A(new_n647), .B(new_n650), .C1(new_n652), .C2(new_n344), .ZN(new_n653));
  INV_X1    g467(.A(new_n650), .ZN(new_n654));
  AOI21_X1  g468(.A(KEYINPUT93), .B1(new_n402), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n646), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n401), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n403), .B1(new_n657), .B2(new_n651), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n647), .B1(new_n658), .B2(new_n650), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n402), .A2(KEYINPUT93), .A3(new_n654), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(KEYINPUT94), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n613), .A2(new_n614), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n645), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT37), .B(G110), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G12));
  AND2_X1   g480(.A1(new_n656), .A2(new_n661), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n581), .A2(G900), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n577), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n637), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n456), .B1(new_n455), .B2(new_n457), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n465), .A2(KEYINPUT32), .A3(new_n466), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n482), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n538), .A2(new_n674), .A3(new_n339), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n667), .A2(new_n671), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  XNOR2_X1  g491(.A(new_n642), .B(KEYINPUT38), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n653), .A2(new_n655), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n678), .A2(new_n680), .A3(new_n187), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n462), .A2(new_n473), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n441), .A2(new_n473), .A3(new_n477), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n300), .ZN(new_n684));
  OAI21_X1  g498(.A(G472), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n468), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n619), .A3(new_n636), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n688), .A2(KEYINPUT95), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(KEYINPUT95), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n516), .A2(new_n526), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n531), .A2(G469), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n536), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n669), .B(KEYINPUT39), .Z(new_n695));
  OR2_X1    g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT96), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT40), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n696), .B(KEYINPUT96), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT40), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n689), .A2(new_n690), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n274), .ZN(G45));
  NOR2_X1   g518(.A1(new_n630), .A2(new_n670), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n675), .A2(new_n656), .A3(new_n661), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT97), .B(G146), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G48));
  INV_X1    g522(.A(new_n524), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT98), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n709), .A2(new_n710), .A3(G469), .ZN(new_n711));
  INV_X1    g525(.A(G469), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT98), .B1(new_n524), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n691), .A3(new_n536), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n716), .A2(new_n632), .A3(new_n483), .A4(new_n631), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  NAND4_X1  g533(.A1(new_n716), .A2(new_n632), .A3(new_n483), .A4(new_n638), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  AOI21_X1  g535(.A(new_n609), .B1(new_n468), .B2(new_n482), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n715), .A2(new_n327), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n722), .A2(new_n723), .A3(new_n656), .A4(new_n661), .ZN(new_n724));
  XOR2_X1   g538(.A(KEYINPUT99), .B(G119), .Z(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G21));
  NAND2_X1  g540(.A1(new_n619), .A2(new_n636), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n715), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n405), .ZN(new_n729));
  OR2_X1    g543(.A1(new_n478), .A2(new_n446), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n463), .A2(new_n464), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n466), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT100), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n613), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g548(.A(KEYINPUT100), .B(G472), .C1(new_n465), .C2(G902), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n732), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n728), .A2(new_n632), .A3(new_n729), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NAND4_X1  g552(.A1(new_n723), .A2(new_n679), .A3(new_n705), .A4(new_n736), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G125), .ZN(G27));
  NOR2_X1   g554(.A1(new_n325), .A2(new_n326), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n537), .A2(new_n329), .ZN(new_n742));
  INV_X1    g556(.A(new_n691), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT101), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n528), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n527), .A2(KEYINPUT101), .A3(new_n517), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n529), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n712), .B1(new_n747), .B2(new_n300), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n741), .B(new_n742), .C1(new_n743), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n674), .A2(new_n729), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(KEYINPUT42), .B1(new_n751), .B2(new_n705), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n747), .A2(new_n300), .ZN(new_n753));
  AOI22_X1  g567(.A1(new_n753), .A2(G469), .B1(new_n516), .B2(new_n526), .ZN(new_n754));
  INV_X1    g568(.A(new_n742), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n754), .A2(new_n642), .A3(new_n755), .ZN(new_n756));
  AND4_X1   g570(.A1(KEYINPUT42), .A2(new_n756), .A3(new_n483), .A4(new_n705), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n752), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g572(.A(KEYINPUT102), .B(G131), .Z(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(G33));
  INV_X1    g574(.A(KEYINPUT103), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n574), .A2(new_n761), .A3(new_n636), .A4(new_n669), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT103), .B1(new_n637), .B2(new_n670), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n756), .A2(new_n483), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G134), .ZN(G36));
  NOR2_X1   g580(.A1(new_n642), .A2(new_n329), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(KEYINPUT104), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT43), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n769), .B1(new_n574), .B2(new_n629), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n619), .A2(KEYINPUT43), .A3(new_n628), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n663), .A3(new_n679), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT44), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n768), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT105), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n773), .A2(new_n774), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n768), .B(KEYINPUT105), .C1(new_n773), .C2(new_n774), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n780), .A2(KEYINPUT106), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n530), .A2(new_n782), .ZN(new_n783));
  OAI211_X1 g597(.A(G469), .B(new_n783), .C1(new_n747), .C2(new_n782), .ZN(new_n784));
  NAND2_X1  g598(.A1(G469), .A2(G902), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT46), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n743), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n785), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n536), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n695), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n780), .A2(KEYINPUT106), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n781), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  INV_X1    g608(.A(KEYINPUT47), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n790), .B(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n674), .A2(new_n729), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n796), .A2(new_n705), .A3(new_n767), .A4(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  NOR4_X1   g613(.A1(new_n678), .A2(new_n405), .A3(new_n686), .A4(new_n755), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n714), .A2(new_n691), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT49), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n800), .A2(new_n574), .A3(new_n629), .A4(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT108), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n636), .A2(KEYINPUT107), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n636), .A2(KEYINPUT107), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n574), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n619), .A2(new_n628), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n342), .A2(new_n584), .A3(new_n616), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n611), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n804), .B1(new_n811), .B2(new_n664), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n694), .B1(new_n328), .B2(new_n341), .ZN(new_n813));
  INV_X1    g627(.A(new_n663), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n667), .A2(new_n813), .A3(new_n610), .A4(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(KEYINPUT108), .A3(new_n611), .A4(new_n810), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n724), .A2(new_n737), .A3(new_n717), .A4(new_n720), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n756), .A2(new_n679), .A3(new_n705), .A4(new_n736), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n807), .A2(new_n642), .A3(new_n329), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n674), .A3(new_n538), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n656), .A2(new_n661), .A3(new_n669), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n819), .B(new_n765), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n758), .A2(new_n818), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n817), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT109), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT109), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n817), .A2(new_n824), .A3(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n667), .B(new_n675), .C1(new_n671), .C2(new_n705), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n339), .A2(new_n619), .A3(new_n636), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n670), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n754), .A2(new_n658), .A3(new_n650), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(new_n536), .A3(new_n686), .A4(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n829), .A2(KEYINPUT52), .A3(new_n739), .A4(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n676), .A2(new_n706), .A3(new_n833), .A4(new_n739), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n826), .A2(new_n828), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n837), .A2(KEYINPUT110), .A3(new_n834), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n834), .A2(KEYINPUT110), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n817), .A2(new_n824), .A3(KEYINPUT53), .ZN(new_n842));
  OAI22_X1  g656(.A1(new_n838), .A2(KEYINPUT53), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(KEYINPUT54), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n838), .A2(KEYINPUT111), .A3(KEYINPUT53), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT111), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n837), .A2(new_n834), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n817), .A2(new_n824), .A3(new_n827), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n827), .B1(new_n817), .B2(new_n824), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n846), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n841), .B1(new_n826), .B2(new_n828), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n845), .B(new_n852), .C1(KEYINPUT53), .C2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n844), .B1(new_n854), .B2(KEYINPUT54), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n715), .A2(new_n329), .A3(new_n642), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n770), .A2(new_n771), .A3(new_n577), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n856), .A2(new_n857), .A3(new_n483), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT48), .ZN(new_n859));
  INV_X1    g673(.A(new_n686), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n856), .A2(new_n729), .A3(new_n578), .A4(new_n860), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n859), .B(new_n575), .C1(new_n630), .C2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n857), .A2(new_n729), .A3(new_n736), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n678), .A2(new_n187), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(new_n716), .A3(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n866), .A2(KEYINPUT50), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n866), .A2(KEYINPUT50), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n861), .A2(new_n619), .A3(new_n629), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n801), .A2(new_n537), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n768), .B(new_n864), .C1(new_n796), .C2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n856), .A2(new_n857), .A3(new_n679), .A4(new_n736), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT112), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n870), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n863), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI211_X1 g691(.A(new_n862), .B(new_n877), .C1(new_n863), .C2(new_n875), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n864), .A2(new_n723), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n855), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(G952), .A2(G953), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n803), .B1(new_n880), .B2(new_n881), .ZN(G75));
  INV_X1    g696(.A(KEYINPUT56), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n843), .A2(G902), .ZN(new_n884));
  INV_X1    g698(.A(G210), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n335), .A2(new_n309), .A3(new_n321), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n324), .ZN(new_n888));
  XNOR2_X1  g702(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n888), .B(new_n889), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n886), .A2(new_n890), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n289), .A2(G952), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(G51));
  NOR2_X1   g708(.A1(new_n841), .A2(new_n842), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n850), .B2(new_n851), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT54), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n785), .B(KEYINPUT57), .ZN(new_n898));
  OAI22_X1  g712(.A1(new_n897), .A2(new_n898), .B1(new_n514), .B2(new_n510), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n784), .B(KEYINPUT115), .Z(new_n900));
  NAND3_X1  g714(.A1(new_n843), .A2(G902), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n893), .B1(new_n899), .B2(new_n901), .ZN(G54));
  NAND2_X1  g716(.A1(KEYINPUT58), .A2(G475), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n896), .A2(new_n300), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n555), .A2(new_n565), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT116), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT116), .ZN(new_n907));
  INV_X1    g721(.A(new_n905), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n907), .B(new_n908), .C1(new_n884), .C2(new_n903), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n893), .B1(new_n904), .B2(new_n905), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n906), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT117), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT117), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n906), .A2(new_n909), .A3(new_n910), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(G60));
  NAND2_X1  g729(.A1(new_n623), .A2(new_n626), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  XOR2_X1   g731(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n918));
  NAND2_X1  g732(.A1(G478), .A2(G902), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n917), .B1(new_n855), .B2(new_n920), .ZN(new_n921));
  OR3_X1    g735(.A1(new_n897), .A2(new_n917), .A3(new_n920), .ZN(new_n922));
  INV_X1    g736(.A(new_n893), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(G63));
  XNOR2_X1  g738(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT120), .ZN(new_n927));
  NAND2_X1  g741(.A1(G217), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT119), .Z(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT60), .Z(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n927), .B1(new_n896), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n826), .A2(new_n828), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT53), .B1(new_n933), .B2(new_n847), .ZN(new_n934));
  OAI211_X1 g748(.A(KEYINPUT120), .B(new_n930), .C1(new_n934), .C2(new_n895), .ZN(new_n935));
  INV_X1    g749(.A(new_n396), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n932), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n923), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n649), .B1(new_n932), .B2(new_n935), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n926), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n932), .A2(new_n935), .ZN(new_n941));
  INV_X1    g755(.A(new_n649), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n943), .A2(new_n923), .A3(new_n925), .A4(new_n937), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n940), .A2(new_n944), .ZN(G66));
  INV_X1    g759(.A(G224), .ZN(new_n946));
  OAI21_X1  g760(.A(G953), .B1(new_n580), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n817), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n948), .A2(new_n818), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n947), .B1(new_n949), .B2(G953), .ZN(new_n950));
  XNOR2_X1  g764(.A(KEYINPUT122), .B(KEYINPUT123), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n335), .B(new_n321), .C1(G898), .C2(new_n289), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n952), .B(new_n953), .Z(G69));
  NOR2_X1   g768(.A1(new_n750), .A2(new_n830), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n791), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n829), .A2(new_n739), .ZN(new_n957));
  AOI211_X1 g771(.A(new_n758), .B(new_n957), .C1(new_n751), .C2(new_n764), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n793), .A2(new_n798), .A3(new_n956), .A4(new_n958), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n959), .A2(KEYINPUT126), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(KEYINPUT126), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n960), .A2(new_n289), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(G900), .A2(G953), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n461), .B(new_n547), .Z(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  XOR2_X1   g780(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n703), .B2(new_n957), .ZN(new_n968));
  INV_X1    g782(.A(new_n957), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT62), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n970), .A2(KEYINPUT124), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n689), .A2(new_n690), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n699), .A2(new_n702), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n969), .B(new_n972), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n793), .A2(new_n968), .A3(new_n975), .A4(new_n798), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n698), .A2(new_n483), .A3(new_n767), .A4(new_n809), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n289), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n964), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(KEYINPUT125), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT125), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n979), .A2(new_n982), .A3(new_n964), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n966), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n289), .B1(G227), .B2(G900), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n985), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n966), .A2(new_n987), .A3(new_n981), .A4(new_n983), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n986), .A2(new_n988), .ZN(G72));
  NAND3_X1  g803(.A1(new_n960), .A2(new_n949), .A3(new_n961), .ZN(new_n990));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT63), .Z(new_n992));
  AOI211_X1 g806(.A(new_n446), .B(new_n472), .C1(new_n990), .C2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n949), .ZN(new_n994));
  OR3_X1    g808(.A1(new_n976), .A2(new_n994), .A3(new_n978), .ZN(new_n995));
  AOI211_X1 g809(.A(new_n473), .B(new_n462), .C1(new_n995), .C2(new_n992), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n470), .B(new_n474), .C1(new_n473), .C2(new_n472), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n992), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT127), .Z(new_n999));
  AND2_X1   g813(.A1(new_n854), .A2(new_n999), .ZN(new_n1000));
  NOR4_X1   g814(.A1(new_n993), .A2(new_n996), .A3(new_n893), .A4(new_n1000), .ZN(G57));
endmodule


