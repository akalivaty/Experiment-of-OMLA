//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n569, new_n570, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1185, new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT64), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT65), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n454), .A2(new_n448), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G137), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT66), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NOR3_X1   g048(.A1(new_n468), .A2(new_n473), .A3(KEYINPUT68), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n475));
  INV_X1    g050(.A(G137), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n463), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT66), .B(G2105), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n475), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n465), .B1(new_n474), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g058(.A(KEYINPUT67), .B1(new_n466), .B2(new_n467), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n478), .A2(new_n485), .A3(new_n479), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n484), .A2(new_n486), .A3(G125), .ZN(new_n487));
  NAND2_X1  g062(.A1(G113), .A2(G2104), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n481), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n483), .A2(new_n489), .ZN(G160));
  NOR2_X1   g065(.A1(new_n466), .A2(new_n467), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(new_n481), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  OAI221_X1 g068(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n481), .C2(G112), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n491), .A2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G136), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n493), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G162));
  AND2_X1   g073(.A1(G126), .A2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(new_n466), .B2(new_n467), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT69), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G114), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n469), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n500), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AND3_X1   g082(.A1(new_n470), .A2(new_n472), .A3(G138), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n508), .A2(new_n509), .A3(new_n484), .A4(new_n486), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n470), .A2(new_n472), .A3(G138), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT4), .B1(new_n511), .B2(new_n491), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n507), .B1(new_n510), .B2(new_n512), .ZN(G164));
  XNOR2_X1  g088(.A(KEYINPUT5), .B(G543), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT70), .A2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT70), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT71), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n516), .A2(KEYINPUT6), .A3(new_n517), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n524), .A2(KEYINPUT6), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n523), .A2(G543), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n521), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n523), .A2(new_n514), .A3(new_n525), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G88), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n529), .B1(new_n520), .B2(KEYINPUT71), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n527), .A2(new_n530), .ZN(G166));
  NAND3_X1  g106(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n526), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G51), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n528), .A2(G89), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n534), .A2(new_n536), .A3(new_n537), .A4(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(G168));
  NAND2_X1  g116(.A1(new_n535), .A2(G52), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n519), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n528), .A2(G90), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n542), .A2(new_n544), .A3(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  NAND2_X1  g122(.A1(new_n535), .A2(G43), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n519), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n528), .A2(G81), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  NAND3_X1  g133(.A1(new_n535), .A2(KEYINPUT9), .A3(G53), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n526), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n528), .A2(G91), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n514), .A2(G65), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n559), .A2(new_n562), .A3(new_n563), .A4(new_n567), .ZN(G299));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n540), .B(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(G286));
  OR2_X1    g146(.A1(new_n527), .A2(new_n530), .ZN(G303));
  NAND2_X1  g147(.A1(new_n535), .A2(G49), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n528), .A2(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  NAND4_X1  g151(.A1(new_n523), .A2(new_n514), .A3(G86), .A4(new_n525), .ZN(new_n577));
  AND2_X1   g152(.A1(G48), .A2(G543), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n523), .A2(new_n525), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n581));
  AND2_X1   g156(.A1(KEYINPUT5), .A2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(KEYINPUT5), .A2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(G61), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n581), .B1(new_n586), .B2(new_n518), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n580), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n519), .B1(new_n584), .B2(new_n585), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(new_n581), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n590), .ZN(G305));
  NAND2_X1  g166(.A1(new_n528), .A2(G85), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  XNOR2_X1  g168(.A(KEYINPUT75), .B(G47), .ZN(new_n594));
  OAI221_X1 g169(.A(new_n592), .B1(new_n519), .B2(new_n593), .C1(new_n526), .C2(new_n594), .ZN(G290));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NOR2_X1   g171(.A1(G301), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n528), .A2(G92), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT10), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n514), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n524), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(G54), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n526), .B2(KEYINPUT76), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(KEYINPUT76), .B2(new_n526), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n602), .A2(KEYINPUT77), .A3(new_n605), .ZN(new_n609));
  AND2_X1   g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n597), .B1(new_n610), .B2(new_n596), .ZN(G284));
  AOI21_X1  g186(.A(new_n597), .B1(new_n610), .B2(new_n596), .ZN(G321));
  NAND2_X1  g187(.A1(new_n570), .A2(G868), .ZN(new_n613));
  XNOR2_X1  g188(.A(G299), .B(KEYINPUT78), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(G868), .B2(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT79), .ZN(G297));
  XNOR2_X1  g191(.A(new_n615), .B(KEYINPUT80), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n610), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND3_X1  g194(.A1(new_n608), .A2(new_n618), .A3(new_n609), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  OR3_X1    g196(.A1(new_n621), .A2(KEYINPUT81), .A3(new_n596), .ZN(new_n622));
  OAI21_X1  g197(.A(KEYINPUT81), .B1(new_n621), .B2(new_n596), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n622), .B(new_n623), .C1(G868), .C2(new_n553), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g200(.A1(new_n484), .A2(new_n486), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(new_n464), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  INV_X1    g204(.A(G2100), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n492), .A2(G123), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT82), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n636), .B(new_n637), .C1(new_n481), .C2(G111), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n495), .A2(G135), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n633), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT83), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2096), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n631), .A2(new_n632), .A3(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2430), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(KEYINPUT14), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT85), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(new_n645), .B2(new_n646), .ZN(new_n650));
  XOR2_X1   g225(.A(G2451), .B(G2454), .Z(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT86), .Z(new_n660));
  INV_X1    g235(.A(G14), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n656), .B2(new_n658), .ZN(new_n662));
  AND2_X1   g237(.A1(new_n660), .A2(new_n662), .ZN(G401));
  INV_X1    g238(.A(KEYINPUT18), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(KEYINPUT17), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(new_n630), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n667), .B2(KEYINPUT18), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(G2096), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(G227));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n678), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT87), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n680), .A2(new_n681), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT20), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT88), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT89), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n695), .B(new_n696), .Z(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G229));
  XOR2_X1   g273(.A(KEYINPUT90), .B(G29), .Z(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n641), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT31), .B(G11), .Z(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT30), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(G28), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n705), .A2(KEYINPUT96), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n704), .B2(G28), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(KEYINPUT96), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n702), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G1961), .ZN(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n711), .A2(G5), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G301), .B2(G16), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n701), .B(new_n709), .C1(new_n710), .C2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(G21), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G168), .B2(new_n711), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n714), .B1(G1966), .B2(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(G1966), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT97), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n703), .A2(G33), .ZN(new_n722));
  NAND2_X1  g297(.A1(G115), .A2(G2104), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n486), .ZN(new_n724));
  INV_X1    g299(.A(G127), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n481), .B1(new_n726), .B2(KEYINPUT95), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(KEYINPUT95), .B2(new_n726), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n481), .A2(G103), .A3(G2104), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT25), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G139), .B2(new_n495), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n722), .B1(new_n732), .B2(new_n703), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(G2072), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n703), .A2(G32), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT26), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n492), .B2(G129), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n495), .A2(G141), .B1(G105), .B2(new_n464), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n735), .B1(new_n741), .B2(new_n703), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT27), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1996), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n699), .A2(G27), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G164), .B2(new_n699), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2078), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n710), .B2(new_n713), .ZN(new_n748));
  NAND2_X1  g323(.A1(G160), .A2(G29), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT24), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n750), .A2(G34), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(G34), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n699), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G2084), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n734), .A2(new_n744), .A3(new_n748), .A4(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(KEYINPUT98), .B1(new_n721), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G16), .A2(G19), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n553), .B2(G16), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT94), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(G1341), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n711), .A2(G20), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT23), .ZN(new_n763));
  INV_X1    g338(.A(G299), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n711), .ZN(new_n765));
  INV_X1    g340(.A(G1956), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n699), .A2(G26), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT28), .Z(new_n769));
  AOI22_X1  g344(.A1(G128), .A2(new_n492), .B1(new_n495), .B2(G140), .ZN(new_n770));
  OAI221_X1 g345(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n481), .C2(G116), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n769), .B1(new_n772), .B2(G29), .ZN(new_n773));
  INV_X1    g348(.A(G2067), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(G162), .A2(new_n700), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G35), .B2(new_n700), .ZN(new_n777));
  INV_X1    g352(.A(G2090), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n781));
  OR3_X1    g356(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n779), .B2(new_n780), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n775), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n761), .A2(new_n767), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n711), .A2(G4), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n610), .B2(new_n711), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n787), .A2(G1348), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(G1348), .ZN(new_n789));
  NOR3_X1   g364(.A1(new_n785), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n719), .B(KEYINPUT97), .ZN(new_n791));
  INV_X1    g366(.A(new_n756), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT98), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n757), .A2(new_n790), .A3(new_n794), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT93), .B(KEYINPUT36), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n699), .A2(G25), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT91), .Z(new_n798));
  NAND2_X1  g373(.A1(new_n492), .A2(G119), .ZN(new_n799));
  OAI221_X1 g374(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n481), .C2(G107), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n495), .A2(G131), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n798), .B1(new_n802), .B2(new_n700), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT35), .B(G1991), .Z(new_n804));
  XOR2_X1   g379(.A(new_n803), .B(new_n804), .Z(new_n805));
  AND2_X1   g380(.A1(new_n711), .A2(G24), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G290), .B2(G16), .ZN(new_n807));
  INV_X1    g382(.A(G1986), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n805), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(G16), .A2(G22), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G303), .B2(new_n711), .ZN(new_n813));
  INV_X1    g388(.A(G1971), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n711), .A2(G6), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G305), .B2(G16), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT32), .B(G1981), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n813), .A2(new_n814), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n815), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n711), .A2(G23), .ZN(new_n823));
  INV_X1    g398(.A(G288), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n824), .B2(new_n711), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT33), .B(G1976), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n825), .B(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n817), .A2(new_n819), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(KEYINPUT92), .B1(new_n822), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n821), .A2(new_n820), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n828), .A2(new_n829), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT92), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n832), .A2(new_n833), .A3(new_n834), .A4(new_n815), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT34), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n811), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n831), .A2(KEYINPUT34), .A3(new_n835), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n796), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n795), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT36), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(KEYINPUT93), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n838), .A2(new_n843), .A3(new_n839), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n841), .A2(KEYINPUT100), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(KEYINPUT100), .B1(new_n841), .B2(new_n844), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(G311));
  NAND2_X1  g422(.A1(new_n841), .A2(new_n844), .ZN(G150));
  NAND2_X1  g423(.A1(new_n535), .A2(G55), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n528), .A2(G93), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n849), .B(new_n850), .C1(new_n519), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(G860), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT37), .Z(new_n854));
  INV_X1    g429(.A(KEYINPUT102), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n610), .A2(G559), .ZN(new_n856));
  XNOR2_X1  g431(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n852), .B(new_n552), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n860), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n855), .B1(new_n863), .B2(KEYINPUT39), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n865));
  AOI211_X1 g440(.A(KEYINPUT102), .B(new_n865), .C1(new_n861), .C2(new_n862), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(G860), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(new_n863), .B2(KEYINPUT39), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n854), .B1(new_n867), .B2(new_n869), .ZN(G145));
  XNOR2_X1  g445(.A(G164), .B(KEYINPUT103), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n732), .B(new_n871), .ZN(new_n872));
  AOI22_X1  g447(.A1(G130), .A2(new_n492), .B1(new_n495), .B2(G142), .ZN(new_n873));
  OAI221_X1 g448(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n481), .C2(G118), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n628), .B(new_n875), .Z(new_n876));
  XNOR2_X1  g451(.A(new_n872), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n772), .B(new_n740), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n802), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n877), .A2(new_n879), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n641), .B(G162), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(G160), .Z(new_n883));
  OR3_X1    g458(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n883), .B1(new_n880), .B2(new_n881), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g463(.A(new_n620), .B(new_n860), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT104), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n606), .A2(new_n764), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n602), .A2(G299), .A3(new_n605), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n892), .A2(new_n890), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT41), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n891), .A2(new_n892), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n896), .A2(KEYINPUT41), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n889), .A2(new_n895), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n889), .A2(new_n895), .A3(new_n897), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n893), .A2(new_n894), .ZN(new_n901));
  OAI21_X1  g476(.A(KEYINPUT105), .B1(new_n889), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n899), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT42), .ZN(new_n904));
  XNOR2_X1  g479(.A(G303), .B(G305), .ZN(new_n905));
  XNOR2_X1  g480(.A(G290), .B(G288), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n905), .B(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT42), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n909), .B(new_n899), .C1(new_n900), .C2(new_n902), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n904), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n908), .B1(new_n904), .B2(new_n910), .ZN(new_n912));
  OAI21_X1  g487(.A(G868), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n852), .A2(new_n596), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(G295));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n914), .ZN(G331));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n907), .B(KEYINPUT107), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n570), .A2(G171), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n540), .A2(G301), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n860), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n919), .A2(new_n920), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n859), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n925), .A2(new_n895), .A3(new_n897), .ZN(new_n926));
  INV_X1    g501(.A(new_n901), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n922), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n921), .A2(KEYINPUT106), .A3(new_n860), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n927), .A2(new_n929), .A3(new_n924), .A4(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n918), .B1(new_n926), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n907), .A3(new_n926), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n885), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n917), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n927), .A2(new_n924), .A3(new_n922), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n929), .A2(new_n924), .A3(new_n930), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n896), .A2(KEYINPUT41), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(new_n927), .B2(KEYINPUT41), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n936), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n918), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n942), .A2(new_n885), .A3(new_n933), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n935), .B1(new_n943), .B2(new_n917), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT44), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n942), .A2(new_n917), .A3(new_n885), .A4(new_n933), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT43), .B1(new_n932), .B2(new_n934), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n945), .A2(new_n950), .ZN(G397));
  INV_X1    g526(.A(new_n489), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT68), .B1(new_n468), .B2(new_n473), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n480), .A2(new_n475), .A3(new_n481), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n952), .A2(G40), .A3(new_n465), .A4(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(G164), .B2(G1384), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(G1996), .A3(new_n740), .ZN(new_n960));
  OR2_X1    g535(.A1(new_n960), .A2(KEYINPUT108), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(KEYINPUT108), .ZN(new_n962));
  INV_X1    g537(.A(G1996), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n961), .A2(new_n962), .B1(new_n741), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n772), .A2(G2067), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n770), .A2(new_n774), .A3(new_n771), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n959), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT109), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n966), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n802), .B(new_n804), .Z(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n959), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  OR2_X1    g551(.A1(new_n976), .A2(KEYINPUT127), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(KEYINPUT127), .ZN(new_n978));
  NOR2_X1   g553(.A1(G290), .A2(G1986), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n959), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT48), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n977), .A2(new_n978), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n959), .B1(new_n969), .B2(new_n740), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n965), .A2(KEYINPUT46), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n984), .A2(KEYINPUT126), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(KEYINPUT126), .ZN(new_n986));
  OAI221_X1 g561(.A(new_n983), .B1(KEYINPUT46), .B2(new_n965), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT47), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n799), .A2(new_n800), .A3(new_n801), .A4(new_n804), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n968), .B1(new_n972), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n959), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n982), .A2(new_n988), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G40), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n483), .A2(new_n993), .A3(new_n489), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n994), .A2(new_n995), .A3(KEYINPUT117), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n997));
  INV_X1    g572(.A(G1384), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n511), .A2(KEYINPUT4), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n478), .A2(new_n479), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n1000), .A2(new_n481), .A3(G138), .ZN(new_n1001));
  AOI22_X1  g576(.A1(new_n626), .A2(new_n999), .B1(new_n1001), .B2(KEYINPUT4), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n997), .B(new_n998), .C1(new_n1002), .C2(new_n507), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n996), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT117), .B1(new_n994), .B2(new_n995), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n766), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1007));
  NOR2_X1   g582(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1008), .B(KEYINPUT120), .ZN(new_n1009));
  NAND3_X1  g584(.A1(G299), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1009), .B1(G299), .B2(new_n1007), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(KEYINPUT45), .B(new_n998), .C1(new_n1002), .C2(new_n507), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n994), .A2(new_n958), .A3(new_n1015), .ZN(new_n1016));
  XOR2_X1   g591(.A(KEYINPUT56), .B(G2072), .Z(new_n1017));
  OR2_X1    g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1006), .A2(new_n1014), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1014), .B1(new_n1006), .B2(new_n1018), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n994), .A2(new_n995), .A3(new_n1003), .ZN(new_n1021));
  INV_X1    g596(.A(G1348), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(G164), .A2(G1384), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n994), .A2(new_n774), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(new_n606), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1019), .B1(new_n1020), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT61), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1006), .A2(new_n1014), .A3(new_n1018), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1030), .B1(new_n1031), .B2(new_n1020), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1006), .A2(new_n1018), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n1013), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1034), .A2(KEYINPUT61), .A3(new_n1019), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n994), .A2(new_n1024), .ZN(new_n1037));
  XOR2_X1   g612(.A(KEYINPUT58), .B(G1341), .Z(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n994), .A2(new_n958), .A3(new_n1015), .A4(new_n963), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1039), .A2(KEYINPUT121), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT121), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n553), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT60), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n606), .B1(new_n1026), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n1047), .B2(new_n1026), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n553), .B(new_n1044), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1027), .A2(KEYINPUT60), .A3(new_n606), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1046), .A2(new_n1049), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1029), .B1(new_n1036), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n540), .A2(G8), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1015), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n502), .A2(new_n504), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G2105), .ZN(new_n1058));
  INV_X1    g633(.A(new_n506), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1058), .A2(new_n1059), .B1(new_n1000), .B2(new_n499), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n481), .A2(new_n509), .A3(G138), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n724), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n509), .B1(new_n508), .B2(new_n1000), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1060), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1064), .A2(KEYINPUT118), .A3(KEYINPUT45), .A4(new_n998), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1056), .A2(new_n994), .A3(new_n958), .A4(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1966), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n994), .A2(new_n995), .A3(new_n1003), .ZN(new_n1068));
  INV_X1    g643(.A(G2084), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1066), .A2(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G8), .ZN(new_n1071));
  OAI211_X1 g646(.A(KEYINPUT51), .B(new_n1054), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1065), .A2(new_n994), .A3(new_n958), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT118), .B1(new_n1024), .B2(KEYINPUT45), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1067), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n994), .A2(new_n995), .A3(new_n1003), .A4(new_n1069), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1073), .B(G8), .C1(new_n1078), .C2(new_n540), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1054), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT123), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT123), .ZN(new_n1082));
  AOI211_X1 g657(.A(new_n1082), .B(new_n1054), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1072), .B(new_n1079), .C1(new_n1081), .C2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(new_n1016), .B2(G2078), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1021), .A2(new_n710), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1085), .A2(G2078), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1086), .B(new_n1087), .C1(new_n1016), .C2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G171), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1086), .B(new_n1087), .C1(new_n1088), .C2(new_n1066), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1090), .B(KEYINPUT54), .C1(G171), .C2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1084), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G1976), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1037), .B(G8), .C1(new_n1094), .C2(G288), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT52), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT52), .B1(G288), .B2(new_n1094), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1096), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n577), .A2(new_n579), .ZN(new_n1100));
  INV_X1    g675(.A(G1981), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n514), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT74), .B1(new_n1102), .B2(new_n519), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n590), .A2(new_n1100), .A3(new_n1101), .A4(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT113), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n588), .A2(KEYINPUT113), .A3(new_n1101), .A4(new_n590), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT115), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT114), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n577), .A2(new_n1110), .A3(new_n579), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1110), .B1(new_n577), .B2(new_n579), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1111), .A2(new_n1112), .A3(new_n589), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1109), .B1(new_n1113), .B2(new_n1101), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n589), .B1(new_n580), .B2(KEYINPUT114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n577), .A2(new_n1110), .A3(new_n579), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1117), .A2(KEYINPUT115), .A3(G1981), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1108), .A2(new_n1114), .A3(KEYINPUT49), .A4(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT116), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1101), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1106), .A2(new_n1107), .B1(new_n1122), .B2(KEYINPUT115), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1123), .A2(KEYINPUT116), .A3(KEYINPUT49), .A4(new_n1114), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1037), .A2(G8), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1123), .A2(new_n1114), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT49), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1099), .B1(new_n1125), .B2(new_n1129), .ZN(new_n1130));
  XOR2_X1   g705(.A(KEYINPUT110), .B(G1971), .Z(new_n1131));
  NAND2_X1  g706(.A1(new_n1016), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT111), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1132), .A2(new_n1133), .B1(new_n1068), .B2(new_n778), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1016), .A2(KEYINPUT111), .A3(new_n1131), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1071), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(G166), .A2(new_n1071), .ZN(new_n1137));
  XNOR2_X1  g712(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1137), .B(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT117), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n997), .B1(new_n1064), .B2(new_n998), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1141), .B1(new_n1142), .B2(new_n956), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1143), .A2(new_n1003), .A3(new_n996), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1132), .B1(new_n1144), .B2(G2090), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(G8), .ZN(new_n1146));
  XOR2_X1   g721(.A(new_n1137), .B(new_n1138), .Z(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1130), .A2(new_n1140), .A3(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1093), .A2(new_n1149), .ZN(new_n1150));
  OR3_X1    g725(.A1(new_n1089), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1151));
  OAI21_X1  g726(.A(KEYINPUT124), .B1(new_n1089), .B2(G171), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1091), .A2(G171), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT54), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1053), .A2(new_n1150), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1125), .A2(new_n1129), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1099), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1159), .A2(new_n1160), .A3(new_n1136), .A4(new_n1139), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1108), .ZN(new_n1162));
  NOR2_X1   g737(.A1(G288), .A2(G1976), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1162), .B1(new_n1159), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1161), .B1(new_n1164), .B2(new_n1126), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1070), .A2(new_n1071), .A3(G286), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1130), .A2(new_n1148), .A3(new_n1140), .A4(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT63), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1166), .A2(KEYINPUT63), .ZN(new_n1170));
  OR2_X1    g745(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1170), .A2(new_n1171), .A3(new_n1130), .A4(new_n1140), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1165), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1157), .A2(new_n1158), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1158), .B1(new_n1157), .B2(new_n1173), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1149), .A2(new_n1153), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1176), .B1(KEYINPUT62), .B2(new_n1084), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1177), .B1(KEYINPUT62), .B2(new_n1084), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n1174), .A2(new_n1175), .A3(new_n1178), .ZN(new_n1179));
  AND2_X1   g754(.A1(G290), .A2(G1986), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n959), .B1(new_n1180), .B2(new_n979), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n973), .A2(new_n1181), .A3(new_n975), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n992), .B1(new_n1179), .B2(new_n1182), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g758(.A1(G227), .A2(new_n461), .ZN(new_n1185));
  NAND2_X1  g759(.A1(new_n697), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g760(.A(new_n1186), .B1(new_n660), .B2(new_n662), .ZN(new_n1187));
  AND3_X1   g761(.A1(new_n1187), .A2(new_n887), .A3(new_n948), .ZN(G308));
  NAND3_X1  g762(.A1(new_n1187), .A2(new_n887), .A3(new_n948), .ZN(G225));
endmodule


