//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942;
  XNOR2_X1  g000(.A(G127gat), .B(G155gat), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206));
  OR2_X1    g005(.A1(new_n206), .A2(G1gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT16), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n208), .B2(G1gat), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT91), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n207), .A2(KEYINPUT91), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(G8gat), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT92), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n211), .A2(KEYINPUT92), .A3(G8gat), .A4(new_n212), .ZN(new_n216));
  INV_X1    g015(.A(G8gat), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n215), .A2(new_n216), .B1(new_n217), .B2(new_n210), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT21), .ZN(new_n219));
  XNOR2_X1  g018(.A(G57gat), .B(G64gat), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g021(.A(G71gat), .B(G78gat), .Z(new_n223));
  OR2_X1    g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n223), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n218), .B1(new_n219), .B2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(G183gat), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(G183gat), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n229), .A2(G231gat), .A3(G233gat), .A4(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n230), .ZN(new_n232));
  INV_X1    g031(.A(G231gat), .ZN(new_n233));
  INV_X1    g032(.A(G233gat), .ZN(new_n234));
  OAI22_X1  g033(.A1(new_n232), .A2(new_n228), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n205), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n226), .A2(new_n219), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n238), .B(new_n239), .Z(new_n240));
  NAND3_X1  g039(.A1(new_n231), .A2(new_n235), .A3(new_n205), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n237), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n240), .ZN(new_n243));
  INV_X1    g042(.A(new_n241), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n243), .B1(new_n244), .B2(new_n236), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(G29gat), .A2(G36gat), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n247), .A2(KEYINPUT14), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(KEYINPUT14), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT87), .B(G29gat), .Z(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(G36gat), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n248), .B(new_n249), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT88), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G43gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(G50gat), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(G50gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(KEYINPUT15), .A3(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n255), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT90), .B(G50gat), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n257), .B1(new_n262), .B2(new_n256), .ZN(new_n263));
  XOR2_X1   g062(.A(KEYINPUT89), .B(KEYINPUT15), .Z(new_n264));
  OR3_X1    g063(.A1(new_n253), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  OR2_X1    g065(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n267));
  NAND2_X1  g066(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n267), .A2(G85gat), .A3(G92gat), .A4(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n270));
  NAND2_X1  g069(.A1(G85gat), .A2(G92gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(G99gat), .A2(G106gat), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n270), .A2(new_n271), .B1(new_n272), .B2(KEYINPUT8), .ZN(new_n273));
  OR2_X1    g072(.A1(G85gat), .A2(G92gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n269), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  OR2_X1    g074(.A1(G99gat), .A2(G106gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n272), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n272), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n269), .A2(new_n273), .A3(new_n278), .A4(new_n274), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT41), .ZN(new_n282));
  NAND2_X1  g081(.A1(G232gat), .A2(G233gat), .ZN(new_n283));
  OAI22_X1  g082(.A1(new_n266), .A2(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n261), .A2(KEYINPUT17), .A3(new_n265), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT17), .B1(new_n261), .B2(new_n265), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n284), .B1(new_n287), .B2(new_n281), .ZN(new_n288));
  XOR2_X1   g087(.A(G190gat), .B(G218gat), .Z(new_n289));
  XNOR2_X1  g088(.A(new_n289), .B(KEYINPUT96), .ZN(new_n290));
  XOR2_X1   g089(.A(new_n288), .B(new_n290), .Z(new_n291));
  XOR2_X1   g090(.A(G134gat), .B(G162gat), .Z(new_n292));
  NAND2_X1  g091(.A1(new_n283), .A2(new_n282), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n291), .B(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G120gat), .B(G148gat), .ZN(new_n296));
  INV_X1    g095(.A(G176gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G204gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n280), .B(new_n226), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT97), .B1(new_n303), .B2(KEYINPUT10), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n280), .A2(KEYINPUT10), .A3(new_n225), .A4(new_n224), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT97), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT10), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n302), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n304), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT98), .ZN(new_n310));
  NAND2_X1  g109(.A1(G230gat), .A2(G233gat), .ZN(new_n311));
  AND3_X1   g110(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n310), .B1(new_n309), .B2(new_n311), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n302), .A2(new_n311), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n301), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  AOI211_X1 g116(.A(new_n315), .B(new_n300), .C1(new_n309), .C2(new_n311), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NOR3_X1   g119(.A1(new_n246), .A2(new_n295), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n218), .B1(new_n285), .B2(new_n286), .ZN(new_n322));
  OR2_X1    g121(.A1(new_n218), .A2(new_n266), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G229gat), .A2(G233gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n325), .B(KEYINPUT93), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT18), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT18), .ZN(new_n328));
  INV_X1    g127(.A(new_n326), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n322), .A2(new_n323), .A3(new_n328), .A4(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT94), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n218), .A2(new_n266), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n218), .A2(new_n266), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XOR2_X1   g134(.A(new_n326), .B(KEYINPUT13), .Z(new_n336));
  OAI21_X1  g135(.A(new_n332), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n336), .ZN(new_n338));
  OAI211_X1 g137(.A(KEYINPUT94), .B(new_n338), .C1(new_n333), .C2(new_n334), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n331), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT11), .B(G169gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(G197gat), .ZN(new_n343));
  XOR2_X1   g142(.A(G113gat), .B(G141gat), .Z(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(KEYINPUT12), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n340), .A3(new_n346), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT72), .ZN(new_n351));
  NAND3_X1  g150(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n352), .B1(G183gat), .B2(G190gat), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT64), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT23), .ZN(new_n356));
  INV_X1    g155(.A(G169gat), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(new_n357), .A3(new_n297), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n358), .A2(new_n359), .B1(G169gat), .B2(G176gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n354), .ZN(new_n361));
  OR2_X1    g160(.A1(G183gat), .A2(G190gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT64), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n361), .A2(new_n362), .A3(new_n363), .A4(new_n352), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n355), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT25), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT65), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT65), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n365), .A2(new_n369), .A3(new_n366), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n361), .A2(KEYINPUT66), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT66), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n354), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n371), .A2(new_n352), .A3(new_n362), .A4(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n374), .A2(KEYINPUT25), .A3(new_n360), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n368), .A2(new_n370), .A3(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT27), .B(G183gat), .ZN(new_n377));
  INV_X1    g176(.A(G190gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  XOR2_X1   g178(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G183gat), .A2(G190gat), .ZN(new_n382));
  OR3_X1    g181(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n383), .B(new_n384), .C1(new_n357), .C2(new_n297), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n381), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n376), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(G113gat), .ZN(new_n388));
  OR3_X1    g187(.A1(new_n388), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT69), .B1(new_n388), .B2(G120gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT70), .B(G113gat), .ZN(new_n391));
  INV_X1    g190(.A(G120gat), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n389), .B(new_n390), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT1), .ZN(new_n394));
  OR2_X1    g193(.A1(G127gat), .A2(G134gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(G127gat), .A2(G134gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n393), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT68), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n395), .A2(KEYINPUT68), .A3(new_n396), .ZN(new_n401));
  XNOR2_X1  g200(.A(G113gat), .B(G120gat), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n400), .B(new_n401), .C1(KEYINPUT1), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n387), .B(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G227gat), .A2(G233gat), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n351), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT34), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT34), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n351), .B(new_n410), .C1(new_n405), .C2(new_n407), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G15gat), .B(G43gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(G71gat), .ZN(new_n414));
  INV_X1    g213(.A(G99gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  OR2_X1    g216(.A1(new_n417), .A2(KEYINPUT71), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(KEYINPUT71), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n418), .A2(KEYINPUT33), .A3(new_n419), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n387), .A2(new_n404), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n387), .A2(new_n404), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(KEYINPUT32), .B(new_n420), .C1(new_n423), .C2(new_n406), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT32), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n405), .A2(new_n407), .B1(new_n425), .B2(KEYINPUT33), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n424), .B1(new_n426), .B2(new_n417), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT33), .ZN(new_n429));
  OAI22_X1  g228(.A1(new_n423), .A2(new_n406), .B1(KEYINPUT32), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n416), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n431), .A2(new_n424), .A3(new_n409), .A4(new_n411), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT36), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n428), .A2(new_n432), .A3(KEYINPUT36), .ZN(new_n436));
  XNOR2_X1  g235(.A(G8gat), .B(G36gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(G92gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT75), .ZN(new_n439));
  INV_X1    g238(.A(G64gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G226gat), .A2(G233gat), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT74), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n365), .A2(new_n369), .A3(new_n366), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n369), .B1(new_n365), .B2(new_n366), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n374), .A2(KEYINPUT25), .A3(new_n360), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n386), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n443), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n376), .A2(KEYINPUT74), .A3(new_n386), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n442), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT73), .ZN(new_n452));
  XNOR2_X1  g251(.A(G197gat), .B(G204gat), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT22), .ZN(new_n454));
  INV_X1    g253(.A(G218gat), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n454), .B1(new_n203), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G211gat), .B(G218gat), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n452), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n457), .A2(new_n459), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n458), .A2(new_n453), .A3(new_n456), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n460), .B1(new_n463), .B2(new_n452), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n442), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n466), .A2(KEYINPUT29), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n387), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NOR3_X1   g268(.A1(new_n451), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n449), .A2(new_n450), .A3(new_n467), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n376), .A2(new_n386), .A3(new_n466), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n464), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n441), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(new_n472), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n465), .ZN(new_n476));
  INV_X1    g275(.A(new_n450), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT74), .B1(new_n376), .B2(new_n386), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n466), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n479), .A2(new_n464), .A3(new_n468), .ZN(new_n480));
  INV_X1    g279(.A(new_n441), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n476), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n474), .A2(new_n482), .A3(KEYINPUT30), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n470), .A2(new_n473), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT30), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n485), .A3(new_n481), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n487));
  NAND2_X1  g286(.A1(G225gat), .A2(G233gat), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT5), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G155gat), .B(G162gat), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G141gat), .B(G148gat), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n492), .B1(KEYINPUT2), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT77), .ZN(new_n495));
  AND2_X1   g294(.A1(KEYINPUT76), .A2(G148gat), .ZN(new_n496));
  NOR2_X1   g295(.A1(KEYINPUT76), .A2(G148gat), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n495), .B(G141gat), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(G141gat), .ZN(new_n499));
  OR2_X1    g298(.A1(KEYINPUT76), .A2(G148gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(KEYINPUT76), .A2(G148gat), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n499), .A2(G148gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT77), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n498), .B(new_n491), .C1(new_n502), .C2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G162gat), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT2), .B1(new_n506), .B2(KEYINPUT78), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n494), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT3), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n496), .A2(new_n497), .ZN(new_n511));
  OAI211_X1 g310(.A(KEYINPUT77), .B(new_n503), .C1(new_n511), .C2(new_n499), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n512), .A2(new_n491), .A3(new_n507), .A4(new_n498), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT3), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n514), .A3(new_n494), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n510), .A2(new_n404), .A3(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n513), .A2(new_n398), .A3(new_n494), .A4(new_n403), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(KEYINPUT4), .A3(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT79), .B(KEYINPUT4), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n490), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n517), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n522), .B1(new_n516), .B2(new_n519), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT4), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n488), .B1(new_n517), .B2(new_n524), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n404), .A2(new_n509), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT80), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(new_n528), .A3(new_n517), .ZN(new_n529));
  INV_X1    g328(.A(new_n488), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n404), .A2(new_n509), .A3(KEYINPUT80), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n532), .A2(KEYINPUT5), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n521), .B1(new_n526), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT0), .B(G57gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(G85gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(G1gat), .B(G29gat), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n536), .B(new_n537), .Z(new_n538));
  AOI21_X1  g337(.A(new_n487), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n521), .ZN(new_n540));
  OAI211_X1 g339(.A(KEYINPUT5), .B(new_n532), .C1(new_n523), .C2(new_n525), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n538), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n542), .A2(new_n543), .A3(new_n487), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n483), .A2(new_n486), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT29), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n465), .B1(new_n548), .B2(new_n515), .ZN(new_n549));
  NAND2_X1  g348(.A1(G228gat), .A2(G233gat), .ZN(new_n550));
  INV_X1    g349(.A(new_n509), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT3), .B1(new_n463), .B2(new_n548), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  OR3_X1    g353(.A1(new_n464), .A2(KEYINPUT82), .A3(KEYINPUT29), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT82), .B1(new_n464), .B2(KEYINPUT29), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(new_n514), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n549), .B1(new_n557), .B2(new_n509), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n554), .B1(new_n558), .B2(new_n550), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT31), .B(G50gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n560), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n562), .B(new_n554), .C1(new_n558), .C2(new_n550), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G78gat), .B(G106gat), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n565), .B(G22gat), .Z(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n561), .A2(new_n566), .A3(new_n563), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n435), .B(new_n436), .C1(new_n547), .C2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n570), .ZN(new_n572));
  AND3_X1   g371(.A1(new_n483), .A2(KEYINPUT83), .A3(new_n486), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT83), .B1(new_n483), .B2(new_n486), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT85), .B1(new_n534), .B2(new_n538), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT85), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n542), .A2(new_n577), .A3(new_n543), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT39), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n530), .B1(new_n529), .B2(new_n531), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT84), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n518), .A2(new_n520), .ZN(new_n584));
  OAI221_X1 g383(.A(new_n583), .B1(new_n582), .B2(new_n581), .C1(new_n488), .C2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n488), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n543), .B1(new_n586), .B2(new_n580), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(KEYINPUT40), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n579), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT40), .B1(new_n585), .B2(new_n587), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n572), .B1(new_n575), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n577), .B1(new_n542), .B2(new_n543), .ZN(new_n593));
  AOI211_X1 g392(.A(KEYINPUT85), .B(new_n538), .C1(new_n540), .C2(new_n541), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n539), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n595), .A2(new_n546), .A3(new_n482), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT37), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n476), .A2(new_n480), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n475), .A2(new_n464), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n479), .A2(new_n465), .A3(new_n468), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n600), .A3(KEYINPUT37), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT38), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n598), .A2(new_n601), .A3(new_n602), .A4(new_n441), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT86), .B1(new_n596), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n546), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n606), .B1(new_n579), .B2(new_n539), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT86), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n607), .A2(new_n608), .A3(new_n482), .A4(new_n603), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n484), .A2(new_n597), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n598), .A2(new_n441), .ZN(new_n611));
  OAI21_X1  g410(.A(KEYINPUT38), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n605), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n571), .B1(new_n592), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT35), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n432), .A2(new_n428), .B1(new_n568), .B2(new_n569), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n615), .B1(new_n616), .B2(new_n547), .ZN(new_n617));
  INV_X1    g416(.A(new_n607), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n615), .B(new_n618), .C1(new_n573), .C2(new_n574), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n617), .B1(new_n620), .B2(new_n616), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n321), .B(new_n350), .C1(new_n614), .C2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n574), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n483), .A2(KEYINPUT83), .A3(new_n486), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n625), .A2(new_n591), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n613), .A2(new_n570), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n571), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n625), .A2(new_n626), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n631), .A2(new_n615), .A3(new_n618), .A4(new_n616), .ZN(new_n632));
  INV_X1    g431(.A(new_n617), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n635), .A2(KEYINPUT99), .A3(new_n321), .A4(new_n350), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n624), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n545), .A2(new_n546), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G1gat), .ZN(G1324gat));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n642), .B1(new_n637), .B2(new_n575), .ZN(new_n643));
  AOI211_X1 g442(.A(KEYINPUT101), .B(new_n631), .C1(new_n624), .C2(new_n636), .ZN(new_n644));
  OR3_X1    g443(.A1(new_n643), .A2(new_n644), .A3(new_n217), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT16), .B(G8gat), .Z(new_n646));
  NAND4_X1  g445(.A1(new_n637), .A2(KEYINPUT42), .A3(new_n575), .A4(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n646), .B1(new_n643), .B2(new_n644), .ZN(new_n648));
  NAND2_X1  g447(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n645), .B(new_n647), .C1(new_n650), .C2(new_n651), .ZN(G1325gat));
  INV_X1    g451(.A(G15gat), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n637), .A2(new_n653), .A3(new_n433), .ZN(new_n654));
  INV_X1    g453(.A(new_n637), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n435), .A2(new_n436), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n656), .B(KEYINPUT102), .Z(new_n657));
  NOR2_X1   g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n654), .B1(new_n658), .B2(new_n653), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT103), .ZN(G1326gat));
  NAND2_X1  g459(.A1(new_n637), .A2(new_n572), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT43), .B(G22gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT104), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n661), .B(new_n663), .ZN(G1327gat));
  NAND2_X1  g463(.A1(new_n242), .A2(new_n245), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(new_n320), .ZN(new_n666));
  AND4_X1   g465(.A1(new_n295), .A2(new_n635), .A3(new_n350), .A4(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n667), .A2(new_n639), .A3(new_n251), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT45), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT45), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n667), .A2(new_n670), .A3(new_n639), .A4(new_n251), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673));
  AOI22_X1  g472(.A1(new_n628), .A2(new_n629), .B1(new_n632), .B2(new_n633), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n291), .B(new_n294), .Z(new_n675));
  OAI21_X1  g474(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n331), .A2(new_n340), .A3(new_n346), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n346), .B1(new_n331), .B2(new_n340), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n348), .A2(KEYINPUT105), .A3(new_n349), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI211_X1 g481(.A(KEYINPUT44), .B(new_n295), .C1(new_n614), .C2(new_n621), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n676), .A2(new_n682), .A3(new_n683), .A4(new_n666), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n250), .B1(new_n684), .B2(new_n638), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n672), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(KEYINPUT106), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n672), .A2(new_n688), .A3(new_n685), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n689), .ZN(G1328gat));
  NAND3_X1  g489(.A1(new_n667), .A2(new_n252), .A3(new_n575), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT107), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n667), .A2(new_n693), .A3(new_n252), .A4(new_n575), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT108), .B1(new_n695), .B2(KEYINPUT46), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(KEYINPUT46), .ZN(new_n697));
  OAI21_X1  g496(.A(G36gat), .B1(new_n684), .B2(new_n631), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n692), .A2(new_n699), .A3(new_n700), .A4(new_n694), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n696), .A2(new_n697), .A3(new_n698), .A4(new_n701), .ZN(G1329gat));
  OR3_X1    g501(.A1(new_n684), .A2(KEYINPUT109), .A3(new_n656), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT109), .B1(new_n684), .B2(new_n656), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(G43gat), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n667), .A2(new_n256), .A3(new_n433), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n705), .A2(KEYINPUT47), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G43gat), .B1(new_n684), .B2(new_n657), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n708), .A2(new_n706), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n707), .B1(KEYINPUT47), .B2(new_n709), .ZN(G1330gat));
  OAI21_X1  g509(.A(new_n262), .B1(new_n684), .B2(new_n570), .ZN(new_n711));
  INV_X1    g510(.A(new_n262), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n667), .A2(new_n712), .A3(new_n572), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT48), .B1(new_n713), .B2(KEYINPUT110), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1331gat));
  NOR2_X1   g515(.A1(new_n682), .A2(new_n319), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n635), .A2(new_n665), .A3(new_n675), .A4(new_n717), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n718), .A2(KEYINPUT111), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(KEYINPUT111), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(new_n638), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT112), .B(G57gat), .Z(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1332gat));
  NOR2_X1   g523(.A1(new_n721), .A2(new_n631), .ZN(new_n725));
  NOR2_X1   g524(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n726));
  AND2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(new_n725), .B2(new_n726), .ZN(G1333gat));
  OAI21_X1  g528(.A(G71gat), .B1(new_n721), .B2(new_n657), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT50), .ZN(new_n731));
  INV_X1    g530(.A(G71gat), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n719), .A2(new_n732), .A3(new_n433), .A4(new_n720), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n731), .B1(new_n730), .B2(new_n733), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(G1334gat));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n570), .ZN(new_n737));
  XNOR2_X1  g536(.A(KEYINPUT113), .B(G78gat), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1335gat));
  NOR2_X1   g538(.A1(new_n682), .A2(new_n665), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n676), .A2(new_n320), .A3(new_n683), .A4(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(G85gat), .B1(new_n741), .B2(new_n638), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n295), .B(new_n740), .C1(new_n614), .C2(new_n621), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(KEYINPUT51), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n319), .A2(G85gat), .A3(new_n638), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT114), .Z(new_n750));
  OAI21_X1  g549(.A(new_n742), .B1(new_n748), .B2(new_n750), .ZN(G1336gat));
  OR2_X1    g550(.A1(new_n741), .A2(new_n631), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G92gat), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n631), .A2(new_n319), .A3(G92gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT115), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(new_n745), .B2(new_n747), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n753), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT117), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n747), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n743), .A2(KEYINPUT117), .A3(new_n759), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  AOI22_X1  g564(.A1(new_n752), .A2(G92gat), .B1(new_n765), .B2(new_n755), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n758), .B1(new_n757), .B2(new_n766), .ZN(G1337gat));
  OAI21_X1  g566(.A(G99gat), .B1(new_n741), .B2(new_n657), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n320), .A2(new_n415), .A3(new_n433), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT118), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n748), .B2(new_n770), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT119), .Z(G1338gat));
  OAI21_X1  g571(.A(G106gat), .B1(new_n741), .B2(new_n570), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT53), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n319), .A2(G106gat), .A3(new_n570), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n773), .B(new_n774), .C1(new_n748), .C2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT120), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n765), .A2(new_n775), .ZN(new_n779));
  AOI211_X1 g578(.A(new_n778), .B(new_n774), .C1(new_n779), .C2(new_n773), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n743), .A2(KEYINPUT117), .A3(new_n759), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT117), .B1(new_n743), .B2(new_n759), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n781), .A2(new_n782), .A3(new_n747), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n773), .B1(new_n783), .B2(new_n776), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT120), .B1(new_n784), .B2(KEYINPUT53), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n777), .B1(new_n780), .B2(new_n785), .ZN(G1339gat));
  AND2_X1   g585(.A1(new_n680), .A2(new_n681), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n321), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n341), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n329), .B1(new_n322), .B2(new_n323), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n790), .A2(KEYINPUT122), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n335), .A2(new_n336), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(KEYINPUT122), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n789), .A2(new_n346), .B1(new_n345), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(new_n312), .B2(new_n313), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n309), .A2(new_n311), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n309), .A2(new_n311), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(KEYINPUT54), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n797), .A2(new_n300), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n318), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n799), .A2(KEYINPUT98), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n301), .B1(new_n806), .B2(new_n796), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n807), .A2(KEYINPUT121), .A3(KEYINPUT55), .A4(new_n800), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n797), .A2(KEYINPUT55), .A3(new_n800), .A4(new_n300), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT121), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n795), .A2(new_n803), .A3(new_n808), .A4(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(new_n675), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n320), .A2(new_n795), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n803), .A2(new_n808), .A3(new_n811), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n787), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n813), .B1(new_n816), .B2(new_n675), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n788), .B1(new_n817), .B2(new_n665), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n575), .A2(new_n638), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n818), .A2(new_n616), .A3(new_n819), .ZN(new_n820));
  OR3_X1    g619(.A1(new_n820), .A2(new_n391), .A3(new_n787), .ZN(new_n821));
  INV_X1    g620(.A(new_n350), .ZN(new_n822));
  INV_X1    g621(.A(new_n820), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT123), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT123), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n820), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n822), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n821), .B1(new_n827), .B2(new_n388), .ZN(G1340gat));
  NAND3_X1  g627(.A1(new_n823), .A2(new_n392), .A3(new_n320), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n319), .B1(new_n824), .B2(new_n826), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(new_n392), .ZN(G1341gat));
  AOI21_X1  g630(.A(G127gat), .B1(new_n823), .B2(new_n665), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n246), .B1(new_n824), .B2(new_n826), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(new_n833), .B2(G127gat), .ZN(G1342gat));
  AND2_X1   g633(.A1(new_n818), .A2(new_n616), .ZN(new_n835));
  INV_X1    g634(.A(G134gat), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(new_n836), .A3(new_n819), .ZN(new_n837));
  OR3_X1    g636(.A1(new_n837), .A2(KEYINPUT56), .A3(new_n675), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT56), .B1(new_n837), .B2(new_n675), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n675), .B1(new_n824), .B2(new_n826), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n838), .B(new_n839), .C1(new_n840), .C2(new_n836), .ZN(G1343gat));
  NAND4_X1  g640(.A1(new_n803), .A2(new_n808), .A3(new_n350), .A4(new_n811), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n295), .B1(new_n842), .B2(new_n814), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n246), .B1(new_n843), .B2(new_n813), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n570), .B1(new_n844), .B2(new_n788), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n819), .A2(new_n656), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n818), .A2(new_n846), .A3(new_n572), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n499), .B1(new_n850), .B2(new_n350), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n818), .A2(new_n572), .A3(new_n657), .A4(new_n819), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(G141gat), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n350), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n847), .A2(new_n682), .A3(new_n849), .A4(new_n848), .ZN(new_n857));
  AOI22_X1  g656(.A1(new_n857), .A2(G141gat), .B1(new_n853), .B2(new_n350), .ZN(new_n858));
  OAI22_X1  g657(.A1(new_n851), .A2(new_n856), .B1(new_n858), .B2(new_n855), .ZN(G1344gat));
  NAND4_X1  g658(.A1(new_n847), .A2(new_n320), .A3(new_n849), .A4(new_n848), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n511), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n803), .A2(new_n808), .A3(new_n811), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n682), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n295), .B1(new_n865), .B2(new_n814), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n246), .B1(new_n866), .B2(new_n813), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n570), .B1(new_n867), .B2(new_n788), .ZN(new_n868));
  INV_X1    g667(.A(new_n511), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n868), .A2(new_n869), .A3(new_n657), .A4(new_n819), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT124), .B1(new_n870), .B2(new_n319), .ZN(new_n871));
  INV_X1    g670(.A(new_n852), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n872), .A2(new_n873), .A3(new_n869), .A4(new_n320), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n321), .A2(new_n787), .ZN(new_n876));
  INV_X1    g675(.A(new_n813), .ZN(new_n877));
  AOI22_X1  g676(.A1(new_n864), .A2(new_n682), .B1(new_n320), .B2(new_n795), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n295), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n876), .B1(new_n879), .B2(new_n246), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT57), .B1(new_n880), .B2(new_n570), .ZN(new_n881));
  INV_X1    g680(.A(new_n844), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n321), .A2(new_n822), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n846), .B(new_n572), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT125), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n848), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n881), .A2(new_n320), .A3(new_n884), .A4(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n848), .A2(new_n885), .ZN(new_n888));
  OAI211_X1 g687(.A(KEYINPUT59), .B(G148gat), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n863), .A2(new_n875), .A3(new_n889), .ZN(G1345gat));
  AOI21_X1  g689(.A(G155gat), .B1(new_n872), .B2(new_n665), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n246), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n891), .B1(new_n893), .B2(G155gat), .ZN(G1346gat));
  XNOR2_X1  g693(.A(KEYINPUT78), .B(G162gat), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n872), .A2(new_n295), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n892), .A2(new_n675), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(new_n895), .ZN(G1347gat));
  NOR2_X1   g697(.A1(new_n631), .A2(new_n639), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n835), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(G169gat), .B1(new_n900), .B2(new_n822), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n835), .A2(new_n357), .A3(new_n899), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n787), .B2(new_n902), .ZN(G1348gat));
  NOR2_X1   g702(.A1(new_n900), .A2(new_n319), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(new_n297), .ZN(G1349gat));
  NAND4_X1  g704(.A1(new_n835), .A2(new_n665), .A3(new_n377), .A4(new_n899), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n818), .A2(new_n665), .A3(new_n616), .A4(new_n899), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(G183gat), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g709(.A1(new_n835), .A2(new_n295), .A3(new_n899), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n911), .A2(new_n912), .A3(new_n378), .ZN(new_n913));
  XOR2_X1   g712(.A(KEYINPUT61), .B(G190gat), .Z(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n911), .B2(new_n914), .ZN(G1351gat));
  AND2_X1   g714(.A1(new_n657), .A2(new_n899), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n881), .A2(new_n884), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(G197gat), .B1(new_n917), .B2(new_n822), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n818), .A2(new_n572), .A3(new_n657), .A4(new_n899), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n919), .A2(G197gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n918), .B1(new_n787), .B2(new_n920), .ZN(G1352gat));
  INV_X1    g720(.A(new_n919), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n299), .A3(new_n320), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n923), .A2(KEYINPUT62), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n881), .A2(new_n320), .A3(new_n884), .ZN(new_n925));
  INV_X1    g724(.A(new_n916), .ZN(new_n926));
  OAI21_X1  g725(.A(G204gat), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n923), .A2(KEYINPUT62), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n924), .A2(new_n927), .A3(new_n928), .ZN(G1353gat));
  NAND3_X1  g728(.A1(new_n922), .A2(new_n203), .A3(new_n665), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n881), .A2(new_n665), .A3(new_n884), .A4(new_n916), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n931), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n932));
  AOI21_X1  g731(.A(KEYINPUT63), .B1(new_n931), .B2(G211gat), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(G1354gat));
  NAND4_X1  g733(.A1(new_n881), .A2(KEYINPUT127), .A3(new_n884), .A4(new_n916), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n935), .A2(G218gat), .A3(new_n295), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT127), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n917), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n455), .B1(new_n919), .B2(new_n675), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g740(.A(KEYINPUT126), .B(new_n455), .C1(new_n919), .C2(new_n675), .ZN(new_n942));
  AOI22_X1  g741(.A1(new_n936), .A2(new_n938), .B1(new_n941), .B2(new_n942), .ZN(G1355gat));
endmodule


