

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755;

  INV_X1 U372 ( .A(n621), .ZN(n683) );
  NOR2_X1 U373 ( .A1(n667), .A2(n569), .ZN(n563) );
  INV_X1 U374 ( .A(G953), .ZN(n744) );
  XNOR2_X2 U375 ( .A(n689), .B(n425), .ZN(n611) );
  NOR2_X2 U376 ( .A1(n752), .A2(n573), .ZN(n447) );
  XNOR2_X2 U377 ( .A(n415), .B(KEYINPUT35), .ZN(n752) );
  NOR2_X1 U378 ( .A1(n602), .A2(n596), .ZN(n588) );
  XNOR2_X2 U379 ( .A(n614), .B(KEYINPUT38), .ZN(n596) );
  XNOR2_X2 U380 ( .A(n741), .B(G146), .ZN(n524) );
  INV_X2 U381 ( .A(G143), .ZN(n424) );
  NAND2_X1 U382 ( .A1(G234), .A2(G237), .ZN(n549) );
  XNOR2_X1 U383 ( .A(n370), .B(KEYINPUT41), .ZN(n701) );
  NOR2_X1 U384 ( .A1(n590), .A2(n680), .ZN(n591) );
  XNOR2_X1 U385 ( .A(n543), .B(n723), .ZN(n368) );
  NOR2_X1 U386 ( .A1(n423), .A2(n628), .ZN(n663) );
  AND2_X1 U387 ( .A1(n400), .A2(n399), .ZN(n398) );
  NOR2_X1 U388 ( .A1(n428), .A2(n616), .ZN(n656) );
  XNOR2_X1 U389 ( .A(n548), .B(n449), .ZN(n600) );
  NAND2_X2 U390 ( .A1(n376), .A2(n372), .ZN(n689) );
  XNOR2_X1 U391 ( .A(n368), .B(n369), .ZN(n708) );
  XNOR2_X1 U392 ( .A(n582), .B(KEYINPUT79), .ZN(n590) );
  XOR2_X1 U393 ( .A(KEYINPUT72), .B(G137), .Z(n460) );
  XNOR2_X2 U394 ( .A(KEYINPUT4), .B(KEYINPUT65), .ZN(n738) );
  XNOR2_X1 U395 ( .A(n402), .B(n359), .ZN(n571) );
  NOR2_X1 U396 ( .A1(G953), .A2(n699), .ZN(n553) );
  XNOR2_X1 U397 ( .A(n497), .B(n439), .ZN(n567) );
  XNOR2_X1 U398 ( .A(n498), .B(n440), .ZN(n439) );
  INV_X1 U399 ( .A(G475), .ZN(n440) );
  INV_X1 U400 ( .A(G469), .ZN(n527) );
  XNOR2_X1 U401 ( .A(n510), .B(n511), .ZN(n719) );
  XOR2_X1 U402 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n457) );
  INV_X1 U403 ( .A(n659), .ZN(n452) );
  NOR2_X1 U404 ( .A1(n613), .A2(n612), .ZN(n620) );
  NAND2_X1 U405 ( .A1(n611), .A2(n668), .ZN(n612) );
  XNOR2_X1 U406 ( .A(n489), .B(n353), .ZN(n568) );
  OR2_X1 U407 ( .A1(n500), .A2(n373), .ZN(n372) );
  AND2_X1 U408 ( .A1(n378), .A2(n377), .ZN(n376) );
  NAND2_X1 U409 ( .A1(n375), .A2(n374), .ZN(n373) );
  NAND2_X1 U410 ( .A1(n619), .A2(KEYINPUT73), .ZN(n393) );
  OR2_X1 U411 ( .A1(G237), .A2(G902), .ZN(n545) );
  XNOR2_X1 U412 ( .A(G902), .B(KEYINPUT15), .ZN(n544) );
  NOR2_X1 U413 ( .A1(G953), .A2(G237), .ZN(n490) );
  XNOR2_X1 U414 ( .A(n594), .B(n529), .ZN(n621) );
  NAND2_X1 U415 ( .A1(n590), .A2(KEYINPUT78), .ZN(n381) );
  NAND2_X1 U416 ( .A1(n386), .A2(n385), .ZN(n384) );
  XNOR2_X1 U417 ( .A(n443), .B(n441), .ZN(n495) );
  XNOR2_X1 U418 ( .A(n539), .B(n542), .ZN(n369) );
  BUF_X1 U419 ( .A(n621), .Z(n428) );
  NOR2_X2 U420 ( .A1(n600), .A2(n355), .ZN(n448) );
  XNOR2_X1 U421 ( .A(n513), .B(KEYINPUT25), .ZN(n453) );
  OR2_X2 U422 ( .A1(n719), .A2(G902), .ZN(n454) );
  INV_X1 U423 ( .A(n567), .ZN(n438) );
  NAND2_X1 U424 ( .A1(n571), .A2(n428), .ZN(n574) );
  INV_X1 U425 ( .A(KEYINPUT6), .ZN(n425) );
  XNOR2_X1 U426 ( .A(n481), .B(n419), .ZN(n483) );
  XNOR2_X1 U427 ( .A(n525), .B(n526), .ZN(n712) );
  XNOR2_X1 U428 ( .A(n524), .B(n523), .ZN(n525) );
  NOR2_X1 U429 ( .A1(n664), .A2(n663), .ZN(n666) );
  AND2_X1 U430 ( .A1(n649), .A2(KEYINPUT80), .ZN(n437) );
  INV_X1 U431 ( .A(KEYINPUT46), .ZN(n598) );
  XNOR2_X1 U432 ( .A(n685), .B(n418), .ZN(n686) );
  XNOR2_X1 U433 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n418) );
  XNOR2_X1 U434 ( .A(KEYINPUT108), .B(n499), .ZN(n672) );
  OR2_X1 U435 ( .A1(n651), .A2(n653), .ZN(n499) );
  XNOR2_X1 U436 ( .A(n540), .B(n455), .ZN(n509) );
  XNOR2_X1 U437 ( .A(KEYINPUT10), .B(KEYINPUT71), .ZN(n455) );
  XNOR2_X1 U438 ( .A(n444), .B(KEYINPUT11), .ZN(n443) );
  NAND2_X1 U439 ( .A1(n490), .A2(G214), .ZN(n444) );
  XNOR2_X1 U440 ( .A(n491), .B(n442), .ZN(n441) );
  XNOR2_X1 U441 ( .A(G113), .B(G104), .ZN(n491) );
  XNOR2_X1 U442 ( .A(KEYINPUT102), .B(KEYINPUT12), .ZN(n442) );
  XOR2_X1 U443 ( .A(KEYINPUT103), .B(KEYINPUT101), .Z(n493) );
  XNOR2_X1 U444 ( .A(G143), .B(G122), .ZN(n492) );
  XNOR2_X1 U445 ( .A(n456), .B(G125), .ZN(n540) );
  INV_X1 U446 ( .A(G146), .ZN(n456) );
  XNOR2_X1 U447 ( .A(n538), .B(KEYINPUT17), .ZN(n539) );
  XOR2_X1 U448 ( .A(KEYINPUT18), .B(KEYINPUT89), .Z(n537) );
  NAND2_X1 U449 ( .A1(n391), .A2(n350), .ZN(n390) );
  INV_X1 U450 ( .A(KEYINPUT48), .ZN(n401) );
  XNOR2_X1 U451 ( .A(n693), .B(n416), .ZN(n694) );
  XNOR2_X1 U452 ( .A(n417), .B(KEYINPUT51), .ZN(n416) );
  INV_X1 U453 ( .A(KEYINPUT118), .ZN(n417) );
  OR2_X2 U454 ( .A1(n596), .A2(n371), .ZN(n674) );
  INV_X1 U455 ( .A(G902), .ZN(n374) );
  INV_X1 U456 ( .A(G472), .ZN(n375) );
  NAND2_X1 U457 ( .A1(G902), .A2(G472), .ZN(n377) );
  XOR2_X1 U458 ( .A(KEYINPUT76), .B(KEYINPUT99), .Z(n468) );
  INV_X1 U459 ( .A(KEYINPUT5), .ZN(n469) );
  XNOR2_X1 U460 ( .A(G131), .B(KEYINPUT100), .ZN(n470) );
  XNOR2_X1 U461 ( .A(n738), .B(G101), .ZN(n519) );
  XNOR2_X1 U462 ( .A(n518), .B(n517), .ZN(n724) );
  XNOR2_X1 U463 ( .A(G110), .B(G107), .ZN(n517) );
  XOR2_X1 U464 ( .A(KEYINPUT77), .B(G104), .Z(n518) );
  XNOR2_X1 U465 ( .A(n482), .B(n420), .ZN(n419) );
  INV_X1 U466 ( .A(KEYINPUT7), .ZN(n420) );
  XNOR2_X1 U467 ( .A(G116), .B(G107), .ZN(n482) );
  INV_X1 U468 ( .A(G134), .ZN(n435) );
  AND2_X1 U469 ( .A1(n742), .A2(n629), .ZN(n432) );
  INV_X1 U470 ( .A(KEYINPUT94), .ZN(n520) );
  XNOR2_X1 U471 ( .A(n433), .B(n724), .ZN(n543) );
  XNOR2_X1 U472 ( .A(n519), .B(KEYINPUT75), .ZN(n433) );
  NOR2_X1 U473 ( .A1(n732), .A2(KEYINPUT2), .ZN(n660) );
  XNOR2_X1 U474 ( .A(n427), .B(n426), .ZN(n699) );
  INV_X1 U475 ( .A(KEYINPUT91), .ZN(n426) );
  NOR2_X1 U476 ( .A1(n383), .A2(n380), .ZN(n379) );
  INV_X1 U477 ( .A(KEYINPUT19), .ZN(n449) );
  NOR2_X1 U478 ( .A1(n592), .A2(n609), .ZN(n593) );
  NAND2_X1 U479 ( .A1(n623), .A2(n434), .ZN(n659) );
  INV_X1 U480 ( .A(n614), .ZN(n434) );
  INV_X1 U481 ( .A(KEYINPUT40), .ZN(n429) );
  AND2_X1 U482 ( .A1(n620), .A2(n614), .ZN(n615) );
  INV_X1 U483 ( .A(n603), .ZN(n564) );
  NOR2_X1 U484 ( .A1(n574), .A2(n689), .ZN(n572) );
  NOR2_X1 U485 ( .A1(n568), .A2(n438), .ZN(n653) );
  AND2_X1 U486 ( .A1(n568), .A2(n438), .ZN(n651) );
  NOR2_X1 U487 ( .A1(n611), .A2(n574), .ZN(n575) );
  INV_X1 U488 ( .A(KEYINPUT124), .ZN(n412) );
  XNOR2_X1 U489 ( .A(n716), .B(n414), .ZN(n718) );
  XNOR2_X1 U490 ( .A(n717), .B(KEYINPUT122), .ZN(n414) );
  INV_X1 U491 ( .A(KEYINPUT60), .ZN(n404) );
  XNOR2_X1 U492 ( .A(n710), .B(n430), .ZN(n713) );
  INV_X1 U493 ( .A(KEYINPUT56), .ZN(n406) );
  AND2_X1 U494 ( .A1(n705), .A2(n403), .ZN(n706) );
  AND2_X1 U495 ( .A1(n704), .A2(n744), .ZN(n403) );
  NOR2_X1 U496 ( .A1(n619), .A2(KEYINPUT73), .ZN(n350) );
  NOR2_X1 U497 ( .A1(n570), .A2(n451), .ZN(n351) );
  OR2_X1 U498 ( .A1(n560), .A2(n559), .ZN(n352) );
  XOR2_X1 U499 ( .A(KEYINPUT107), .B(G478), .Z(n353) );
  XOR2_X1 U500 ( .A(n506), .B(n505), .Z(n354) );
  AND2_X1 U501 ( .A1(n554), .A2(n581), .ZN(n355) );
  AND2_X1 U502 ( .A1(n637), .A2(n352), .ZN(n356) );
  XOR2_X1 U503 ( .A(G131), .B(G140), .Z(n523) );
  NOR2_X1 U504 ( .A1(n680), .A2(n671), .ZN(n357) );
  NOR2_X1 U505 ( .A1(n751), .A2(n452), .ZN(n358) );
  INV_X1 U506 ( .A(n679), .ZN(n451) );
  XOR2_X1 U507 ( .A(KEYINPUT68), .B(KEYINPUT22), .Z(n359) );
  XOR2_X1 U508 ( .A(KEYINPUT32), .B(KEYINPUT67), .Z(n360) );
  XOR2_X1 U509 ( .A(n555), .B(KEYINPUT0), .Z(n361) );
  XOR2_X1 U510 ( .A(n500), .B(n478), .Z(n362) );
  XOR2_X1 U511 ( .A(n714), .B(n459), .Z(n363) );
  XOR2_X1 U512 ( .A(n708), .B(n707), .Z(n364) );
  XNOR2_X1 U513 ( .A(n719), .B(KEYINPUT123), .ZN(n365) );
  NOR2_X1 U514 ( .A1(G952), .A2(n744), .ZN(n722) );
  INV_X1 U515 ( .A(n722), .ZN(n421) );
  NAND2_X1 U516 ( .A1(n398), .A2(n395), .ZN(n388) );
  XNOR2_X1 U517 ( .A(n387), .B(n401), .ZN(n624) );
  NAND2_X1 U518 ( .A1(n571), .A2(n351), .ZN(n450) );
  NAND2_X1 U519 ( .A1(n389), .A2(n388), .ZN(n387) );
  NAND2_X1 U520 ( .A1(n366), .A2(n679), .ZN(n609) );
  XNOR2_X1 U521 ( .A(n591), .B(KEYINPUT74), .ZN(n366) );
  NAND2_X1 U522 ( .A1(n367), .A2(n606), .ZN(n608) );
  NAND2_X1 U523 ( .A1(n437), .A2(n672), .ZN(n367) );
  NOR2_X1 U524 ( .A1(n708), .A2(n629), .ZN(n547) );
  XNOR2_X2 U525 ( .A(n535), .B(KEYINPUT16), .ZN(n723) );
  INV_X1 U526 ( .A(n596), .ZN(n669) );
  NOR2_X2 U527 ( .A1(n674), .A2(n671), .ZN(n370) );
  INV_X1 U528 ( .A(n668), .ZN(n371) );
  NAND2_X1 U529 ( .A1(n500), .A2(G472), .ZN(n378) );
  NAND2_X1 U530 ( .A1(n379), .A2(n585), .ZN(n602) );
  NAND2_X1 U531 ( .A1(n382), .A2(n381), .ZN(n380) );
  NAND2_X1 U532 ( .A1(n583), .A2(KEYINPUT78), .ZN(n382) );
  NOR2_X1 U533 ( .A1(n583), .A2(n384), .ZN(n383) );
  INV_X1 U534 ( .A(KEYINPUT78), .ZN(n385) );
  INV_X1 U535 ( .A(n590), .ZN(n386) );
  NAND2_X1 U536 ( .A1(n684), .A2(n594), .ZN(n583) );
  NAND2_X1 U537 ( .A1(n392), .A2(n390), .ZN(n389) );
  INV_X1 U538 ( .A(n618), .ZN(n391) );
  AND2_X1 U539 ( .A1(n394), .A2(n393), .ZN(n392) );
  NAND2_X1 U540 ( .A1(n618), .A2(KEYINPUT73), .ZN(n394) );
  NAND2_X1 U541 ( .A1(n397), .A2(n396), .ZN(n395) );
  INV_X1 U542 ( .A(n755), .ZN(n396) );
  NOR2_X1 U543 ( .A1(n754), .A2(n598), .ZN(n397) );
  NAND2_X1 U544 ( .A1(n754), .A2(n598), .ZN(n399) );
  NAND2_X1 U545 ( .A1(n755), .A2(n598), .ZN(n400) );
  NAND2_X1 U546 ( .A1(n557), .A2(n357), .ZN(n402) );
  NAND2_X1 U547 ( .A1(n565), .A2(n564), .ZN(n415) );
  XNOR2_X1 U548 ( .A(n627), .B(KEYINPUT84), .ZN(n423) );
  XNOR2_X1 U549 ( .A(n405), .B(n404), .ZN(G60) );
  NAND2_X1 U550 ( .A1(n409), .A2(n421), .ZN(n405) );
  XNOR2_X1 U551 ( .A(n407), .B(n406), .ZN(G51) );
  NAND2_X1 U552 ( .A1(n410), .A2(n421), .ZN(n407) );
  XNOR2_X1 U553 ( .A(n408), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U554 ( .A1(n411), .A2(n421), .ZN(n408) );
  XNOR2_X1 U555 ( .A(n715), .B(n363), .ZN(n409) );
  XNOR2_X1 U556 ( .A(n709), .B(n364), .ZN(n410) );
  XNOR2_X1 U557 ( .A(n636), .B(n362), .ZN(n411) );
  XNOR2_X1 U558 ( .A(n413), .B(n412), .ZN(G66) );
  NAND2_X1 U559 ( .A1(n422), .A2(n421), .ZN(n413) );
  XNOR2_X2 U560 ( .A(n448), .B(n361), .ZN(n557) );
  NOR2_X2 U561 ( .A1(G902), .A2(n712), .ZN(n528) );
  NOR2_X1 U562 ( .A1(n566), .A2(n561), .ZN(n562) );
  XNOR2_X1 U563 ( .A(n721), .B(n365), .ZN(n422) );
  INV_X1 U564 ( .A(n557), .ZN(n569) );
  BUF_X2 U565 ( .A(n586), .Z(n614) );
  XNOR2_X2 U566 ( .A(n424), .B(G128), .ZN(n541) );
  XNOR2_X2 U567 ( .A(n445), .B(n577), .ZN(n732) );
  NAND2_X1 U568 ( .A1(n586), .A2(n668), .ZN(n548) );
  XNOR2_X1 U569 ( .A(n547), .B(n546), .ZN(n586) );
  NAND2_X1 U570 ( .A1(n552), .A2(G952), .ZN(n427) );
  XNOR2_X2 U571 ( .A(n589), .B(n429), .ZN(n755) );
  XNOR2_X1 U572 ( .A(n712), .B(n711), .ZN(n430) );
  NAND2_X1 U573 ( .A1(n617), .A2(n431), .ZN(n618) );
  XNOR2_X1 U574 ( .A(n656), .B(KEYINPUT85), .ZN(n431) );
  NAND2_X1 U575 ( .A1(n432), .A2(n732), .ZN(n632) );
  XNOR2_X2 U576 ( .A(n484), .B(n460), .ZN(n741) );
  XNOR2_X2 U577 ( .A(n541), .B(n435), .ZN(n484) );
  NAND2_X1 U578 ( .A1(n672), .A2(n436), .ZN(n607) );
  AND2_X1 U579 ( .A1(n649), .A2(KEYINPUT47), .ZN(n436) );
  NAND2_X1 U580 ( .A1(n446), .A2(n356), .ZN(n445) );
  XNOR2_X1 U581 ( .A(n447), .B(KEYINPUT44), .ZN(n446) );
  XNOR2_X2 U582 ( .A(n450), .B(n360), .ZN(n753) );
  AND2_X2 U583 ( .A1(n624), .A2(n358), .ZN(n742) );
  NOR2_X2 U584 ( .A1(n599), .A2(n600), .ZN(n649) );
  XNOR2_X2 U585 ( .A(n454), .B(n453), .ZN(n679) );
  XNOR2_X1 U586 ( .A(n509), .B(n457), .ZN(n510) );
  XNOR2_X1 U587 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U588 ( .A(n496), .B(n737), .ZN(n714) );
  XNOR2_X1 U589 ( .A(n543), .B(n522), .ZN(n526) );
  XNOR2_X1 U590 ( .A(KEYINPUT36), .B(KEYINPUT87), .ZN(n458) );
  XNOR2_X1 U591 ( .A(KEYINPUT59), .B(KEYINPUT121), .ZN(n459) );
  XNOR2_X1 U592 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U593 ( .A(n472), .B(n471), .ZN(n473) );
  INV_X1 U594 ( .A(KEYINPUT88), .ZN(n555) );
  XNOR2_X1 U595 ( .A(n521), .B(n520), .ZN(n522) );
  INV_X1 U596 ( .A(KEYINPUT39), .ZN(n587) );
  INV_X1 U597 ( .A(G116), .ZN(n461) );
  NAND2_X1 U598 ( .A1(G113), .A2(n461), .ZN(n464) );
  INV_X1 U599 ( .A(G113), .ZN(n462) );
  NAND2_X1 U600 ( .A1(n462), .A2(G116), .ZN(n463) );
  NAND2_X1 U601 ( .A1(n464), .A2(n463), .ZN(n466) );
  XNOR2_X1 U602 ( .A(KEYINPUT3), .B(G119), .ZN(n465) );
  XNOR2_X1 U603 ( .A(n466), .B(n465), .ZN(n530) );
  XNOR2_X1 U604 ( .A(n519), .B(n530), .ZN(n474) );
  NAND2_X1 U605 ( .A1(n490), .A2(G210), .ZN(n467) );
  XNOR2_X1 U606 ( .A(n468), .B(n467), .ZN(n472) );
  XNOR2_X1 U607 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U608 ( .A(n524), .B(n475), .ZN(n500) );
  XOR2_X1 U609 ( .A(KEYINPUT90), .B(KEYINPUT111), .Z(n477) );
  XNOR2_X1 U610 ( .A(KEYINPUT62), .B(KEYINPUT110), .ZN(n476) );
  XNOR2_X1 U611 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U612 ( .A(KEYINPUT105), .B(KEYINPUT9), .Z(n480) );
  XNOR2_X1 U613 ( .A(G122), .B(KEYINPUT106), .ZN(n479) );
  XNOR2_X1 U614 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U615 ( .A(n484), .B(n483), .Z(n488) );
  XOR2_X1 U616 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n486) );
  NAND2_X1 U617 ( .A1(G234), .A2(n744), .ZN(n485) );
  XNOR2_X1 U618 ( .A(n486), .B(n485), .ZN(n507) );
  NAND2_X1 U619 ( .A1(G217), .A2(n507), .ZN(n487) );
  XNOR2_X1 U620 ( .A(n488), .B(n487), .ZN(n717) );
  NOR2_X1 U621 ( .A1(G902), .A2(n717), .ZN(n489) );
  XNOR2_X1 U622 ( .A(KEYINPUT13), .B(KEYINPUT104), .ZN(n498) );
  XNOR2_X1 U623 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U624 ( .A(n509), .B(n523), .Z(n737) );
  NOR2_X1 U625 ( .A1(G902), .A2(n714), .ZN(n497) );
  XOR2_X1 U626 ( .A(n672), .B(KEYINPUT80), .Z(n560) );
  INV_X1 U627 ( .A(n689), .ZN(n592) );
  XOR2_X1 U628 ( .A(G110), .B(G119), .Z(n502) );
  XNOR2_X1 U629 ( .A(G128), .B(G137), .ZN(n501) );
  XNOR2_X1 U630 ( .A(n502), .B(n501), .ZN(n506) );
  XOR2_X1 U631 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n504) );
  XNOR2_X1 U632 ( .A(G140), .B(KEYINPUT97), .ZN(n503) );
  XNOR2_X1 U633 ( .A(n504), .B(n503), .ZN(n505) );
  NAND2_X1 U634 ( .A1(n507), .A2(G221), .ZN(n508) );
  XNOR2_X1 U635 ( .A(n354), .B(n508), .ZN(n511) );
  NAND2_X1 U636 ( .A1(G234), .A2(n544), .ZN(n512) );
  XNOR2_X1 U637 ( .A(KEYINPUT20), .B(n512), .ZN(n514) );
  NAND2_X1 U638 ( .A1(G217), .A2(n514), .ZN(n513) );
  NAND2_X1 U639 ( .A1(n514), .A2(G221), .ZN(n515) );
  XOR2_X1 U640 ( .A(KEYINPUT98), .B(n515), .Z(n516) );
  XOR2_X1 U641 ( .A(KEYINPUT21), .B(n516), .Z(n680) );
  NOR2_X1 U642 ( .A1(n679), .A2(n680), .ZN(n684) );
  NAND2_X1 U643 ( .A1(G227), .A2(n744), .ZN(n521) );
  XNOR2_X2 U644 ( .A(n528), .B(n527), .ZN(n594) );
  XNOR2_X1 U645 ( .A(KEYINPUT1), .B(KEYINPUT69), .ZN(n529) );
  NAND2_X1 U646 ( .A1(n684), .A2(n683), .ZN(n561) );
  NOR2_X1 U647 ( .A1(n592), .A2(n561), .ZN(n692) );
  NAND2_X1 U648 ( .A1(G214), .A2(n545), .ZN(n668) );
  NAND2_X1 U649 ( .A1(n530), .A2(G122), .ZN(n534) );
  INV_X1 U650 ( .A(n530), .ZN(n532) );
  INV_X1 U651 ( .A(G122), .ZN(n531) );
  NAND2_X1 U652 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U653 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U654 ( .A1(G224), .A2(n744), .ZN(n536) );
  XOR2_X1 U655 ( .A(n537), .B(n536), .Z(n538) );
  XNOR2_X1 U656 ( .A(n541), .B(n540), .ZN(n542) );
  INV_X1 U657 ( .A(n544), .ZN(n629) );
  NAND2_X1 U658 ( .A1(G210), .A2(n545), .ZN(n546) );
  XNOR2_X1 U659 ( .A(n549), .B(KEYINPUT14), .ZN(n552) );
  NAND2_X1 U660 ( .A1(G902), .A2(n552), .ZN(n578) );
  INV_X1 U661 ( .A(n578), .ZN(n550) );
  NOR2_X1 U662 ( .A1(G898), .A2(n744), .ZN(n727) );
  NAND2_X1 U663 ( .A1(n550), .A2(n727), .ZN(n551) );
  XOR2_X1 U664 ( .A(KEYINPUT93), .B(n551), .Z(n554) );
  XOR2_X1 U665 ( .A(KEYINPUT92), .B(n553), .Z(n581) );
  NAND2_X1 U666 ( .A1(n692), .A2(n557), .ZN(n556) );
  XNOR2_X1 U667 ( .A(n556), .B(KEYINPUT31), .ZN(n654) );
  OR2_X1 U668 ( .A1(n569), .A2(n583), .ZN(n558) );
  NOR2_X1 U669 ( .A1(n689), .A2(n558), .ZN(n639) );
  NOR2_X1 U670 ( .A1(n654), .A2(n639), .ZN(n559) );
  INV_X1 U671 ( .A(n611), .ZN(n566) );
  XNOR2_X1 U672 ( .A(n562), .B(KEYINPUT33), .ZN(n667) );
  XNOR2_X1 U673 ( .A(n563), .B(KEYINPUT34), .ZN(n565) );
  OR2_X1 U674 ( .A1(n568), .A2(n567), .ZN(n603) );
  NAND2_X1 U675 ( .A1(n566), .A2(n683), .ZN(n570) );
  NAND2_X1 U676 ( .A1(n568), .A2(n567), .ZN(n671) );
  NAND2_X1 U677 ( .A1(n679), .A2(n572), .ZN(n643) );
  NAND2_X1 U678 ( .A1(n753), .A2(n643), .ZN(n573) );
  XNOR2_X1 U679 ( .A(n575), .B(KEYINPUT86), .ZN(n576) );
  NAND2_X1 U680 ( .A1(n576), .A2(n451), .ZN(n637) );
  XNOR2_X1 U681 ( .A(KEYINPUT45), .B(KEYINPUT64), .ZN(n577) );
  INV_X1 U682 ( .A(n732), .ZN(n628) );
  NOR2_X1 U683 ( .A1(G900), .A2(n578), .ZN(n579) );
  NAND2_X1 U684 ( .A1(G953), .A2(n579), .ZN(n580) );
  NAND2_X1 U685 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U686 ( .A1(n689), .A2(n668), .ZN(n584) );
  XOR2_X1 U687 ( .A(KEYINPUT30), .B(n584), .Z(n585) );
  XNOR2_X1 U688 ( .A(n588), .B(n587), .ZN(n625) );
  NAND2_X1 U689 ( .A1(n625), .A2(n651), .ZN(n589) );
  XNOR2_X1 U690 ( .A(KEYINPUT28), .B(n593), .ZN(n595) );
  NAND2_X1 U691 ( .A1(n595), .A2(n594), .ZN(n599) );
  NOR2_X1 U692 ( .A1(n599), .A2(n701), .ZN(n597) );
  XNOR2_X1 U693 ( .A(n597), .B(KEYINPUT42), .ZN(n754) );
  NOR2_X1 U694 ( .A1(n672), .A2(KEYINPUT80), .ZN(n601) );
  NAND2_X1 U695 ( .A1(n601), .A2(n649), .ZN(n605) );
  NOR2_X1 U696 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U697 ( .A1(n614), .A2(n604), .ZN(n648) );
  NAND2_X1 U698 ( .A1(n605), .A2(n648), .ZN(n619) );
  INV_X1 U699 ( .A(KEYINPUT47), .ZN(n606) );
  NAND2_X1 U700 ( .A1(n608), .A2(n607), .ZN(n617) );
  INV_X1 U701 ( .A(n609), .ZN(n610) );
  NAND2_X1 U702 ( .A1(n651), .A2(n610), .ZN(n613) );
  XNOR2_X1 U703 ( .A(n615), .B(n458), .ZN(n616) );
  NAND2_X1 U704 ( .A1(n428), .A2(n620), .ZN(n622) );
  XNOR2_X1 U705 ( .A(n622), .B(KEYINPUT43), .ZN(n623) );
  AND2_X1 U706 ( .A1(n625), .A2(n653), .ZN(n626) );
  XOR2_X1 U707 ( .A(KEYINPUT109), .B(n626), .Z(n751) );
  NAND2_X1 U708 ( .A1(n742), .A2(KEYINPUT2), .ZN(n627) );
  INV_X1 U709 ( .A(n663), .ZN(n635) );
  XOR2_X1 U710 ( .A(n629), .B(KEYINPUT83), .Z(n630) );
  NAND2_X1 U711 ( .A1(n630), .A2(KEYINPUT2), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U713 ( .A(n633), .B(KEYINPUT66), .ZN(n634) );
  AND2_X2 U714 ( .A1(n635), .A2(n634), .ZN(n720) );
  NAND2_X1 U715 ( .A1(n720), .A2(G472), .ZN(n636) );
  XNOR2_X1 U716 ( .A(G101), .B(n637), .ZN(G3) );
  NAND2_X1 U717 ( .A1(n639), .A2(n651), .ZN(n638) );
  XNOR2_X1 U718 ( .A(n638), .B(G104), .ZN(G6) );
  XOR2_X1 U719 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n641) );
  NAND2_X1 U720 ( .A1(n639), .A2(n653), .ZN(n640) );
  XNOR2_X1 U721 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U722 ( .A(G107), .B(n642), .ZN(G9) );
  XNOR2_X1 U723 ( .A(G110), .B(KEYINPUT112), .ZN(n644) );
  XNOR2_X1 U724 ( .A(n644), .B(n643), .ZN(G12) );
  XOR2_X1 U725 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n646) );
  NAND2_X1 U726 ( .A1(n649), .A2(n653), .ZN(n645) );
  XNOR2_X1 U727 ( .A(n646), .B(n645), .ZN(n647) );
  XOR2_X1 U728 ( .A(G128), .B(n647), .Z(G30) );
  XNOR2_X1 U729 ( .A(G143), .B(n648), .ZN(G45) );
  NAND2_X1 U730 ( .A1(n649), .A2(n651), .ZN(n650) );
  XNOR2_X1 U731 ( .A(n650), .B(G146), .ZN(G48) );
  NAND2_X1 U732 ( .A1(n654), .A2(n651), .ZN(n652) );
  XNOR2_X1 U733 ( .A(n652), .B(G113), .ZN(G15) );
  NAND2_X1 U734 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U735 ( .A(n655), .B(G116), .ZN(G18) );
  XNOR2_X1 U736 ( .A(n656), .B(KEYINPUT114), .ZN(n657) );
  XNOR2_X1 U737 ( .A(n657), .B(KEYINPUT37), .ZN(n658) );
  XNOR2_X1 U738 ( .A(G125), .B(n658), .ZN(G27) );
  XNOR2_X1 U739 ( .A(G140), .B(n659), .ZN(G42) );
  XNOR2_X1 U740 ( .A(n660), .B(KEYINPUT81), .ZN(n662) );
  OR2_X1 U741 ( .A1(KEYINPUT2), .A2(n742), .ZN(n661) );
  NAND2_X1 U742 ( .A1(n662), .A2(n661), .ZN(n664) );
  INV_X1 U743 ( .A(KEYINPUT82), .ZN(n665) );
  XNOR2_X1 U744 ( .A(n666), .B(n665), .ZN(n705) );
  NOR2_X1 U745 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U746 ( .A1(n671), .A2(n670), .ZN(n676) );
  INV_X1 U747 ( .A(n672), .ZN(n673) );
  NOR2_X1 U748 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U749 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U750 ( .A(KEYINPUT119), .B(n677), .Z(n678) );
  NOR2_X1 U751 ( .A1(n667), .A2(n678), .ZN(n696) );
  NAND2_X1 U752 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U753 ( .A(n681), .B(KEYINPUT49), .ZN(n682) );
  XNOR2_X1 U754 ( .A(KEYINPUT115), .B(n682), .ZN(n687) );
  OR2_X1 U755 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U756 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U757 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U758 ( .A(KEYINPUT117), .B(n690), .Z(n691) );
  NOR2_X1 U759 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U760 ( .A1(n701), .A2(n694), .ZN(n695) );
  NOR2_X1 U761 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U762 ( .A(n697), .B(KEYINPUT52), .ZN(n698) );
  NOR2_X1 U763 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U764 ( .A(n700), .B(KEYINPUT120), .ZN(n703) );
  NOR2_X1 U765 ( .A1(n667), .A2(n701), .ZN(n702) );
  NOR2_X1 U766 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U767 ( .A(n706), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U768 ( .A1(n720), .A2(G210), .ZN(n709) );
  XOR2_X1 U769 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n707) );
  XOR2_X1 U770 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n711) );
  NAND2_X1 U771 ( .A1(n720), .A2(G469), .ZN(n710) );
  NOR2_X1 U772 ( .A1(n722), .A2(n713), .ZN(G54) );
  NAND2_X1 U773 ( .A1(n720), .A2(G475), .ZN(n715) );
  NAND2_X1 U774 ( .A1(n720), .A2(G478), .ZN(n716) );
  NOR2_X1 U775 ( .A1(n722), .A2(n718), .ZN(G63) );
  NAND2_X1 U776 ( .A1(n720), .A2(G217), .ZN(n721) );
  XOR2_X1 U777 ( .A(KEYINPUT126), .B(n723), .Z(n726) );
  XNOR2_X1 U778 ( .A(G101), .B(n724), .ZN(n725) );
  XNOR2_X1 U779 ( .A(n726), .B(n725), .ZN(n728) );
  NOR2_X1 U780 ( .A1(n728), .A2(n727), .ZN(n736) );
  XOR2_X1 U781 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n730) );
  NAND2_X1 U782 ( .A1(G224), .A2(G953), .ZN(n729) );
  XNOR2_X1 U783 ( .A(n730), .B(n729), .ZN(n731) );
  NAND2_X1 U784 ( .A1(n731), .A2(G898), .ZN(n734) );
  NAND2_X1 U785 ( .A1(n732), .A2(n744), .ZN(n733) );
  NAND2_X1 U786 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U787 ( .A(n736), .B(n735), .ZN(G69) );
  XNOR2_X1 U788 ( .A(n737), .B(KEYINPUT127), .ZN(n739) );
  XNOR2_X1 U789 ( .A(n738), .B(n739), .ZN(n740) );
  XOR2_X1 U790 ( .A(n741), .B(n740), .Z(n746) );
  INV_X1 U791 ( .A(n746), .ZN(n743) );
  XOR2_X1 U792 ( .A(n743), .B(n742), .Z(n745) );
  NAND2_X1 U793 ( .A1(n745), .A2(n744), .ZN(n750) );
  XOR2_X1 U794 ( .A(G227), .B(n746), .Z(n747) );
  NAND2_X1 U795 ( .A1(n747), .A2(G900), .ZN(n748) );
  NAND2_X1 U796 ( .A1(n748), .A2(G953), .ZN(n749) );
  NAND2_X1 U797 ( .A1(n750), .A2(n749), .ZN(G72) );
  XOR2_X1 U798 ( .A(G134), .B(n751), .Z(G36) );
  XOR2_X1 U799 ( .A(n752), .B(G122), .Z(G24) );
  XNOR2_X1 U800 ( .A(G119), .B(n753), .ZN(G21) );
  XOR2_X1 U801 ( .A(n754), .B(G137), .Z(G39) );
  XOR2_X1 U802 ( .A(n755), .B(G131), .Z(G33) );
endmodule

