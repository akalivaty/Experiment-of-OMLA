

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584;

  NOR2_X1 U324 ( .A1(n567), .A2(n466), .ZN(n547) );
  XOR2_X1 U325 ( .A(n337), .B(n336), .Z(n573) );
  XNOR2_X2 U326 ( .A(n451), .B(KEYINPUT121), .ZN(n561) );
  NAND2_X1 U327 ( .A1(n509), .A2(n568), .ZN(n358) );
  XNOR2_X1 U328 ( .A(n573), .B(n338), .ZN(n509) );
  XNOR2_X1 U329 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n342) );
  XNOR2_X1 U330 ( .A(n471), .B(KEYINPUT37), .ZN(n472) );
  XOR2_X1 U331 ( .A(n374), .B(n373), .Z(n557) );
  XNOR2_X1 U332 ( .A(n411), .B(n410), .ZN(n546) );
  XOR2_X1 U333 ( .A(n332), .B(n331), .Z(n292) );
  XNOR2_X1 U334 ( .A(KEYINPUT45), .B(KEYINPUT115), .ZN(n377) );
  INV_X1 U335 ( .A(KEYINPUT8), .ZN(n343) );
  XNOR2_X1 U336 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U337 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U338 ( .A(n346), .B(n345), .ZN(n370) );
  INV_X1 U339 ( .A(KEYINPUT104), .ZN(n471) );
  XNOR2_X1 U340 ( .A(n333), .B(n292), .ZN(n334) );
  INV_X1 U341 ( .A(KEYINPUT41), .ZN(n338) );
  XNOR2_X1 U342 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U343 ( .A(n473), .B(n472), .ZN(n521) );
  XOR2_X1 U344 ( .A(n330), .B(n304), .Z(n523) );
  XOR2_X1 U345 ( .A(KEYINPUT106), .B(n477), .Z(n506) );
  XNOR2_X1 U346 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n481) );
  XNOR2_X1 U347 ( .A(n478), .B(G43GAT), .ZN(n479) );
  XNOR2_X1 U348 ( .A(n482), .B(n481), .ZN(G1351GAT) );
  XNOR2_X1 U349 ( .A(n480), .B(n479), .ZN(G1330GAT) );
  XNOR2_X1 U350 ( .A(G176GAT), .B(G92GAT), .ZN(n293) );
  XNOR2_X1 U351 ( .A(n293), .B(G64GAT), .ZN(n330) );
  XOR2_X1 U352 ( .A(G169GAT), .B(G8GAT), .Z(n354) );
  XOR2_X1 U353 ( .A(G190GAT), .B(KEYINPUT76), .Z(n363) );
  XNOR2_X1 U354 ( .A(n354), .B(n363), .ZN(n303) );
  XOR2_X1 U355 ( .A(G218GAT), .B(G204GAT), .Z(n295) );
  NAND2_X1 U356 ( .A1(G226GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U357 ( .A(n295), .B(n294), .ZN(n297) );
  XNOR2_X1 U358 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n296) );
  XNOR2_X1 U359 ( .A(n296), .B(G211GAT), .ZN(n422) );
  XOR2_X1 U360 ( .A(n297), .B(n422), .Z(n301) );
  XOR2_X1 U361 ( .A(G183GAT), .B(KEYINPUT19), .Z(n299) );
  XNOR2_X1 U362 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n298) );
  XNOR2_X1 U363 ( .A(n299), .B(n298), .ZN(n443) );
  XNOR2_X1 U364 ( .A(n443), .B(G36GAT), .ZN(n300) );
  XNOR2_X1 U365 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U366 ( .A(n303), .B(n302), .ZN(n304) );
  INV_X1 U367 ( .A(n523), .ZN(n454) );
  XOR2_X1 U368 ( .A(G211GAT), .B(G155GAT), .Z(n306) );
  XNOR2_X1 U369 ( .A(G22GAT), .B(G78GAT), .ZN(n305) );
  XNOR2_X1 U370 ( .A(n306), .B(n305), .ZN(n310) );
  XOR2_X1 U371 ( .A(G71GAT), .B(G183GAT), .Z(n308) );
  XNOR2_X1 U372 ( .A(G8GAT), .B(G127GAT), .ZN(n307) );
  XNOR2_X1 U373 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U374 ( .A(n310), .B(n309), .Z(n315) );
  XOR2_X1 U375 ( .A(KEYINPUT77), .B(KEYINPUT79), .Z(n312) );
  NAND2_X1 U376 ( .A1(G231GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U377 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U378 ( .A(KEYINPUT78), .B(n313), .ZN(n314) );
  XNOR2_X1 U379 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U380 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n317) );
  XNOR2_X1 U381 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n316) );
  XNOR2_X1 U382 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U383 ( .A(n319), .B(n318), .Z(n323) );
  XNOR2_X1 U384 ( .A(G15GAT), .B(G1GAT), .ZN(n320) );
  XNOR2_X1 U385 ( .A(n320), .B(KEYINPUT69), .ZN(n352) );
  XNOR2_X1 U386 ( .A(G57GAT), .B(KEYINPUT72), .ZN(n321) );
  XNOR2_X1 U387 ( .A(n321), .B(KEYINPUT13), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n352), .B(n329), .ZN(n322) );
  XNOR2_X1 U389 ( .A(n323), .B(n322), .ZN(n576) );
  XOR2_X1 U390 ( .A(G120GAT), .B(G71GAT), .Z(n436) );
  XOR2_X1 U391 ( .A(G99GAT), .B(G85GAT), .Z(n361) );
  INV_X1 U392 ( .A(n361), .ZN(n324) );
  XOR2_X1 U393 ( .A(n436), .B(n324), .Z(n337) );
  XOR2_X1 U394 ( .A(G78GAT), .B(G148GAT), .Z(n326) );
  XNOR2_X1 U395 ( .A(G106GAT), .B(G204GAT), .ZN(n325) );
  XNOR2_X1 U396 ( .A(n326), .B(n325), .ZN(n419) );
  XNOR2_X1 U397 ( .A(n419), .B(KEYINPUT74), .ZN(n328) );
  AND2_X1 U398 ( .A1(G230GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U399 ( .A(n328), .B(n327), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n330), .B(n329), .ZN(n333) );
  XOR2_X1 U401 ( .A(KEYINPUT73), .B(KEYINPUT33), .Z(n332) );
  XNOR2_X1 U402 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n331) );
  XOR2_X1 U403 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n340) );
  NAND2_X1 U404 ( .A1(G229GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U405 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U406 ( .A(n341), .B(KEYINPUT68), .Z(n351) );
  XNOR2_X1 U407 ( .A(n342), .B(G29GAT), .ZN(n346) );
  XNOR2_X1 U408 ( .A(G43GAT), .B(G50GAT), .ZN(n344) );
  XOR2_X1 U409 ( .A(KEYINPUT70), .B(KEYINPUT67), .Z(n348) );
  XNOR2_X1 U410 ( .A(G197GAT), .B(G113GAT), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n370), .B(n349), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n351), .B(n350), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n356) );
  XOR2_X1 U415 ( .A(G141GAT), .B(G22GAT), .Z(n425) );
  XNOR2_X1 U416 ( .A(n425), .B(n354), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n510) );
  INV_X1 U418 ( .A(n510), .ZN(n568) );
  XOR2_X1 U419 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n357) );
  XOR2_X1 U420 ( .A(n358), .B(n357), .Z(n359) );
  NOR2_X1 U421 ( .A1(n576), .A2(n359), .ZN(n360) );
  XNOR2_X1 U422 ( .A(n360), .B(KEYINPUT114), .ZN(n375) );
  XNOR2_X1 U423 ( .A(G106GAT), .B(G92GAT), .ZN(n362) );
  XOR2_X1 U424 ( .A(n362), .B(n361), .Z(n374) );
  XOR2_X1 U425 ( .A(G134GAT), .B(KEYINPUT75), .Z(n394) );
  XOR2_X1 U426 ( .A(n363), .B(n394), .Z(n365) );
  NAND2_X1 U427 ( .A1(G232GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U428 ( .A(n365), .B(n364), .ZN(n369) );
  XOR2_X1 U429 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n367) );
  XNOR2_X1 U430 ( .A(KEYINPUT65), .B(KEYINPUT9), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U432 ( .A(n369), .B(n368), .Z(n372) );
  XOR2_X1 U433 ( .A(G218GAT), .B(G162GAT), .Z(n424) );
  XNOR2_X1 U434 ( .A(n370), .B(n424), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n373) );
  INV_X1 U436 ( .A(n557), .ZN(n483) );
  NAND2_X1 U437 ( .A1(n375), .A2(n483), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n376), .B(KEYINPUT47), .ZN(n382) );
  XOR2_X1 U439 ( .A(KEYINPUT36), .B(n483), .Z(n579) );
  NAND2_X1 U440 ( .A1(n576), .A2(n579), .ZN(n378) );
  INV_X1 U441 ( .A(n573), .ZN(n474) );
  NAND2_X1 U442 ( .A1(n379), .A2(n474), .ZN(n380) );
  XNOR2_X1 U443 ( .A(n510), .B(KEYINPUT71), .ZN(n559) );
  NOR2_X1 U444 ( .A1(n380), .A2(n559), .ZN(n381) );
  NOR2_X1 U445 ( .A1(n382), .A2(n381), .ZN(n385) );
  XNOR2_X1 U446 ( .A(KEYINPUT64), .B(KEYINPUT116), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n383), .B(KEYINPUT48), .ZN(n384) );
  XNOR2_X1 U448 ( .A(n385), .B(n384), .ZN(n549) );
  NOR2_X1 U449 ( .A1(n454), .A2(n549), .ZN(n386) );
  XOR2_X1 U450 ( .A(KEYINPUT54), .B(n386), .Z(n412) );
  XOR2_X1 U451 ( .A(G57GAT), .B(G120GAT), .Z(n388) );
  XNOR2_X1 U452 ( .A(G141GAT), .B(G1GAT), .ZN(n387) );
  XNOR2_X1 U453 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U454 ( .A(G85GAT), .B(G162GAT), .Z(n390) );
  XNOR2_X1 U455 ( .A(G29GAT), .B(G148GAT), .ZN(n389) );
  XNOR2_X1 U456 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U457 ( .A(n392), .B(n391), .ZN(n411) );
  XNOR2_X1 U458 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n393) );
  XNOR2_X1 U459 ( .A(n393), .B(G127GAT), .ZN(n445) );
  XOR2_X1 U460 ( .A(n394), .B(n445), .Z(n396) );
  NAND2_X1 U461 ( .A1(G225GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U462 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U463 ( .A(n397), .B(KEYINPUT92), .Z(n401) );
  XOR2_X1 U464 ( .A(G155GAT), .B(KEYINPUT87), .Z(n399) );
  XNOR2_X1 U465 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n398) );
  XNOR2_X1 U466 ( .A(n399), .B(n398), .ZN(n418) );
  XNOR2_X1 U467 ( .A(n418), .B(KEYINPUT91), .ZN(n400) );
  XNOR2_X1 U468 ( .A(n401), .B(n400), .ZN(n409) );
  XOR2_X1 U469 ( .A(KEYINPUT90), .B(KEYINPUT94), .Z(n403) );
  XNOR2_X1 U470 ( .A(KEYINPUT1), .B(KEYINPUT89), .ZN(n402) );
  XNOR2_X1 U471 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U472 ( .A(KEYINPUT93), .B(KEYINPUT6), .Z(n405) );
  XNOR2_X1 U473 ( .A(KEYINPUT4), .B(KEYINPUT5), .ZN(n404) );
  XNOR2_X1 U474 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U475 ( .A(n407), .B(n406), .Z(n408) );
  XNOR2_X1 U476 ( .A(n409), .B(n408), .ZN(n410) );
  NOR2_X2 U477 ( .A1(n412), .A2(n546), .ZN(n565) );
  XOR2_X1 U478 ( .A(KEYINPUT88), .B(KEYINPUT24), .Z(n414) );
  XNOR2_X1 U479 ( .A(G50GAT), .B(KEYINPUT85), .ZN(n413) );
  XOR2_X1 U480 ( .A(n414), .B(n413), .Z(n429) );
  XOR2_X1 U481 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n416) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U483 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U484 ( .A(n417), .B(KEYINPUT86), .Z(n421) );
  XNOR2_X1 U485 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U486 ( .A(n421), .B(n420), .ZN(n423) );
  XOR2_X1 U487 ( .A(n423), .B(n422), .Z(n427) );
  XNOR2_X1 U488 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U489 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U490 ( .A(n429), .B(n428), .ZN(n464) );
  NAND2_X1 U491 ( .A1(n565), .A2(n464), .ZN(n430) );
  XNOR2_X1 U492 ( .A(n430), .B(KEYINPUT55), .ZN(n450) );
  XOR2_X1 U493 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n432) );
  XNOR2_X1 U494 ( .A(KEYINPUT81), .B(KEYINPUT20), .ZN(n431) );
  XNOR2_X1 U495 ( .A(n432), .B(n431), .ZN(n440) );
  XOR2_X1 U496 ( .A(KEYINPUT80), .B(G99GAT), .Z(n434) );
  XNOR2_X1 U497 ( .A(G15GAT), .B(G134GAT), .ZN(n433) );
  XNOR2_X1 U498 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U499 ( .A(n435), .B(G190GAT), .Z(n438) );
  XNOR2_X1 U500 ( .A(G43GAT), .B(n436), .ZN(n437) );
  XNOR2_X1 U501 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U502 ( .A(n440), .B(n439), .ZN(n449) );
  XOR2_X1 U503 ( .A(KEYINPUT82), .B(G176GAT), .Z(n442) );
  NAND2_X1 U504 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U505 ( .A(n442), .B(n441), .ZN(n444) );
  XOR2_X1 U506 ( .A(n444), .B(n443), .Z(n447) );
  XNOR2_X1 U507 ( .A(G169GAT), .B(n445), .ZN(n446) );
  XNOR2_X1 U508 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U509 ( .A(n449), .B(n448), .Z(n532) );
  INV_X1 U510 ( .A(n532), .ZN(n525) );
  NAND2_X1 U511 ( .A1(n450), .A2(n525), .ZN(n451) );
  NAND2_X1 U512 ( .A1(n561), .A2(n576), .ZN(n453) );
  XNOR2_X1 U513 ( .A(KEYINPUT122), .B(G183GAT), .ZN(n452) );
  XNOR2_X1 U514 ( .A(n453), .B(n452), .ZN(G1350GAT) );
  NOR2_X1 U515 ( .A1(n532), .A2(n454), .ZN(n455) );
  XNOR2_X1 U516 ( .A(KEYINPUT97), .B(n455), .ZN(n456) );
  NAND2_X1 U517 ( .A1(n456), .A2(n464), .ZN(n457) );
  XNOR2_X1 U518 ( .A(KEYINPUT25), .B(n457), .ZN(n461) );
  XNOR2_X1 U519 ( .A(KEYINPUT26), .B(KEYINPUT95), .ZN(n459) );
  NOR2_X1 U520 ( .A1(n525), .A2(n464), .ZN(n458) );
  XNOR2_X1 U521 ( .A(n459), .B(n458), .ZN(n567) );
  XOR2_X1 U522 ( .A(KEYINPUT27), .B(n523), .Z(n466) );
  XNOR2_X1 U523 ( .A(KEYINPUT96), .B(n547), .ZN(n460) );
  NOR2_X1 U524 ( .A1(n461), .A2(n460), .ZN(n462) );
  NOR2_X1 U525 ( .A1(n462), .A2(n546), .ZN(n463) );
  XNOR2_X1 U526 ( .A(n463), .B(KEYINPUT98), .ZN(n469) );
  XOR2_X1 U527 ( .A(n464), .B(KEYINPUT66), .Z(n465) );
  XNOR2_X1 U528 ( .A(KEYINPUT28), .B(n465), .ZN(n529) );
  NOR2_X1 U529 ( .A1(n466), .A2(n529), .ZN(n467) );
  NAND2_X1 U530 ( .A1(n467), .A2(n546), .ZN(n534) );
  NOR2_X1 U531 ( .A1(n534), .A2(n525), .ZN(n468) );
  NOR2_X1 U532 ( .A1(n469), .A2(n468), .ZN(n485) );
  NOR2_X1 U533 ( .A1(n576), .A2(n485), .ZN(n470) );
  NAND2_X1 U534 ( .A1(n579), .A2(n470), .ZN(n473) );
  NAND2_X1 U535 ( .A1(n559), .A2(n474), .ZN(n488) );
  NOR2_X1 U536 ( .A1(n521), .A2(n488), .ZN(n476) );
  XNOR2_X1 U537 ( .A(KEYINPUT38), .B(KEYINPUT105), .ZN(n475) );
  XNOR2_X1 U538 ( .A(n476), .B(n475), .ZN(n477) );
  NAND2_X1 U539 ( .A1(n506), .A2(n525), .ZN(n480) );
  XOR2_X1 U540 ( .A(KEYINPUT40), .B(KEYINPUT109), .Z(n478) );
  NAND2_X1 U541 ( .A1(n557), .A2(n561), .ZN(n482) );
  NAND2_X1 U542 ( .A1(n483), .A2(n576), .ZN(n484) );
  XOR2_X1 U543 ( .A(KEYINPUT16), .B(n484), .Z(n487) );
  INV_X1 U544 ( .A(n485), .ZN(n486) );
  NAND2_X1 U545 ( .A1(n487), .A2(n486), .ZN(n511) );
  NOR2_X1 U546 ( .A1(n488), .A2(n511), .ZN(n498) );
  NAND2_X1 U547 ( .A1(n546), .A2(n498), .ZN(n491) );
  XOR2_X1 U548 ( .A(G1GAT), .B(KEYINPUT34), .Z(n489) );
  XNOR2_X1 U549 ( .A(KEYINPUT99), .B(n489), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(G1324GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n493) );
  NAND2_X1 U552 ( .A1(n498), .A2(n523), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U554 ( .A(G8GAT), .B(n494), .ZN(G1325GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n496) );
  NAND2_X1 U556 ( .A1(n498), .A2(n525), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U558 ( .A(G15GAT), .B(n497), .ZN(G1326GAT) );
  XOR2_X1 U559 ( .A(G22GAT), .B(KEYINPUT103), .Z(n500) );
  NAND2_X1 U560 ( .A1(n498), .A2(n529), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(G1327GAT) );
  NAND2_X1 U562 ( .A1(n546), .A2(n506), .ZN(n503) );
  XNOR2_X1 U563 ( .A(G29GAT), .B(KEYINPUT107), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n501), .B(KEYINPUT39), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  XNOR2_X1 U566 ( .A(G36GAT), .B(KEYINPUT108), .ZN(n505) );
  NAND2_X1 U567 ( .A1(n523), .A2(n506), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(G1329GAT) );
  NAND2_X1 U569 ( .A1(n529), .A2(n506), .ZN(n507) );
  XNOR2_X1 U570 ( .A(n507), .B(KEYINPUT110), .ZN(n508) );
  XNOR2_X1 U571 ( .A(G50GAT), .B(n508), .ZN(G1331GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT42), .B(KEYINPUT111), .Z(n513) );
  NAND2_X1 U573 ( .A1(n510), .A2(n509), .ZN(n520) );
  NOR2_X1 U574 ( .A1(n520), .A2(n511), .ZN(n517) );
  NAND2_X1 U575 ( .A1(n517), .A2(n546), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(n514), .ZN(G1332GAT) );
  NAND2_X1 U578 ( .A1(n517), .A2(n523), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n515), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U580 ( .A1(n517), .A2(n525), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n516), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U583 ( .A1(n517), .A2(n529), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NOR2_X1 U585 ( .A1(n521), .A2(n520), .ZN(n528) );
  NAND2_X1 U586 ( .A1(n528), .A2(n546), .ZN(n522) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(n522), .ZN(G1336GAT) );
  NAND2_X1 U588 ( .A1(n528), .A2(n523), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U590 ( .A1(n528), .A2(n525), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n526), .B(KEYINPUT112), .ZN(n527) );
  XNOR2_X1 U592 ( .A(G99GAT), .B(n527), .ZN(G1338GAT) );
  NAND2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(KEYINPUT44), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  OR2_X1 U596 ( .A1(n532), .A2(n549), .ZN(n533) );
  NOR2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n559), .A2(n541), .ZN(n535) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U601 ( .A1(n541), .A2(n509), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n539) );
  NAND2_X1 U604 ( .A1(n541), .A2(n576), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U608 ( .A1(n541), .A2(n557), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n545) );
  XOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT118), .Z(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  NAND2_X1 U612 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n556) );
  NAND2_X1 U614 ( .A1(n556), .A2(n568), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n550), .B(KEYINPUT120), .ZN(n551) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(n551), .ZN(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n553) );
  NAND2_X1 U618 ( .A1(n556), .A2(n509), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(n554), .ZN(G1345GAT) );
  NAND2_X1 U621 ( .A1(n556), .A2(n576), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U625 ( .A1(n559), .A2(n561), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G169GAT), .B(n560), .ZN(G1348GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n509), .ZN(n563) );
  XOR2_X1 U628 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(n564), .ZN(G1349GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT59), .B(KEYINPUT60), .Z(n570) );
  INV_X1 U632 ( .A(n565), .ZN(n566) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n580) );
  NAND2_X1 U634 ( .A1(n580), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n572) );
  XOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT123), .Z(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT61), .Z(n575) );
  NAND2_X1 U639 ( .A1(n580), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  NAND2_X1 U641 ( .A1(n580), .A2(n576), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(KEYINPUT124), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G211GAT), .B(n578), .ZN(G1354GAT) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(KEYINPUT125), .ZN(n584) );
  XOR2_X1 U645 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n582) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(G1355GAT) );
endmodule

