//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 0 0 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n807,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT3), .ZN(new_n203));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT22), .ZN(new_n205));
  INV_X1    g004(.A(G211gat), .ZN(new_n206));
  INV_X1    g005(.A(G218gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n204), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G211gat), .B(G218gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n212), .A2(KEYINPUT75), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n204), .A3(new_n208), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(KEYINPUT75), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n203), .B1(new_n216), .B2(KEYINPUT29), .ZN(new_n217));
  INV_X1    g016(.A(G141gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT82), .B1(new_n218), .B2(G148gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT82), .ZN(new_n220));
  INV_X1    g019(.A(G148gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(new_n221), .A3(G141gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n218), .A2(G148gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n219), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(G155gat), .A2(G162gat), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(KEYINPUT83), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT83), .ZN(new_n229));
  INV_X1    g028(.A(new_n227), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n229), .B1(new_n230), .B2(new_n225), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n227), .A2(KEYINPUT2), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n224), .A2(new_n228), .A3(new_n231), .A4(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT2), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n218), .A2(G148gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n221), .A2(G141gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT81), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n225), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT81), .B1(G155gat), .B2(G162gat), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n240), .A2(new_n227), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n237), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n233), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n202), .B1(new_n217), .B2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT85), .B(KEYINPUT3), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n233), .A2(new_n242), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT29), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(KEYINPUT90), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(KEYINPUT90), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n216), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n244), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT91), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n233), .A2(new_n242), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n212), .A2(new_n214), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT89), .B1(new_n256), .B2(new_n248), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n257), .A2(new_n245), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n256), .A2(KEYINPUT89), .A3(new_n248), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n255), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n216), .A2(new_n249), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n202), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n253), .A2(new_n254), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n254), .B1(new_n253), .B2(new_n262), .ZN(new_n265));
  OAI21_X1  g064(.A(G50gat), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n265), .ZN(new_n267));
  INV_X1    g066(.A(G50gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n267), .A2(new_n268), .A3(new_n263), .ZN(new_n269));
  XOR2_X1   g068(.A(G78gat), .B(G106gat), .Z(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(G22gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT31), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n266), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n272), .B1(new_n266), .B2(new_n269), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G227gat), .A2(G233gat), .ZN(new_n276));
  XOR2_X1   g075(.A(new_n276), .B(KEYINPUT64), .Z(new_n277));
  XOR2_X1   g076(.A(G127gat), .B(G134gat), .Z(new_n278));
  XNOR2_X1  g077(.A(G113gat), .B(G120gat), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n278), .B1(KEYINPUT1), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G120gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G113gat), .ZN(new_n282));
  INV_X1    g081(.A(G113gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G120gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G127gat), .B(G134gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT1), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n280), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n280), .A2(KEYINPUT72), .A3(new_n288), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT23), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n294), .A2(G176gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT65), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(G169gat), .ZN(new_n297));
  INV_X1    g096(.A(G169gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(KEYINPUT65), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n295), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(G183gat), .A2(G190gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT24), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n305));
  INV_X1    g104(.A(G183gat), .ZN(new_n306));
  INV_X1    g105(.A(G190gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n304), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  OR2_X1    g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310));
  AND2_X1   g109(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n311));
  NOR2_X1   g110(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n300), .A2(new_n301), .A3(new_n309), .A4(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT25), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT67), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n302), .A2(new_n317), .A3(new_n303), .ZN(new_n318));
  OAI211_X1 g117(.A(G183gat), .B(G190gat), .C1(KEYINPUT67), .C2(KEYINPUT24), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(new_n308), .A3(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT23), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n315), .B1(G169gat), .B2(G176gat), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n320), .A2(new_n313), .A3(new_n322), .A4(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n316), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT68), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n313), .A2(new_n322), .A3(new_n323), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n314), .A2(new_n315), .B1(new_n328), .B2(new_n320), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT68), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT27), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT69), .B1(new_n332), .B2(G183gat), .ZN(new_n333));
  AOI21_X1  g132(.A(G190gat), .B1(new_n332), .B2(G183gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT69), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(new_n306), .A3(KEYINPUT27), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n333), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT28), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT70), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT70), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n337), .A2(new_n341), .A3(new_n338), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n307), .B1(new_n306), .B2(KEYINPUT27), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n332), .A2(G183gat), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n343), .A2(new_n344), .A3(new_n338), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n340), .A2(new_n342), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT71), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT26), .B1(new_n310), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT26), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n321), .A2(KEYINPUT71), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n351), .A3(new_n301), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(new_n302), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n347), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n293), .B1(new_n331), .B2(new_n355), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n316), .A2(KEYINPUT68), .A3(new_n324), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT68), .B1(new_n316), .B2(new_n324), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n293), .B(new_n355), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n277), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT33), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT73), .B(G71gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n364), .B(G99gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(G15gat), .B(G43gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n355), .B1(new_n357), .B2(new_n358), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(new_n292), .A3(new_n291), .ZN(new_n370));
  INV_X1    g169(.A(new_n277), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(new_n371), .A3(new_n359), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n361), .A2(KEYINPUT32), .A3(new_n372), .ZN(new_n373));
  XOR2_X1   g172(.A(KEYINPUT74), .B(KEYINPUT34), .Z(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT32), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n370), .A2(new_n376), .A3(new_n371), .A4(new_n359), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n373), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n375), .B1(new_n373), .B2(new_n377), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n368), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n373), .A2(new_n377), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n374), .ZN(new_n383));
  INV_X1    g182(.A(new_n368), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n384), .A3(new_n378), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n275), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT35), .ZN(new_n389));
  NAND2_X1  g188(.A1(G226gat), .A2(G233gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT76), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n392), .B1(new_n355), .B2(new_n325), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n345), .B1(new_n339), .B2(KEYINPUT70), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n353), .B1(new_n394), .B2(new_n342), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n395), .A2(KEYINPUT76), .A3(new_n329), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n391), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n391), .A2(KEYINPUT29), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n369), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n397), .A2(new_n216), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT77), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n397), .A2(KEYINPUT77), .A3(new_n216), .A4(new_n399), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n355), .A2(new_n392), .A3(new_n325), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT76), .B1(new_n395), .B2(new_n329), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n405), .A3(new_n398), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n391), .B(new_n355), .C1(new_n357), .C2(new_n358), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n216), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G8gat), .B(G36gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(G64gat), .B(G92gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n402), .A2(new_n403), .A3(new_n409), .A4(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT80), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT30), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n408), .B1(new_n400), .B2(new_n401), .ZN(new_n419));
  INV_X1    g218(.A(new_n417), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n419), .A2(new_n403), .A3(new_n413), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n415), .A2(new_n416), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AND4_X1   g223(.A1(KEYINPUT78), .A2(new_n402), .A3(new_n403), .A4(new_n409), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT78), .B1(new_n419), .B2(new_n403), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n412), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT79), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n402), .A2(new_n403), .A3(new_n409), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT78), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n419), .A2(KEYINPUT78), .A3(new_n403), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT79), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n434), .A3(new_n412), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n424), .B1(new_n428), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT94), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT84), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n286), .B1(new_n287), .B2(new_n285), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n280), .A2(KEYINPUT84), .A3(new_n288), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n247), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n203), .B1(new_n233), .B2(new_n242), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT86), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n280), .A2(KEYINPUT84), .A3(new_n288), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT84), .B1(new_n280), .B2(new_n288), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n444), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT86), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n448), .A2(new_n449), .A3(new_n450), .A4(new_n247), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n445), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT4), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n243), .A2(new_n289), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n293), .A2(new_n255), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n454), .B1(new_n455), .B2(new_n453), .ZN(new_n456));
  NAND2_X1  g255(.A1(G225gat), .A2(G233gat), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n458), .A2(KEYINPUT5), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n452), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(G1gat), .B(G29gat), .ZN(new_n461));
  INV_X1    g260(.A(G85gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT0), .B(G57gat), .ZN(new_n464));
  XOR2_X1   g263(.A(new_n463), .B(new_n464), .Z(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n292), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT72), .B1(new_n280), .B2(new_n288), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n255), .B(KEYINPUT4), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n453), .B1(new_n243), .B2(new_n289), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(new_n470), .A3(new_n457), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n471), .B1(new_n445), .B2(new_n451), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n243), .A2(new_n289), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n473), .B1(new_n448), .B2(new_n243), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT5), .B1(new_n474), .B2(new_n457), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n460), .B(new_n466), .C1(new_n472), .C2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n475), .ZN(new_n479));
  INV_X1    g278(.A(new_n471), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n452), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n466), .B1(new_n482), .B2(new_n460), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n437), .B1(new_n478), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n475), .B1(new_n452), .B2(new_n480), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n452), .A2(new_n456), .A3(new_n459), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n465), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT88), .B1(new_n487), .B2(new_n477), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n487), .A2(KEYINPUT94), .A3(new_n477), .A4(new_n476), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT88), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n483), .A2(new_n490), .A3(KEYINPUT6), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n484), .A2(new_n488), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n388), .A2(new_n389), .A3(new_n436), .A4(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT87), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n483), .B1(new_n478), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n495), .B1(new_n494), .B2(new_n478), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n488), .A2(new_n491), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n418), .A2(new_n421), .B1(new_n415), .B2(new_n416), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n434), .B1(new_n433), .B2(new_n412), .ZN(new_n500));
  AOI211_X1 g299(.A(KEYINPUT79), .B(new_n413), .C1(new_n431), .C2(new_n432), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n498), .B(new_n499), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT35), .B1(new_n502), .B2(new_n387), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n493), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT36), .ZN(new_n505));
  NOR3_X1   g304(.A1(new_n379), .A2(new_n380), .A3(new_n368), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n384), .B1(new_n383), .B2(new_n378), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n381), .A2(new_n385), .A3(KEYINPUT36), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n275), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n510), .B1(new_n502), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT38), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n414), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT37), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n515), .B1(new_n431), .B2(new_n432), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n419), .A2(new_n515), .A3(new_n403), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n412), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n514), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n406), .A2(new_n216), .A3(new_n407), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT95), .ZN(new_n521));
  INV_X1    g320(.A(new_n216), .ZN(new_n522));
  INV_X1    g321(.A(new_n399), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n390), .B1(new_n404), .B2(new_n405), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT95), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n406), .A2(new_n526), .A3(new_n216), .A4(new_n407), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n521), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT37), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n413), .A2(KEYINPUT38), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n529), .A2(new_n517), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n492), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n519), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n452), .A2(new_n456), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n458), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT39), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n536), .B1(new_n474), .B2(new_n457), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n534), .A2(new_n536), .A3(new_n458), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n539), .A2(KEYINPUT92), .A3(new_n466), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT92), .B1(new_n539), .B2(new_n466), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(KEYINPUT93), .A2(KEYINPUT40), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n543), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n487), .A3(new_n545), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n533), .B(new_n275), .C1(new_n436), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n512), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n504), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G29gat), .A2(G36gat), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NOR3_X1   g351(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(G43gat), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT97), .B1(new_n555), .B2(G50gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT97), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(new_n268), .A3(G43gat), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n556), .B(new_n558), .C1(G43gat), .C2(new_n268), .ZN(new_n559));
  XOR2_X1   g358(.A(KEYINPUT96), .B(KEYINPUT15), .Z(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n268), .A2(G43gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n555), .A2(G50gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT15), .ZN(new_n564));
  OR3_X1    g363(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n554), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n565), .A2(new_n554), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT98), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT98), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n565), .A2(new_n554), .ZN(new_n570));
  NOR3_X1   g369(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n571), .B1(new_n559), .B2(new_n560), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n569), .B(new_n570), .C1(new_n572), .C2(new_n554), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT17), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G15gat), .B(G22gat), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT16), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n577), .B1(new_n578), .B2(G1gat), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n579), .B1(G1gat), .B2(new_n577), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n580), .A2(G8gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(G8gat), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT17), .B1(new_n566), .B2(new_n567), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n576), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G229gat), .A2(G233gat), .ZN(new_n587));
  AOI21_X1  g386(.A(KEYINPUT99), .B1(new_n574), .B2(new_n583), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n574), .A2(new_n583), .A3(KEYINPUT99), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n586), .B(new_n587), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT18), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n588), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n574), .A2(new_n583), .A3(KEYINPUT99), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n595), .A2(KEYINPUT18), .A3(new_n587), .A4(new_n586), .ZN(new_n596));
  OAI22_X1  g395(.A1(new_n589), .A2(new_n588), .B1(new_n574), .B2(new_n583), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n587), .B(KEYINPUT13), .Z(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n592), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G113gat), .B(G141gat), .ZN(new_n601));
  INV_X1    g400(.A(G197gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT11), .B(G169gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT12), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT100), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n592), .A2(new_n596), .A3(new_n599), .A4(new_n606), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n609), .B1(new_n608), .B2(new_n610), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(G64gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(G57gat), .ZN(new_n616));
  XOR2_X1   g415(.A(KEYINPUT102), .B(G57gat), .Z(new_n617));
  OAI21_X1  g416(.A(new_n616), .B1(new_n617), .B2(new_n615), .ZN(new_n618));
  NOR2_X1   g417(.A1(G71gat), .A2(G78gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(KEYINPUT9), .ZN(new_n620));
  NAND2_X1  g419(.A1(G71gat), .A2(G78gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT101), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n621), .B1(new_n619), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n625), .B1(new_n624), .B2(new_n619), .ZN(new_n626));
  INV_X1    g425(.A(new_n616), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n615), .A2(G57gat), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT9), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n623), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT103), .B(KEYINPUT21), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(G127gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(G155gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(new_n306), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G211gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n637), .B(new_n640), .ZN(new_n641));
  AOI22_X1  g440(.A1(new_n618), .A2(new_n622), .B1(new_n626), .B2(new_n629), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n583), .B1(KEYINPUT21), .B2(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n641), .A2(new_n645), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G99gat), .A2(G106gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT8), .ZN(new_n650));
  NAND2_X1  g449(.A1(G85gat), .A2(G92gat), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT7), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(G92gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n462), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n650), .A2(new_n653), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT104), .ZN(new_n658));
  AOI22_X1  g457(.A1(KEYINPUT8), .A2(new_n649), .B1(new_n462), .B2(new_n654), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n659), .A2(new_n660), .A3(new_n653), .A4(new_n656), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(G99gat), .B(G106gat), .Z(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n658), .A2(new_n663), .A3(new_n661), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(KEYINPUT105), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n668));
  INV_X1    g467(.A(new_n666), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n663), .B1(new_n658), .B2(new_n661), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n576), .A2(new_n585), .A3(new_n667), .A4(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n667), .ZN(new_n673));
  AND2_X1   g472(.A1(G232gat), .A2(G233gat), .ZN(new_n674));
  AOI22_X1  g473(.A1(new_n673), .A2(new_n574), .B1(KEYINPUT41), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g475(.A(G134gat), .B(G162gat), .Z(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n676), .B(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n674), .A2(KEYINPUT41), .ZN(new_n680));
  XNOR2_X1  g479(.A(G190gat), .B(G218gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n679), .A2(new_n682), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n648), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(G230gat), .A2(G233gat), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n631), .B1(new_n669), .B2(new_n670), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n665), .A2(new_n642), .A3(new_n666), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT10), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n642), .A2(KEYINPUT10), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n691), .B1(new_n671), .B2(new_n667), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n687), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n687), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n688), .A2(new_n689), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(G120gat), .B(G148gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(G176gat), .B(G204gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n693), .A2(new_n695), .A3(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n693), .A2(new_n702), .ZN(new_n703));
  OAI211_X1 g502(.A(KEYINPUT106), .B(new_n687), .C1(new_n690), .C2(new_n692), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(new_n695), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n701), .B1(new_n705), .B2(new_n698), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n614), .A2(new_n686), .A3(new_n707), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n549), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n498), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G1gat), .ZN(G1324gat));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n713));
  INV_X1    g512(.A(new_n436), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g514(.A(KEYINPUT16), .B(G8gat), .Z(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT42), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n713), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n715), .A2(KEYINPUT108), .A3(KEYINPUT42), .A4(new_n716), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n709), .ZN(new_n722));
  OAI21_X1  g521(.A(G8gat), .B1(new_n722), .B2(new_n436), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT107), .B1(new_n717), .B2(new_n718), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n717), .A2(KEYINPUT107), .A3(new_n718), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n721), .B(new_n723), .C1(new_n724), .C2(new_n725), .ZN(G1325gat));
  AOI21_X1  g525(.A(G15gat), .B1(new_n709), .B2(new_n386), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n510), .A2(G15gat), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n727), .B1(new_n709), .B2(new_n728), .ZN(G1326gat));
  NAND2_X1  g528(.A1(new_n709), .A2(new_n511), .ZN(new_n730));
  XNOR2_X1  g529(.A(KEYINPUT43), .B(G22gat), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1327gat));
  AOI21_X1  g531(.A(new_n685), .B1(new_n504), .B2(new_n548), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n614), .A2(new_n648), .A3(new_n707), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n735), .A2(G29gat), .A3(new_n498), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n736), .B(KEYINPUT45), .Z(new_n737));
  AND3_X1   g536(.A1(new_n512), .A2(KEYINPUT110), .A3(new_n547), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT110), .B1(new_n512), .B2(new_n547), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n504), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n685), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI211_X1 g543(.A(new_n743), .B(new_n685), .C1(new_n504), .C2(new_n548), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n648), .B(KEYINPUT109), .Z(new_n747));
  NAND2_X1  g546(.A1(new_n608), .A2(new_n610), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n747), .A2(new_n748), .A3(new_n706), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n744), .A2(new_n710), .A3(new_n746), .A4(new_n750), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n751), .A2(KEYINPUT111), .ZN(new_n752));
  OAI21_X1  g551(.A(G29gat), .B1(new_n751), .B2(KEYINPUT111), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n737), .B1(new_n752), .B2(new_n753), .ZN(G1328gat));
  NOR3_X1   g553(.A1(new_n735), .A2(G36gat), .A3(new_n436), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT46), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n744), .A2(new_n714), .A3(new_n746), .A4(new_n750), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(G36gat), .B1(new_n757), .B2(new_n758), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n756), .B1(new_n759), .B2(new_n760), .ZN(G1329gat));
  NAND4_X1  g560(.A1(new_n733), .A2(new_n555), .A3(new_n386), .A4(new_n734), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT44), .B1(new_n740), .B2(new_n741), .ZN(new_n763));
  INV_X1    g562(.A(new_n510), .ZN(new_n764));
  NOR4_X1   g563(.A1(new_n763), .A2(new_n764), .A3(new_n745), .A4(new_n749), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n762), .B1(new_n765), .B2(new_n555), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g567(.A(KEYINPUT47), .B(new_n762), .C1(new_n765), .C2(new_n555), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(G1330gat));
  NOR2_X1   g569(.A1(new_n275), .A2(G50gat), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n733), .A2(new_n734), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT48), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI211_X1 g575(.A(KEYINPUT114), .B(KEYINPUT48), .C1(new_n772), .C2(new_n773), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR4_X1   g577(.A1(new_n763), .A2(new_n275), .A3(new_n745), .A4(new_n749), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n772), .B1(new_n779), .B2(new_n268), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n744), .A2(new_n746), .A3(new_n750), .ZN(new_n782));
  OAI21_X1  g581(.A(G50gat), .B1(new_n782), .B2(new_n275), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n776), .A2(new_n777), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(new_n784), .A3(new_n772), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n781), .A2(new_n785), .ZN(G1331gat));
  NOR3_X1   g585(.A1(new_n686), .A2(new_n748), .A3(new_n706), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n740), .A2(new_n787), .ZN(new_n788));
  OR3_X1    g587(.A1(new_n788), .A2(KEYINPUT115), .A3(new_n498), .ZN(new_n789));
  OAI21_X1  g588(.A(KEYINPUT115), .B1(new_n788), .B2(new_n498), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(new_n617), .ZN(G1332gat));
  INV_X1    g591(.A(new_n788), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n436), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT116), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n793), .A2(new_n797), .A3(new_n794), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n799), .B(new_n800), .ZN(G1333gat));
  OAI21_X1  g600(.A(G71gat), .B1(new_n788), .B2(new_n764), .ZN(new_n802));
  INV_X1    g601(.A(G71gat), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n386), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n788), .B2(new_n804), .ZN(new_n805));
  XOR2_X1   g604(.A(new_n805), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g605(.A1(new_n788), .A2(new_n275), .ZN(new_n807));
  XOR2_X1   g606(.A(KEYINPUT117), .B(G78gat), .Z(new_n808));
  XNOR2_X1  g607(.A(new_n807), .B(new_n808), .ZN(G1335gat));
  INV_X1    g608(.A(new_n648), .ZN(new_n810));
  INV_X1    g609(.A(new_n748), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT118), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n740), .A2(new_n741), .A3(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n740), .A2(KEYINPUT51), .A3(new_n741), .A4(new_n813), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n818), .A2(new_n710), .A3(new_n707), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n813), .A2(new_n707), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n763), .A2(new_n745), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n498), .A2(new_n462), .ZN(new_n822));
  AOI22_X1  g621(.A1(new_n819), .A2(new_n462), .B1(new_n821), .B2(new_n822), .ZN(G1336gat));
  INV_X1    g622(.A(new_n820), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n744), .A2(new_n714), .A3(new_n746), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(G92gat), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n436), .A2(G92gat), .A3(new_n706), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n818), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n826), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  XOR2_X1   g629(.A(new_n827), .B(KEYINPUT119), .Z(new_n831));
  AOI22_X1  g630(.A1(G92gat), .A2(new_n825), .B1(new_n818), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n830), .B1(new_n832), .B2(new_n829), .ZN(G1337gat));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n386), .A3(new_n707), .ZN(new_n834));
  INV_X1    g633(.A(G99gat), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n764), .A2(new_n835), .ZN(new_n836));
  AOI22_X1  g635(.A1(new_n834), .A2(new_n835), .B1(new_n821), .B2(new_n836), .ZN(G1338gat));
  INV_X1    g636(.A(G106gat), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n838), .B1(new_n821), .B2(new_n511), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n275), .A2(G106gat), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  AOI211_X1 g640(.A(new_n706), .B(new_n841), .C1(new_n816), .C2(new_n817), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT53), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n744), .A2(new_n746), .A3(new_n824), .ZN(new_n844));
  OAI21_X1  g643(.A(G106gat), .B1(new_n844), .B2(new_n275), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n818), .A2(new_n707), .A3(new_n840), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n843), .A2(new_n848), .ZN(G1339gat));
  NAND2_X1  g648(.A1(new_n436), .A2(new_n710), .ZN(new_n850));
  OR3_X1    g649(.A1(new_n690), .A2(new_n692), .A3(new_n687), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n693), .A3(KEYINPUT54), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n703), .A2(new_n704), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT120), .B1(new_n855), .B2(new_n698), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT54), .B1(new_n703), .B2(new_n704), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n857), .A2(new_n858), .A3(new_n699), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n852), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT55), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n701), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n852), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n855), .A2(KEYINPUT120), .A3(new_n698), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n858), .B1(new_n857), .B2(new_n699), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT55), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n862), .A2(new_n748), .A3(new_n867), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n597), .A2(new_n598), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n587), .B1(new_n595), .B2(new_n586), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n605), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n872), .A2(new_n610), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n707), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n741), .B1(new_n868), .B2(new_n874), .ZN(new_n875));
  AND4_X1   g674(.A1(new_n741), .A2(new_n862), .A3(new_n867), .A4(new_n873), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n747), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n686), .A2(new_n707), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n811), .ZN(new_n879));
  AOI211_X1 g678(.A(new_n387), .B(new_n850), .C1(new_n877), .C2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n283), .A3(new_n748), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n880), .A2(new_n613), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(new_n283), .ZN(G1340gat));
  NAND2_X1  g682(.A1(new_n880), .A2(new_n707), .ZN(new_n884));
  XOR2_X1   g683(.A(KEYINPUT121), .B(G120gat), .Z(new_n885));
  XNOR2_X1  g684(.A(new_n884), .B(new_n885), .ZN(G1341gat));
  AOI21_X1  g685(.A(G127gat), .B1(new_n880), .B2(new_n648), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n747), .A2(new_n634), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n880), .B2(new_n888), .ZN(G1342gat));
  NAND2_X1  g688(.A1(new_n880), .A2(new_n741), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(G134gat), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n893), .B1(KEYINPUT56), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n895), .B1(KEYINPUT56), .B2(new_n894), .ZN(G1343gat));
  NOR2_X1   g695(.A1(new_n850), .A2(new_n510), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n275), .B1(new_n877), .B2(new_n879), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n700), .B1(new_n866), .B2(KEYINPUT55), .ZN(new_n902));
  AOI211_X1 g701(.A(new_n861), .B(new_n863), .C1(new_n864), .C2(new_n865), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n741), .A3(new_n873), .ZN(new_n905));
  INV_X1    g704(.A(new_n874), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n906), .B1(new_n904), .B2(new_n613), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n905), .B1(new_n907), .B2(new_n741), .ZN(new_n908));
  AOI22_X1  g707(.A1(new_n908), .A2(new_n810), .B1(new_n811), .B2(new_n878), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT57), .B1(new_n909), .B2(new_n275), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n901), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(G141gat), .B1(new_n911), .B2(new_n614), .ZN(new_n912));
  INV_X1    g711(.A(new_n899), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n913), .A2(new_n898), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n614), .A2(G141gat), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT58), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(new_n911), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n748), .ZN(new_n919));
  AOI22_X1  g718(.A1(new_n919), .A2(G141gat), .B1(new_n914), .B2(new_n915), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT58), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(G1344gat));
  NAND3_X1  g721(.A1(new_n914), .A2(new_n221), .A3(new_n707), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n275), .A2(KEYINPUT57), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n613), .A2(new_n862), .A3(new_n867), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n741), .B1(new_n926), .B2(new_n874), .ZN(new_n927));
  OAI21_X1  g726(.A(KEYINPUT122), .B1(new_n927), .B2(new_n876), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n929), .B(new_n905), .C1(new_n907), .C2(new_n741), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n928), .A2(new_n930), .A3(new_n810), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n878), .A2(new_n614), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n925), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n877), .A2(new_n879), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n900), .B1(new_n934), .B2(new_n511), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n897), .A2(new_n707), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n933), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  OAI211_X1 g736(.A(KEYINPUT123), .B(KEYINPUT59), .C1(new_n937), .C2(new_n221), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n221), .A2(KEYINPUT59), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n939), .B1(new_n911), .B2(new_n706), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n931), .A2(new_n932), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n924), .ZN(new_n943));
  INV_X1    g742(.A(new_n935), .ZN(new_n944));
  INV_X1    g743(.A(new_n936), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G148gat), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT123), .B1(new_n947), .B2(KEYINPUT59), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n923), .B1(new_n941), .B2(new_n948), .ZN(G1345gat));
  AOI21_X1  g748(.A(G155gat), .B1(new_n914), .B2(new_n648), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n747), .A2(new_n636), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(new_n918), .B2(new_n951), .ZN(G1346gat));
  OAI21_X1  g751(.A(G162gat), .B1(new_n911), .B2(new_n685), .ZN(new_n953));
  INV_X1    g752(.A(G162gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n914), .A2(new_n954), .A3(new_n741), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(new_n955), .ZN(G1347gat));
  NOR3_X1   g755(.A1(new_n436), .A2(new_n387), .A3(new_n710), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n934), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(G169gat), .B1(new_n958), .B2(new_n614), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT124), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n748), .B1(new_n297), .B2(new_n299), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n960), .B1(new_n958), .B2(new_n961), .ZN(G1348gat));
  INV_X1    g761(.A(new_n958), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(new_n707), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(G176gat), .ZN(G1349gat));
  OAI21_X1  g764(.A(G183gat), .B1(new_n958), .B2(new_n747), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n306), .A2(KEYINPUT27), .ZN(new_n967));
  OR3_X1    g766(.A1(new_n810), .A2(new_n344), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n966), .B1(new_n958), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g769(.A(new_n957), .ZN(new_n971));
  AOI211_X1 g770(.A(new_n685), .B(new_n971), .C1(new_n877), .C2(new_n879), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(new_n307), .ZN(new_n973));
  OAI211_X1 g772(.A(KEYINPUT125), .B(KEYINPUT61), .C1(new_n972), .C2(new_n307), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT61), .ZN(new_n975));
  OAI211_X1 g774(.A(new_n975), .B(G190gat), .C1(new_n958), .C2(new_n685), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(G190gat), .B1(new_n958), .B2(new_n685), .ZN(new_n978));
  AOI21_X1  g777(.A(KEYINPUT125), .B1(new_n978), .B2(KEYINPUT61), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n973), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(KEYINPUT126), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n982));
  OAI211_X1 g781(.A(new_n982), .B(new_n973), .C1(new_n977), .C2(new_n979), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n981), .A2(new_n983), .ZN(G1351gat));
  NOR3_X1   g783(.A1(new_n510), .A2(new_n436), .A3(new_n710), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n899), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n986), .A2(new_n602), .A3(new_n748), .ZN(new_n987));
  AND3_X1   g786(.A1(new_n943), .A2(new_n944), .A3(new_n985), .ZN(new_n988));
  AND2_X1   g787(.A1(new_n988), .A2(new_n613), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n987), .B1(new_n989), .B2(new_n602), .ZN(G1352gat));
  INV_X1    g789(.A(G204gat), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n986), .A2(new_n991), .A3(new_n707), .ZN(new_n992));
  XOR2_X1   g791(.A(new_n992), .B(KEYINPUT62), .Z(new_n993));
  NAND4_X1  g792(.A1(new_n943), .A2(new_n944), .A3(new_n707), .A4(new_n985), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n995));
  AND2_X1   g794(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g795(.A(G204gat), .B1(new_n994), .B2(new_n995), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n993), .B1(new_n996), .B2(new_n997), .ZN(G1353gat));
  NAND3_X1  g797(.A1(new_n986), .A2(new_n206), .A3(new_n648), .ZN(new_n999));
  NAND4_X1  g798(.A1(new_n943), .A2(new_n944), .A3(new_n648), .A4(new_n985), .ZN(new_n1000));
  AND3_X1   g799(.A1(new_n1000), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1001));
  AOI21_X1  g800(.A(KEYINPUT63), .B1(new_n1000), .B2(G211gat), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n999), .B1(new_n1001), .B2(new_n1002), .ZN(G1354gat));
  AOI21_X1  g802(.A(G218gat), .B1(new_n986), .B2(new_n741), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n685), .A2(new_n207), .ZN(new_n1005));
  AOI21_X1  g804(.A(new_n1004), .B1(new_n988), .B2(new_n1005), .ZN(G1355gat));
endmodule


