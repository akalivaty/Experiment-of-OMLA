//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n562, new_n563, new_n564,
    new_n565, new_n567, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n467));
  AND3_X1   g042(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n467), .B1(new_n464), .B2(new_n466), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n463), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT65), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n462), .B1(new_n472), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G137), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n480), .B1(new_n474), .B2(new_n476), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n483), .A2(new_n459), .A3(KEYINPUT3), .ZN(new_n484));
  AOI21_X1  g059(.A(KEYINPUT67), .B1(new_n465), .B2(G2104), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n465), .A2(G2104), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(KEYINPUT68), .B1(new_n482), .B2(new_n487), .ZN(new_n488));
  NOR3_X1   g063(.A1(new_n465), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n483), .B1(new_n459), .B2(KEYINPUT3), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(new_n464), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n491), .A2(new_n492), .A3(new_n481), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n479), .A2(new_n494), .ZN(G160));
  OAI221_X1 g070(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n477), .C2(G112), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n491), .A2(new_n473), .ZN(new_n497));
  INV_X1    g072(.A(G136), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n487), .A2(new_n477), .ZN(new_n500));
  XNOR2_X1  g075(.A(new_n500), .B(KEYINPUT69), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n499), .B1(new_n501), .B2(G124), .ZN(G162));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(new_n473), .B2(G114), .ZN(new_n504));
  NOR2_X1   g079(.A1(G102), .A2(G2105), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(G126), .A2(G2105), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G138), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n510), .B1(new_n474), .B2(new_n476), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n509), .B1(new_n511), .B2(KEYINPUT4), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n507), .B1(new_n512), .B2(new_n487), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT66), .B1(new_n486), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(KEYINPUT4), .B1(new_n517), .B2(new_n511), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n503), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n511), .B1(new_n468), .B2(new_n469), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT4), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI211_X1 g097(.A(new_n521), .B(new_n510), .C1(new_n474), .C2(new_n476), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n491), .B1(new_n523), .B2(new_n509), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n522), .A2(KEYINPUT70), .A3(new_n524), .A4(new_n507), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n519), .A2(new_n525), .ZN(G164));
  NAND2_X1  g101(.A1(G75), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT5), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT5), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G543), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G62), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n527), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G651), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n529), .A2(new_n531), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT6), .B(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G88), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G50), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n539), .A2(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n536), .A2(new_n543), .ZN(G166));
  AND2_X1   g119(.A1(new_n537), .A2(new_n538), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G89), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n538), .A2(G543), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G51), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n537), .A2(G63), .A3(G651), .ZN(new_n549));
  NAND3_X1  g124(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT7), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n546), .A2(new_n548), .A3(new_n549), .A4(new_n551), .ZN(G286));
  INV_X1    g127(.A(G286), .ZN(G168));
  AOI22_X1  g128(.A1(new_n537), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G651), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT71), .Z(new_n557));
  AND2_X1   g132(.A1(new_n545), .A2(G90), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n547), .A2(G52), .ZN(new_n559));
  OR3_X1    g134(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(G301));
  INV_X1    g135(.A(G301), .ZN(G171));
  AOI22_X1  g136(.A1(new_n537), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n562));
  OR2_X1    g137(.A1(new_n562), .A2(new_n555), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n545), .A2(G81), .B1(G43), .B2(new_n547), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  AND3_X1   g141(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G36), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(G188));
  NAND2_X1  g146(.A1(new_n547), .A2(G53), .ZN(new_n572));
  XOR2_X1   g147(.A(new_n572), .B(KEYINPUT9), .Z(new_n573));
  NAND3_X1  g148(.A1(new_n545), .A2(KEYINPUT72), .A3(G91), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT72), .ZN(new_n575));
  INV_X1    g150(.A(G91), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n539), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n537), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n574), .B(new_n577), .C1(new_n555), .C2(new_n578), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G299));
  INV_X1    g156(.A(G166), .ZN(G303));
  NAND2_X1  g157(.A1(new_n545), .A2(G87), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n547), .A2(G49), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n537), .B2(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G288));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n532), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G651), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(KEYINPUT73), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT73), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n589), .A2(new_n592), .A3(G651), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n547), .A2(G48), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n545), .A2(G86), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G305));
  AOI22_X1  g172(.A1(new_n537), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n555), .ZN(new_n599));
  INV_X1    g174(.A(G85), .ZN(new_n600));
  INV_X1    g175(.A(G47), .ZN(new_n601));
  OAI22_X1  g176(.A1(new_n539), .A2(new_n600), .B1(new_n541), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT74), .Z(new_n606));
  NAND2_X1  g181(.A1(new_n545), .A2(G92), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT10), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n537), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(new_n555), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n547), .A2(G54), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n606), .B1(G868), .B2(new_n614), .ZN(G284));
  OAI21_X1  g190(.A(new_n606), .B1(G868), .B2(new_n614), .ZN(G321));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NOR2_X1   g192(.A1(G168), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n580), .B2(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(KEYINPUT75), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(KEYINPUT75), .B2(new_n618), .ZN(G297));
  OAI21_X1  g197(.A(new_n621), .B1(KEYINPUT75), .B2(new_n618), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n614), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n614), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n565), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n501), .A2(G123), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT76), .ZN(new_n631));
  OAI221_X1 g206(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n477), .C2(G111), .ZN(new_n632));
  INV_X1    g207(.A(new_n497), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G135), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n517), .A2(new_n460), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT12), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT13), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2100), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n636), .A2(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2435), .ZN(new_n649));
  XOR2_X1   g224(.A(G2427), .B(G2438), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT14), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n647), .B(new_n652), .Z(new_n653));
  AND2_X1   g228(.A1(new_n653), .A2(G14), .ZN(G401));
  XNOR2_X1  g229(.A(KEYINPUT77), .B(KEYINPUT18), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g233(.A1(new_n658), .A2(KEYINPUT17), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n658), .B2(new_n655), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n661), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2096), .B(G2100), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n668), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  AOI22_X1  g249(.A1(new_n672), .A2(KEYINPUT20), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n674), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n676), .A2(new_n668), .A3(new_n671), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n675), .B(new_n677), .C1(KEYINPUT20), .C2(new_n672), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT78), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1981), .B(G1986), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G229));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G23), .ZN(new_n687));
  INV_X1    g262(.A(G288), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n688), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT82), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT33), .B(G1976), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n686), .A2(G22), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G166), .B2(new_n686), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1971), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n686), .A2(G6), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G305), .B2(G16), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT32), .B(G1981), .Z(new_n698));
  AOI21_X1  g273(.A(new_n695), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n692), .B(new_n699), .C1(new_n697), .C2(new_n698), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT34), .Z(new_n701));
  NAND2_X1  g276(.A1(new_n686), .A2(G24), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(new_n603), .B2(new_n686), .ZN(new_n703));
  INV_X1    g278(.A(G1986), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G25), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n633), .A2(G131), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT79), .Z(new_n709));
  NAND2_X1  g284(.A1(new_n501), .A2(G119), .ZN(new_n710));
  OAI221_X1 g285(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n477), .C2(G107), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT80), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n707), .B1(new_n714), .B2(new_n706), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT81), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT35), .B(G1991), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n716), .B(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n701), .A2(new_n705), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT36), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT31), .B(G11), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n614), .A2(new_n686), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G4), .B2(new_n686), .ZN(new_n724));
  INV_X1    g299(.A(G1348), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  NAND2_X1  g302(.A1(G168), .A2(G16), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G16), .B2(G21), .ZN(new_n729));
  INV_X1    g304(.A(G1966), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT87), .ZN(new_n732));
  NOR2_X1   g307(.A1(G5), .A2(G16), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G171), .B2(G16), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G1961), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n726), .A2(new_n727), .A3(new_n732), .A4(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT89), .B(KEYINPUT23), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n686), .A2(G20), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n580), .B2(new_n686), .ZN(new_n740));
  INV_X1    g315(.A(G1956), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n686), .A2(G19), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n565), .B2(new_n686), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G1341), .ZN(new_n745));
  INV_X1    g320(.A(G28), .ZN(new_n746));
  AOI21_X1  g321(.A(G29), .B1(new_n746), .B2(KEYINPUT30), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(KEYINPUT30), .B2(new_n746), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n729), .B2(new_n730), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n742), .B(new_n750), .C1(new_n734), .C2(G1961), .ZN(new_n751));
  NOR2_X1   g326(.A1(G29), .A2(G32), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n501), .A2(G129), .ZN(new_n753));
  NAND3_X1  g328(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT26), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n633), .A2(G141), .B1(G105), .B2(new_n460), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n753), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n752), .B1(new_n759), .B2(G29), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT27), .B(G1996), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT85), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  OR2_X1    g338(.A1(KEYINPUT24), .A2(G34), .ZN(new_n764));
  NAND2_X1  g339(.A1(KEYINPUT24), .A2(G34), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n764), .A2(new_n706), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G160), .B2(new_n706), .ZN(new_n767));
  OAI221_X1 g342(.A(new_n763), .B1(G2084), .B2(new_n767), .C1(new_n635), .C2(new_n706), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n736), .A2(new_n751), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n706), .A2(G35), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G162), .B2(new_n706), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT29), .ZN(new_n772));
  INV_X1    g347(.A(G2090), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G27), .A2(G29), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G164), .B2(G29), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT88), .B(G2078), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n706), .A2(G26), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT28), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n501), .A2(G128), .ZN(new_n781));
  OAI221_X1 g356(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n477), .C2(G116), .ZN(new_n782));
  INV_X1    g357(.A(G140), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n497), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n785), .A2(new_n706), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT83), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n786), .A2(new_n787), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n780), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G2067), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n769), .A2(new_n774), .A3(new_n778), .A4(new_n793), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n517), .A2(G127), .ZN(new_n795));
  AND2_X1   g370(.A1(G115), .A2(G2104), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n478), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n633), .A2(G139), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n477), .A2(G103), .A3(G2104), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT25), .Z(new_n800));
  AND3_X1   g375(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(G29), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G29), .B2(G33), .ZN(new_n803));
  INV_X1    g378(.A(G2072), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT84), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n760), .A2(new_n762), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G2084), .B2(new_n767), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n806), .B(new_n808), .C1(new_n804), .C2(new_n803), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT86), .Z(new_n810));
  NOR2_X1   g385(.A1(new_n794), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n721), .A2(new_n722), .A3(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(G311));
  XOR2_X1   g388(.A(new_n812), .B(KEYINPUT90), .Z(G150));
  NOR2_X1   g389(.A1(new_n613), .A2(new_n624), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT38), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n545), .A2(G93), .B1(G55), .B2(new_n547), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n537), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n555), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n565), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT91), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n819), .B(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n820), .B1(new_n823), .B2(new_n565), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n816), .B(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT39), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT92), .ZN(new_n828));
  INV_X1    g403(.A(G860), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n828), .B(new_n829), .C1(new_n826), .C2(new_n825), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n822), .A2(new_n829), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT94), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT93), .B(KEYINPUT37), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n830), .A2(new_n834), .ZN(G145));
  XNOR2_X1  g410(.A(new_n635), .B(G162), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G160), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n638), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n501), .A2(G130), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT96), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT97), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n843), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n844), .B(new_n845), .C1(G118), .C2(new_n477), .ZN(new_n846));
  INV_X1    g421(.A(G142), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n841), .B(new_n846), .C1(new_n847), .C2(new_n497), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n848), .A2(new_n714), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT98), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n714), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n850), .B1(new_n849), .B2(new_n851), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n839), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n854), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n856), .A2(new_n852), .A3(new_n638), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n855), .A2(new_n857), .A3(KEYINPUT99), .ZN(new_n858));
  AOI21_X1  g433(.A(KEYINPUT99), .B1(new_n855), .B2(new_n857), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT95), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n801), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n785), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n477), .A2(KEYINPUT4), .A3(G138), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(new_n508), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n506), .B1(new_n864), .B2(new_n491), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(new_n522), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n862), .B(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n759), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n858), .A2(new_n859), .A3(new_n868), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n859), .A2(new_n868), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n838), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OR3_X1    g448(.A1(new_n869), .A2(new_n870), .A3(new_n838), .ZN(new_n874));
  INV_X1    g449(.A(G37), .ZN(new_n875));
  OAI211_X1 g450(.A(KEYINPUT100), .B(new_n838), .C1(new_n869), .C2(new_n870), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n873), .A2(new_n874), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(KEYINPUT40), .ZN(new_n878));
  AOI21_X1  g453(.A(G37), .B1(new_n871), .B2(new_n872), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT40), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n879), .A2(new_n880), .A3(new_n874), .A4(new_n876), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n878), .A2(new_n881), .ZN(G395));
  AOI21_X1  g457(.A(KEYINPUT101), .B1(new_n613), .B2(new_n580), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n613), .B(new_n580), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n883), .B1(new_n884), .B2(KEYINPUT101), .ZN(new_n885));
  OR3_X1    g460(.A1(new_n885), .A2(KEYINPUT102), .A3(KEYINPUT41), .ZN(new_n886));
  OAI21_X1  g461(.A(KEYINPUT102), .B1(new_n885), .B2(KEYINPUT41), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n886), .B(new_n887), .C1(new_n888), .C2(new_n884), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n824), .B(new_n626), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n884), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n891), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(G166), .B(G288), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(G305), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n603), .B(KEYINPUT103), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n895), .B(new_n896), .Z(new_n897));
  XNOR2_X1  g472(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n897), .B(new_n898), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n893), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n893), .A2(new_n899), .ZN(new_n901));
  OAI21_X1  g476(.A(G868), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n823), .A2(new_n617), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(G331));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n905));
  XNOR2_X1  g480(.A(G331), .B(new_n905), .ZN(G295));
  INV_X1    g481(.A(new_n897), .ZN(new_n907));
  NAND2_X1  g482(.A1(G286), .A2(KEYINPUT106), .ZN(new_n908));
  NAND2_X1  g483(.A1(G301), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n824), .B(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(G286), .A2(KEYINPUT106), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n910), .B(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n892), .B1(new_n912), .B2(new_n888), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n912), .A2(new_n888), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n907), .B(new_n913), .C1(new_n914), .C2(new_n885), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n892), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n889), .B2(new_n912), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n897), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(new_n918), .A3(new_n875), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n915), .A2(new_n918), .A3(KEYINPUT108), .A4(new_n875), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(KEYINPUT43), .A3(new_n922), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n916), .B(new_n907), .C1(new_n889), .C2(new_n912), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n918), .A2(new_n875), .A3(new_n924), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n925), .A2(KEYINPUT43), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(KEYINPUT44), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(KEYINPUT43), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n915), .A2(new_n918), .A3(new_n929), .A4(new_n875), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT44), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n931), .A2(KEYINPUT107), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n933));
  AOI211_X1 g508(.A(new_n933), .B(KEYINPUT44), .C1(new_n928), .C2(new_n930), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n927), .B1(new_n932), .B2(new_n934), .ZN(G397));
  INV_X1    g510(.A(KEYINPUT127), .ZN(new_n936));
  INV_X1    g511(.A(G1384), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n937), .B1(new_n513), .B2(new_n518), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n938), .A2(KEYINPUT109), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(KEYINPUT109), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n471), .B1(new_n515), .B2(new_n516), .ZN(new_n943));
  INV_X1    g518(.A(new_n463), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n478), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n945), .A2(new_n494), .A3(G40), .A4(new_n461), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n785), .A2(new_n792), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n781), .A2(G2067), .A3(new_n784), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G1996), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n759), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n758), .A2(G1996), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n952), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n714), .A2(new_n718), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n713), .A2(new_n717), .ZN(new_n959));
  OR3_X1    g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(G1986), .B2(G290), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n603), .A2(new_n704), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n948), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n519), .A2(new_n937), .A3(new_n525), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n946), .B1(new_n964), .B2(KEYINPUT50), .ZN(new_n965));
  AOI21_X1  g540(.A(G1384), .B1(new_n865), .B2(new_n522), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n965), .A2(new_n773), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n964), .A2(new_n941), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n946), .B1(KEYINPUT45), .B2(new_n966), .ZN(new_n971));
  AOI21_X1  g546(.A(G1971), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT110), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n965), .A2(new_n773), .A3(new_n968), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n970), .A2(new_n971), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n974), .B(new_n975), .C1(new_n976), .C2(G1971), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n973), .A2(G8), .A3(new_n977), .ZN(new_n978));
  OAI211_X1 g553(.A(KEYINPUT111), .B(G8), .C1(new_n536), .C2(new_n543), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT55), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n983));
  OAI21_X1  g558(.A(G8), .B1(new_n536), .B2(new_n543), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n984), .A2(new_n985), .A3(new_n983), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n982), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n988), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n990), .A2(new_n986), .A3(new_n981), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n978), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(G305), .A2(G1981), .ZN(new_n994));
  INV_X1    g569(.A(G1981), .ZN(new_n995));
  AOI22_X1  g570(.A1(new_n591), .A2(new_n593), .B1(G86), .B2(new_n545), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n995), .B1(new_n996), .B2(new_n595), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT49), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(G305), .A2(G1981), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT49), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n996), .A2(new_n995), .A3(new_n595), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n946), .A2(new_n938), .ZN(new_n1003));
  INV_X1    g578(.A(G8), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT114), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1006), .B(G8), .C1(new_n946), .C2(new_n938), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n998), .A2(new_n1002), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n688), .A2(G1976), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1011));
  INV_X1    g586(.A(G1976), .ZN(new_n1012));
  NAND2_X1  g587(.A1(G288), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1013), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1009), .B(new_n1011), .C1(new_n1014), .C2(KEYINPUT52), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n966), .A2(new_n479), .A3(G40), .A4(new_n494), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1006), .B1(new_n1016), .B2(G8), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1007), .ZN(new_n1018));
  OAI211_X1 g593(.A(KEYINPUT115), .B(new_n1009), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1013), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1008), .B1(new_n1015), .B2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n519), .A2(new_n525), .A3(KEYINPUT45), .A4(new_n937), .ZN(new_n1025));
  INV_X1    g600(.A(new_n946), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n938), .A2(new_n941), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n730), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n964), .A2(KEYINPUT50), .ZN(new_n1030));
  INV_X1    g605(.A(G2084), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1030), .A2(new_n1031), .A3(new_n1026), .A4(new_n968), .ZN(new_n1032));
  AOI211_X1 g607(.A(new_n1004), .B(G286), .C1(new_n1029), .C2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n993), .A2(new_n1024), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT63), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n519), .A2(new_n525), .A3(new_n967), .A4(new_n937), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n938), .A2(KEYINPUT50), .ZN(new_n1037));
  AND4_X1   g612(.A1(new_n773), .A2(new_n1036), .A3(new_n1026), .A4(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(G8), .B1(new_n972), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT63), .B1(new_n1039), .B2(new_n992), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n1033), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT113), .B1(new_n989), .B2(new_n991), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n981), .B1(new_n990), .B2(new_n986), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n987), .A2(new_n982), .A3(new_n988), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1042), .A2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1047), .A2(new_n973), .A3(G8), .A4(new_n977), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1041), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1050));
  OR3_X1    g625(.A1(new_n1008), .A2(G1976), .A3(G288), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n1001), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1049), .A2(new_n1024), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1035), .A2(new_n1053), .ZN(new_n1054));
  AOI221_X4 g629(.A(new_n1008), .B1(new_n1039), .B2(new_n992), .C1(new_n1015), .C2(new_n1023), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(G8), .ZN(new_n1057));
  NOR2_X1   g632(.A1(G168), .A2(new_n1004), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1057), .A2(KEYINPUT51), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1061), .B(G8), .C1(new_n1056), .C2(G286), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT120), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1056), .A2(KEYINPUT120), .A3(new_n1058), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1060), .B(new_n1062), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G2078), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n970), .A2(new_n971), .A3(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1030), .A2(new_n1026), .A3(new_n968), .ZN(new_n1070));
  INV_X1    g645(.A(G1961), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1066), .A2(KEYINPUT53), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .A4(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1069), .A2(new_n1072), .A3(G301), .A4(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT124), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1067), .A2(new_n1068), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1077), .A2(new_n1078), .A3(G301), .A4(new_n1074), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n942), .A2(new_n971), .A3(new_n1073), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1069), .A2(new_n1072), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G171), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1076), .A2(new_n1079), .A3(new_n1082), .A4(KEYINPUT54), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1055), .A2(new_n1065), .A3(new_n1083), .A4(new_n1048), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1069), .A2(new_n1072), .A3(G301), .A4(new_n1080), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT122), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1077), .A2(new_n1087), .A3(G301), .A4(new_n1080), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1069), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G171), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1086), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT123), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(new_n1095), .A3(new_n1092), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1084), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT56), .B(G2072), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n970), .A2(new_n971), .A3(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1036), .A2(new_n1026), .A3(new_n1037), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1100), .A2(new_n1101), .A3(new_n741), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1101), .B1(new_n1100), .B2(new_n741), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1099), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1105), .B1(new_n579), .B2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n580), .B(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1104), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1016), .A2(G2067), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(new_n1070), .B2(new_n725), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1110), .B1(new_n613), .B2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1108), .B(new_n1099), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT118), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1100), .A2(new_n741), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1100), .A2(new_n1101), .A3(new_n741), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1119), .A2(new_n1120), .A3(new_n1108), .A4(new_n1099), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1113), .A2(new_n1115), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1115), .A2(new_n1121), .A3(new_n1110), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1110), .A2(KEYINPUT61), .A3(new_n1114), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n613), .B1(new_n1112), .B2(KEYINPUT60), .ZN(new_n1127));
  AOI21_X1  g702(.A(G1348), .B1(new_n965), .B2(new_n968), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT60), .ZN(new_n1129));
  NOR4_X1   g704(.A1(new_n1128), .A2(new_n614), .A3(new_n1129), .A4(new_n1111), .ZN(new_n1130));
  OAI22_X1  g705(.A1(new_n1127), .A2(new_n1130), .B1(KEYINPUT60), .B2(new_n1112), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n970), .A2(new_n971), .A3(new_n953), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  OR2_X1    g710(.A1(KEYINPUT58), .A2(G1341), .ZN(new_n1136));
  NAND2_X1  g711(.A1(KEYINPUT58), .A2(G1341), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1016), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n970), .A2(new_n971), .A3(KEYINPUT119), .A4(new_n953), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1135), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1132), .B1(new_n1140), .B2(new_n565), .ZN(new_n1141));
  AND3_X1   g716(.A1(new_n1140), .A2(new_n1132), .A3(new_n565), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1126), .B(new_n1131), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1122), .B1(new_n1125), .B2(new_n1143), .ZN(new_n1144));
  AOI211_X1 g719(.A(KEYINPUT125), .B(new_n1054), .C1(new_n1097), .C2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1084), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1144), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1054), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1146), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1145), .A2(new_n1151), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1055), .A2(new_n1048), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n1065), .A2(KEYINPUT62), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1090), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1065), .A2(KEYINPUT62), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n963), .B1(new_n1152), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n950), .B1(new_n956), .B2(new_n959), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1159), .A2(new_n948), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT126), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n948), .A2(new_n962), .ZN(new_n1162));
  XOR2_X1   g737(.A(new_n1162), .B(KEYINPUT48), .Z(new_n1163));
  INV_X1    g738(.A(new_n960), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1163), .B1(new_n1164), .B2(new_n948), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n948), .A2(G1996), .ZN(new_n1166));
  OR2_X1    g741(.A1(new_n1166), .A2(KEYINPUT46), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n947), .B1(new_n952), .B2(new_n758), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1166), .A2(KEYINPUT46), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT47), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1161), .A2(new_n1165), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n936), .B1(new_n1158), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1172), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1157), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1145), .A2(new_n1151), .A3(new_n1175), .ZN(new_n1176));
  OAI211_X1 g751(.A(KEYINPUT127), .B(new_n1174), .C1(new_n1176), .C2(new_n963), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1173), .A2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g753(.A(G319), .ZN(new_n1180));
  AOI211_X1 g754(.A(new_n1180), .B(G229), .C1(new_n928), .C2(new_n930), .ZN(new_n1181));
  NOR2_X1   g755(.A1(G401), .A2(G227), .ZN(new_n1182));
  AND3_X1   g756(.A1(new_n1181), .A2(new_n877), .A3(new_n1182), .ZN(G308));
  NAND3_X1  g757(.A1(new_n1181), .A2(new_n877), .A3(new_n1182), .ZN(G225));
endmodule


