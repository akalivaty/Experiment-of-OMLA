//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT89), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT81), .A2(G104), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT81), .A2(G104), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n192), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT3), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(new_n192), .A3(G104), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT82), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n197), .A2(new_n192), .A3(KEYINPUT82), .A4(G104), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G101), .ZN(new_n203));
  OR2_X1    g017(.A1(KEYINPUT81), .A2(G104), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT81), .A2(G104), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(G107), .A3(new_n205), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n196), .A2(new_n202), .A3(new_n203), .A4(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT4), .ZN(new_n208));
  NOR3_X1   g022(.A1(new_n193), .A2(new_n194), .A3(new_n192), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n209), .B1(KEYINPUT3), .B2(new_n195), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n203), .B1(new_n210), .B2(new_n202), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT2), .A2(G113), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT2), .A2(G113), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n213), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G119), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G116), .ZN(new_n220));
  INV_X1    g034(.A(G116), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G119), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n218), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n221), .A2(G119), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n219), .A2(G116), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n220), .A2(new_n222), .A3(KEYINPUT69), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n227), .B(new_n228), .C1(new_n218), .C2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n217), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n232));
  OAI22_X1  g046(.A1(new_n231), .A2(new_n232), .B1(KEYINPUT2), .B2(G113), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(KEYINPUT68), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n223), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT4), .ZN(new_n236));
  AOI21_X1  g050(.A(G107), .B1(new_n204), .B2(new_n205), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n206), .B1(new_n237), .B2(new_n197), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n200), .A2(new_n201), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n236), .B(G101), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT85), .B1(new_n212), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(G110), .B(G122), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n220), .A2(new_n222), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n233), .A2(new_n244), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n220), .A2(new_n222), .A3(KEYINPUT69), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT69), .B1(new_n220), .B2(new_n222), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT5), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(G113), .B1(new_n220), .B2(KEYINPUT5), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n245), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n192), .A2(G104), .ZN(new_n252));
  OAI21_X1  g066(.A(G101), .B1(new_n237), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n251), .A2(new_n207), .A3(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(G101), .B1(new_n238), .B2(new_n239), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(KEYINPUT4), .A3(new_n207), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT85), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n256), .A2(new_n257), .A3(new_n235), .A4(new_n240), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n242), .A2(new_n243), .A3(new_n254), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n207), .A2(new_n253), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n260), .A2(new_n251), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n244), .A2(new_n262), .ZN(new_n263));
  OAI22_X1  g077(.A1(new_n263), .A2(new_n249), .B1(new_n233), .B2(new_n244), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n207), .A2(new_n264), .A3(new_n253), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n243), .B(KEYINPUT8), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT88), .B1(new_n261), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n260), .A2(new_n251), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT88), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n269), .A2(new_n270), .A3(new_n266), .A4(new_n265), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G146), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G143), .ZN(new_n274));
  INV_X1    g088(.A(G143), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G146), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n274), .A2(KEYINPUT1), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(new_n278), .A3(G128), .ZN(new_n279));
  INV_X1    g093(.A(G125), .ZN(new_n280));
  INV_X1    g094(.A(G128), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n274), .B(new_n276), .C1(KEYINPUT1), .C2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(G143), .B(G146), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(KEYINPUT0), .A3(G128), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT0), .B(G128), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n285), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n283), .B1(new_n287), .B2(new_n280), .ZN(new_n288));
  INV_X1    g102(.A(G953), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G224), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n290), .A2(KEYINPUT7), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n288), .B(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n259), .A2(new_n272), .A3(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n191), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n292), .B1(new_n268), .B2(new_n271), .ZN(new_n297));
  AOI211_X1 g111(.A(KEYINPUT89), .B(G902), .C1(new_n297), .C2(new_n259), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  XOR2_X1   g113(.A(new_n290), .B(KEYINPUT87), .Z(new_n300));
  XNOR2_X1  g114(.A(new_n288), .B(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT6), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n303), .A2(KEYINPUT86), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n259), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n243), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n258), .A2(new_n254), .ZN(new_n307));
  INV_X1    g121(.A(new_n241), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n257), .B1(new_n308), .B2(new_n256), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n306), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n306), .B(new_n304), .C1(new_n307), .C2(new_n309), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n302), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n190), .B1(new_n299), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n294), .A2(new_n295), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT89), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n294), .A2(new_n191), .A3(new_n295), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n311), .A2(new_n312), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n301), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n189), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n188), .B1(new_n314), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G214), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n323), .A2(G237), .A3(G953), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n275), .A2(KEYINPUT90), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT90), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G143), .ZN(new_n328));
  NOR2_X1   g142(.A1(G237), .A2(G953), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n328), .A2(new_n325), .B1(new_n329), .B2(G214), .ZN(new_n330));
  AND2_X1   g144(.A1(KEYINPUT18), .A2(G131), .ZN(new_n331));
  OAI22_X1  g145(.A1(new_n326), .A2(new_n330), .B1(KEYINPUT91), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(KEYINPUT91), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n324), .A2(new_n325), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n328), .A2(new_n325), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n335), .B1(new_n336), .B2(new_n324), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(KEYINPUT91), .A3(new_n331), .ZN(new_n338));
  INV_X1    g152(.A(G140), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G125), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n280), .A2(G140), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n280), .A2(KEYINPUT77), .A3(G140), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n343), .A2(KEYINPUT92), .A3(G146), .A4(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n346));
  XNOR2_X1  g160(.A(G125), .B(G140), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n346), .B1(new_n347), .B2(new_n273), .ZN(new_n348));
  AND4_X1   g162(.A1(new_n346), .A2(new_n340), .A3(new_n341), .A4(new_n273), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n343), .A2(new_n344), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT92), .B1(new_n351), .B2(G146), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n334), .B(new_n338), .C1(new_n350), .C2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(G131), .B1(new_n326), .B2(new_n330), .ZN(new_n354));
  INV_X1    g168(.A(G131), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n355), .B(new_n335), .C1(new_n336), .C2(new_n324), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n343), .A2(KEYINPUT16), .A3(new_n344), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT16), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n340), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G146), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT19), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(new_n343), .B2(new_n344), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n347), .A2(KEYINPUT19), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n273), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n357), .A2(new_n362), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n353), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(G113), .B(G122), .ZN(new_n369));
  XOR2_X1   g183(.A(new_n369), .B(G104), .Z(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n373), .B1(new_n361), .B2(G146), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n358), .A2(KEYINPUT78), .A3(new_n273), .A4(new_n360), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n362), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n337), .A2(KEYINPUT17), .A3(G131), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n377), .B1(new_n357), .B2(KEYINPUT17), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n353), .B(new_n370), .C1(new_n376), .C2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n372), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(G475), .A2(G902), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT20), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT20), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n380), .A2(new_n384), .A3(new_n381), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n353), .B1(new_n376), .B2(new_n378), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n371), .ZN(new_n388));
  AOI21_X1  g202(.A(G902), .B1(new_n388), .B2(new_n379), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G475), .ZN(new_n391));
  INV_X1    g205(.A(G478), .ZN(new_n392));
  NOR2_X1   g206(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n392), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n221), .A2(G122), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n192), .B1(new_n398), .B2(KEYINPUT14), .ZN(new_n399));
  XOR2_X1   g213(.A(G116), .B(G122), .Z(new_n400));
  OR2_X1    g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n400), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n281), .A2(G143), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT93), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n403), .B(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n281), .A2(G143), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n405), .A2(G134), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G134), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n403), .B(KEYINPUT93), .ZN(new_n409));
  INV_X1    g223(.A(new_n406), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n401), .B(new_n402), .C1(new_n407), .C2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n406), .B(KEYINPUT13), .ZN(new_n413));
  OAI21_X1  g227(.A(G134), .B1(new_n413), .B2(new_n405), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n400), .B(G107), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n409), .A2(new_n408), .A3(new_n410), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  XOR2_X1   g232(.A(KEYINPUT76), .B(G217), .Z(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT9), .B(G234), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n419), .A2(G953), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n412), .A2(new_n417), .A3(new_n421), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n397), .B1(new_n425), .B2(new_n295), .ZN(new_n426));
  AOI211_X1 g240(.A(G902), .B(new_n396), .C1(new_n423), .C2(new_n424), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n289), .A2(G952), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(G234), .B2(G237), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(G898), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(G234), .A2(G237), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(G902), .A3(G953), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n431), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n386), .A2(new_n391), .A3(new_n428), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT95), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n383), .A2(new_n385), .B1(new_n390), .B2(G475), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT95), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n439), .A2(new_n440), .A3(new_n428), .A4(new_n436), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(G221), .B1(new_n420), .B2(G902), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  XOR2_X1   g258(.A(KEYINPUT83), .B(G469), .Z(new_n445));
  INV_X1    g259(.A(new_n287), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n256), .A2(new_n446), .A3(new_n240), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT64), .ZN(new_n448));
  INV_X1    g262(.A(G137), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n448), .B1(new_n449), .B2(G134), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n408), .A2(KEYINPUT64), .A3(G137), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT11), .B1(new_n408), .B2(G137), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT11), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(new_n449), .A3(G134), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n355), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n456), .A2(new_n355), .A3(new_n450), .A4(new_n451), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT65), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n452), .A2(KEYINPUT65), .A3(new_n355), .A4(new_n456), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n457), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT10), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n279), .A2(new_n282), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n463), .B1(new_n260), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n464), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n466), .A2(new_n207), .A3(KEYINPUT10), .A4(new_n253), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n447), .A2(new_n462), .A3(new_n465), .A4(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(G110), .B(G140), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(KEYINPUT80), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n289), .A2(G227), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n470), .B(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n260), .B(new_n464), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n460), .A2(new_n461), .ZN(new_n474));
  INV_X1    g288(.A(new_n457), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT12), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n260), .A2(new_n464), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n466), .B1(new_n207), .B2(new_n253), .ZN(new_n479));
  OAI211_X1 g293(.A(KEYINPUT12), .B(new_n476), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n468), .B(new_n472), .C1(new_n477), .C2(new_n481), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n256), .A2(new_n446), .A3(new_n240), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n465), .A2(new_n467), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n476), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n472), .B1(new_n485), .B2(new_n468), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT84), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n482), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI211_X1 g302(.A(KEYINPUT84), .B(new_n472), .C1(new_n485), .C2(new_n468), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n295), .B(new_n445), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n468), .B1(new_n477), .B2(new_n481), .ZN(new_n491));
  INV_X1    g305(.A(new_n472), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n468), .A2(new_n472), .ZN(new_n493));
  AOI22_X1  g307(.A1(new_n491), .A2(new_n492), .B1(new_n493), .B2(new_n485), .ZN(new_n494));
  OAI21_X1  g308(.A(G469), .B1(new_n494), .B2(G902), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n444), .B1(new_n490), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n322), .A2(new_n442), .A3(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n408), .A2(G137), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n449), .A2(G134), .ZN(new_n499));
  OAI21_X1  g313(.A(G131), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n279), .A2(new_n500), .A3(new_n282), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n474), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n235), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n503), .B(new_n504), .C1(new_n462), .C2(new_n287), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT73), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT28), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n506), .B1(new_n505), .B2(new_n507), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XOR2_X1   g324(.A(KEYINPUT26), .B(G101), .Z(new_n511));
  NAND2_X1  g325(.A1(new_n329), .A2(G210), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  XOR2_X1   g329(.A(new_n515), .B(KEYINPUT72), .Z(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n505), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT66), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n476), .B2(new_n446), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n462), .A2(KEYINPUT66), .A3(new_n287), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n503), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n518), .B1(new_n522), .B2(new_n235), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n510), .B(new_n517), .C1(new_n523), .C2(new_n507), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT29), .ZN(new_n525));
  INV_X1    g339(.A(new_n515), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n503), .B(KEYINPUT30), .C1(new_n462), .C2(new_n287), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n235), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT30), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n528), .B1(new_n522), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n526), .B1(new_n530), .B2(new_n518), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n524), .A2(new_n525), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT74), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n462), .A2(new_n287), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n501), .B1(new_n460), .B2(new_n461), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n235), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n505), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n533), .B1(new_n537), .B2(KEYINPUT28), .ZN(new_n538));
  AOI211_X1 g352(.A(KEYINPUT74), .B(new_n507), .C1(new_n536), .C2(new_n505), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n510), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n515), .A2(KEYINPUT29), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n295), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(G472), .B1(new_n532), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT32), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT31), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n505), .A2(KEYINPUT71), .A3(new_n515), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT71), .B1(new_n505), .B2(new_n515), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n545), .B1(new_n548), .B2(new_n530), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n505), .A2(new_n515), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT71), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n505), .A2(KEYINPUT71), .A3(new_n515), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n476), .A2(new_n519), .A3(new_n446), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT66), .B1(new_n462), .B2(new_n287), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n535), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n235), .B(new_n527), .C1(new_n557), .C2(KEYINPUT30), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n554), .A2(new_n558), .A3(KEYINPUT31), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n549), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n522), .A2(new_n235), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n507), .B1(new_n561), .B2(new_n505), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n508), .A2(new_n509), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n516), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(G472), .A2(G902), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n544), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n566), .ZN(new_n568));
  AOI211_X1 g382(.A(KEYINPUT32), .B(new_n568), .C1(new_n560), .C2(new_n564), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n543), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT75), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n510), .B1(new_n523), .B2(new_n507), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n549), .A2(new_n559), .B1(new_n572), .B2(new_n516), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT32), .B1(new_n573), .B2(new_n568), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n565), .A2(new_n544), .A3(new_n566), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT75), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(new_n577), .A3(new_n543), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT23), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n219), .B2(G128), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n281), .A2(KEYINPUT23), .A3(G119), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n580), .B(new_n581), .C1(G119), .C2(new_n281), .ZN(new_n582));
  XNOR2_X1  g396(.A(G119), .B(G128), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT24), .B(G110), .Z(new_n584));
  AOI22_X1  g398(.A1(new_n582), .A2(G110), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n376), .A2(new_n585), .ZN(new_n586));
  OAI22_X1  g400(.A1(new_n582), .A2(G110), .B1(new_n583), .B2(new_n584), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n362), .B(new_n587), .C1(new_n349), .C2(new_n348), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT22), .B(G137), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n289), .A2(G221), .A3(G234), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n586), .A2(new_n588), .A3(new_n592), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n295), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT25), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n419), .B1(G234), .B2(new_n295), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n594), .A2(new_n595), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n599), .A2(G902), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n497), .A2(new_n571), .A3(new_n578), .A4(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  NAND2_X1  g421(.A1(new_n314), .A2(new_n321), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n187), .ZN(new_n609));
  INV_X1    g423(.A(new_n436), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n392), .A2(new_n295), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n425), .A2(new_n295), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n612), .B1(new_n613), .B2(G478), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n425), .B(KEYINPUT33), .Z(new_n615));
  AOI21_X1  g429(.A(new_n614), .B1(new_n615), .B2(G478), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n380), .A2(new_n384), .A3(new_n381), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n384), .B1(new_n380), .B2(new_n381), .ZN(new_n618));
  INV_X1    g432(.A(G475), .ZN(new_n619));
  OAI22_X1  g433(.A1(new_n617), .A2(new_n618), .B1(new_n619), .B2(new_n389), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n609), .A2(new_n610), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n565), .A2(new_n566), .ZN(new_n623));
  OAI21_X1  g437(.A(G472), .B1(new_n573), .B2(G902), .ZN(new_n624));
  AND4_X1   g438(.A1(new_n623), .A2(new_n605), .A3(new_n496), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT34), .B(G104), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT96), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n626), .B(new_n628), .ZN(G6));
  NOR2_X1   g443(.A1(new_n609), .A2(new_n610), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n620), .A2(new_n428), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n625), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  OR2_X1    g448(.A1(new_n593), .A2(KEYINPUT36), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n589), .B(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n602), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n598), .B2(new_n599), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(new_n438), .B2(new_n441), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n322), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n641), .A2(new_n623), .A3(new_n496), .A4(new_n624), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT37), .B(G110), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G12));
  INV_X1    g458(.A(new_n639), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n496), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n571), .A2(new_n578), .A3(new_n322), .A4(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n289), .A2(G900), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(G902), .A3(new_n434), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT97), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n651), .A2(new_n431), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n631), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n647), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G128), .ZN(G30));
  INV_X1    g470(.A(KEYINPUT38), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n608), .B(new_n657), .ZN(new_n658));
  AOI22_X1  g472(.A1(new_n554), .A2(new_n558), .B1(new_n516), .B2(new_n537), .ZN(new_n659));
  OAI21_X1  g473(.A(G472), .B1(new_n659), .B2(G902), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n576), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n439), .A2(new_n428), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n639), .A2(new_n187), .A3(new_n663), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n658), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n653), .B(KEYINPUT39), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n496), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n665), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT98), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G143), .ZN(G45));
  INV_X1    g487(.A(new_n653), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n621), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n647), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n273), .ZN(G48));
  AND3_X1   g492(.A1(new_n571), .A2(new_n578), .A3(new_n605), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n295), .B1(new_n488), .B2(new_n489), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(G469), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n681), .A2(new_n443), .A3(new_n490), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n679), .A2(KEYINPUT99), .A3(new_n622), .A4(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT99), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n571), .A2(new_n578), .A3(new_n605), .A4(new_n682), .ZN(new_n685));
  INV_X1    g499(.A(new_n622), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT41), .B(G113), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G15));
  NAND2_X1  g504(.A1(new_n630), .A2(new_n631), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n221), .ZN(G18));
  NAND4_X1  g507(.A1(new_n571), .A2(new_n641), .A3(new_n578), .A4(new_n682), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G119), .ZN(G21));
  AND3_X1   g509(.A1(new_n608), .A2(new_n187), .A3(new_n663), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT100), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n540), .A2(new_n697), .ZN(new_n698));
  OAI211_X1 g512(.A(KEYINPUT100), .B(new_n510), .C1(new_n538), .C2(new_n539), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n516), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n560), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n566), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n702), .A2(new_n605), .A3(new_n624), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n696), .A2(new_n703), .A3(new_n436), .A4(new_n682), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G122), .ZN(G24));
  NAND4_X1  g519(.A1(new_n702), .A2(new_n624), .A3(new_n645), .A4(new_n675), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n682), .A2(new_n322), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT101), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G125), .ZN(G27));
  NAND2_X1  g524(.A1(G469), .A2(G902), .ZN(new_n711));
  XOR2_X1   g525(.A(new_n711), .B(KEYINPUT102), .Z(new_n712));
  AOI21_X1  g526(.A(new_n712), .B1(new_n494), .B2(G469), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n444), .B1(new_n490), .B2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n314), .A2(new_n321), .A3(new_n187), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n717), .A2(new_n570), .A3(new_n605), .A4(new_n675), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT42), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n571), .A2(new_n578), .A3(new_n605), .A4(new_n717), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n676), .A2(KEYINPUT42), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n719), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n355), .ZN(G33));
  NOR2_X1   g538(.A1(new_n720), .A2(new_n654), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n408), .ZN(G36));
  OR2_X1    g540(.A1(new_n494), .A2(KEYINPUT45), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n494), .A2(KEYINPUT45), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(G469), .A3(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n712), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(KEYINPUT46), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n490), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(KEYINPUT103), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT103), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n731), .A2(new_n734), .A3(new_n490), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n729), .A2(new_n730), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT46), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n733), .A2(new_n735), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n443), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n666), .ZN(new_n742));
  INV_X1    g556(.A(new_n616), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT43), .B1(new_n743), .B2(new_n620), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n616), .A2(new_n745), .A3(new_n439), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n639), .B1(new_n624), .B2(new_n623), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(KEYINPUT44), .A3(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n716), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(KEYINPUT44), .B1(new_n747), .B2(new_n748), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n742), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n449), .ZN(G39));
  NAND2_X1  g569(.A1(new_n741), .A2(KEYINPUT47), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT47), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n740), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n750), .A2(new_n604), .A3(new_n675), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n760), .B1(new_n571), .B2(new_n578), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G140), .ZN(G42));
  INV_X1    g577(.A(KEYINPUT105), .ZN(new_n764));
  INV_X1    g578(.A(new_n720), .ZN(new_n765));
  AOI22_X1  g579(.A1(new_n765), .A2(new_n721), .B1(KEYINPUT42), .B2(new_n718), .ZN(new_n766));
  INV_X1    g580(.A(new_n621), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n630), .B(new_n625), .C1(new_n767), .C2(new_n631), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n606), .A2(new_n768), .A3(new_n642), .ZN(new_n769));
  INV_X1    g583(.A(new_n706), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n717), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n571), .A2(new_n578), .A3(new_n646), .ZN(new_n772));
  INV_X1    g586(.A(new_n428), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n620), .A2(new_n773), .A3(new_n674), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n314), .A2(new_n321), .A3(new_n187), .A4(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT104), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n775), .B(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n771), .B1(new_n772), .B2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n725), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n766), .A2(new_n769), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n704), .B(new_n694), .C1(new_n685), .C2(new_n691), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n688), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n764), .B1(new_n781), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n775), .B(KEYINPUT104), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n786), .A2(new_n571), .A3(new_n578), .A4(new_n646), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n787), .B(new_n771), .C1(new_n654), .C2(new_n720), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n606), .A2(new_n768), .A3(new_n642), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n788), .A2(new_n723), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n782), .B1(new_n687), .B2(new_n683), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(KEYINPUT105), .A3(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n785), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n645), .A2(new_n674), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n696), .A2(new_n661), .A3(new_n714), .A4(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  AND4_X1   g610(.A1(new_n571), .A2(new_n578), .A3(new_n322), .A4(new_n646), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n796), .B1(new_n797), .B2(new_n675), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n798), .A2(new_n709), .A3(new_n655), .A4(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n707), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT101), .B1(new_n770), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT101), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n706), .A2(new_n707), .A3(new_n803), .ZN(new_n804));
  OAI22_X1  g618(.A1(new_n802), .A2(new_n804), .B1(new_n647), .B2(new_n654), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n795), .B1(new_n647), .B2(new_n676), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT52), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT106), .B1(new_n800), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n800), .A2(new_n807), .A3(KEYINPUT106), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT53), .B1(new_n793), .B2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n790), .A2(new_n800), .A3(new_n807), .A4(new_n791), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g629(.A(KEYINPUT107), .B(KEYINPUT54), .C1(new_n812), .C2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT107), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n800), .A2(new_n807), .A3(KEYINPUT106), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n785), .B(new_n792), .C1(new_n818), .C2(new_n808), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n815), .B1(new_n819), .B2(new_n814), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n817), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n723), .A2(new_n778), .A3(new_n725), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n791), .A2(new_n823), .A3(new_n769), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n800), .A2(new_n807), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n814), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT108), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(KEYINPUT108), .B(new_n814), .C1(new_n824), .C2(new_n825), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n824), .A2(new_n814), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n828), .A2(new_n829), .B1(new_n811), .B2(new_n830), .ZN(new_n831));
  XOR2_X1   g645(.A(KEYINPUT109), .B(KEYINPUT54), .Z(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n816), .A2(new_n822), .A3(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n744), .A2(new_n430), .A3(new_n746), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n681), .A2(new_n443), .A3(new_n490), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n716), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AOI211_X1 g652(.A(new_n604), .B(new_n838), .C1(new_n576), .C2(new_n543), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n839), .B(KEYINPUT48), .Z(new_n840));
  AND2_X1   g654(.A1(new_n703), .A2(new_n835), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n801), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n604), .A2(new_n431), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n662), .A2(new_n837), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n767), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n429), .B(KEYINPUT115), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n840), .A2(new_n842), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n681), .A2(new_n490), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n444), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n756), .A2(new_n758), .A3(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n841), .A2(new_n750), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n682), .A2(new_n188), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT111), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(new_n658), .A3(new_n841), .ZN(new_n855));
  NOR2_X1   g669(.A1(KEYINPUT112), .A2(KEYINPUT50), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n854), .A2(new_n658), .A3(new_n856), .A4(new_n841), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n702), .A2(new_n624), .A3(new_n645), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n838), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n616), .A2(new_n620), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n861), .B1(new_n844), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n858), .A2(new_n859), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT114), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT114), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n858), .A2(new_n866), .A3(new_n859), .A4(new_n863), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n852), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT51), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n849), .B(KEYINPUT110), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n756), .A2(new_n758), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT51), .B1(new_n871), .B2(new_n851), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n864), .A2(KEYINPUT113), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n864), .A2(KEYINPUT113), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n847), .B1(new_n869), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT116), .ZN(new_n877));
  OAI22_X1  g691(.A1(new_n834), .A2(new_n877), .B1(G952), .B2(G953), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n848), .B(KEYINPUT49), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n605), .A2(new_n187), .A3(new_n443), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n880), .A2(new_n620), .A3(new_n743), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n879), .A2(new_n881), .A3(new_n658), .A4(new_n662), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n878), .A2(new_n882), .ZN(G75));
  NOR2_X1   g697(.A1(new_n289), .A2(G952), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n830), .B1(new_n818), .B2(new_n808), .ZN(new_n885));
  INV_X1    g699(.A(new_n829), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT108), .B1(new_n813), .B2(new_n814), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n888), .A2(G210), .A3(G902), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT56), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n319), .A2(new_n301), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n892), .A2(new_n313), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT55), .Z(new_n894));
  AOI21_X1  g708(.A(new_n884), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT117), .ZN(new_n896));
  INV_X1    g710(.A(new_n894), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n889), .A2(new_n896), .A3(new_n890), .A4(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n889), .A2(new_n890), .A3(new_n897), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT117), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n895), .A2(new_n898), .A3(new_n900), .ZN(G51));
  XNOR2_X1  g715(.A(new_n712), .B(KEYINPUT57), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n831), .A2(new_n832), .ZN(new_n903));
  INV_X1    g717(.A(new_n832), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n888), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n902), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n488), .A2(new_n489), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OR3_X1    g722(.A1(new_n831), .A2(new_n295), .A3(new_n729), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n884), .B1(new_n908), .B2(new_n909), .ZN(G54));
  AND2_X1   g724(.A1(KEYINPUT58), .A2(G475), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n888), .A2(G902), .A3(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n380), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n884), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n888), .A2(G902), .A3(new_n380), .A4(new_n911), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT118), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n914), .A2(KEYINPUT118), .A3(new_n915), .A4(new_n916), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(G60));
  INV_X1    g735(.A(new_n615), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n611), .B(KEYINPUT59), .Z(new_n923));
  AOI21_X1  g737(.A(new_n922), .B1(new_n834), .B2(new_n923), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n903), .B2(new_n905), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n915), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n924), .A2(new_n927), .ZN(G63));
  NAND2_X1  g742(.A1(G217), .A2(G902), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT60), .ZN(new_n930));
  OR3_X1    g744(.A1(new_n831), .A2(new_n636), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n601), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n831), .B2(new_n930), .ZN(new_n933));
  NOR2_X1   g747(.A1(KEYINPUT119), .A2(KEYINPUT61), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n884), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n931), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(KEYINPUT119), .A2(KEYINPUT61), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT120), .Z(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n931), .A2(new_n938), .A3(new_n933), .A4(new_n935), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(G66));
  AOI21_X1  g756(.A(new_n289), .B1(new_n433), .B2(G224), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n784), .A2(new_n789), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n943), .B1(new_n945), .B2(new_n289), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n311), .B(new_n312), .C1(G898), .C2(new_n289), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n946), .B(new_n947), .Z(G69));
  OAI21_X1  g762(.A(new_n527), .B1(new_n557), .B2(KEYINPUT30), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT121), .Z(new_n950));
  OR2_X1    g764(.A1(new_n364), .A2(new_n365), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n950), .B(new_n951), .Z(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n754), .A2(new_n723), .A3(new_n725), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n805), .A2(new_n677), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT123), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n696), .A2(new_n570), .A3(new_n605), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n956), .B1(new_n742), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n957), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n741), .A2(new_n959), .A3(KEYINPUT123), .A4(new_n666), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n954), .A2(new_n762), .A3(new_n955), .A4(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT124), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n962), .A2(new_n963), .ZN(new_n966));
  AOI21_X1  g780(.A(G953), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n953), .B1(new_n967), .B2(new_n648), .ZN(new_n968));
  INV_X1    g782(.A(new_n754), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n767), .A2(new_n631), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n970), .A2(new_n667), .A3(new_n716), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n679), .A2(new_n971), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n762), .A2(new_n969), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n672), .A2(new_n955), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(KEYINPUT62), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n672), .A2(new_n976), .A3(new_n955), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n973), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT122), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n973), .A2(new_n975), .A3(KEYINPUT122), .A4(new_n977), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n289), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n952), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n289), .B1(G227), .B2(G900), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n968), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n962), .A2(new_n963), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n289), .B1(new_n988), .B2(new_n964), .ZN(new_n989));
  INV_X1    g803(.A(new_n648), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n952), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n953), .B1(new_n982), .B2(new_n289), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n985), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n987), .A2(new_n993), .ZN(G72));
  NOR2_X1   g808(.A1(new_n530), .A2(new_n518), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n980), .A2(new_n944), .A3(new_n981), .ZN(new_n996));
  XNOR2_X1  g810(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n997));
  NAND2_X1  g811(.A1(G472), .A2(G902), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n997), .B(new_n998), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT126), .Z(new_n1000));
  AOI211_X1 g814(.A(new_n526), .B(new_n995), .C1(new_n996), .C2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n995), .A2(new_n526), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n965), .A2(new_n944), .A3(new_n966), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1002), .B1(new_n1003), .B2(new_n1000), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n531), .A2(KEYINPUT127), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1005), .B1(new_n530), .B2(new_n548), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n531), .A2(KEYINPUT127), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n999), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n915), .B1(new_n820), .B2(new_n1008), .ZN(new_n1009));
  NOR3_X1   g823(.A1(new_n1001), .A2(new_n1004), .A3(new_n1009), .ZN(G57));
endmodule


