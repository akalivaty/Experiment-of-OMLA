

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U554 ( .A1(n712), .A2(n711), .ZN(n765) );
  XNOR2_X1 U555 ( .A(n752), .B(n751), .ZN(n753) );
  NOR2_X1 U556 ( .A1(n539), .A2(n538), .ZN(G160) );
  NOR2_X1 U557 ( .A1(n765), .A2(n933), .ZN(n731) );
  NOR2_X1 U558 ( .A1(n964), .A2(n734), .ZN(n736) );
  INV_X1 U559 ( .A(KEYINPUT100), .ZN(n751) );
  INV_X1 U560 ( .A(KEYINPUT101), .ZN(n755) );
  XNOR2_X1 U561 ( .A(n755), .B(KEYINPUT29), .ZN(n756) );
  NOR2_X1 U562 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X2 U563 ( .A1(G2105), .A2(n526), .ZN(n882) );
  NOR2_X1 U564 ( .A1(G651), .A2(n634), .ZN(n640) );
  NOR2_X1 U565 ( .A1(n531), .A2(n530), .ZN(G164) );
  XNOR2_X1 U566 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n521) );
  NOR2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  XNOR2_X2 U568 ( .A(n521), .B(n520), .ZN(n883) );
  NAND2_X1 U569 ( .A1(G138), .A2(n883), .ZN(n523) );
  INV_X1 U570 ( .A(KEYINPUT87), .ZN(n522) );
  XNOR2_X1 U571 ( .A(n523), .B(n522), .ZN(n525) );
  AND2_X1 U572 ( .A1(G2105), .A2(G2104), .ZN(n878) );
  NAND2_X1 U573 ( .A1(n878), .A2(G114), .ZN(n524) );
  NAND2_X1 U574 ( .A1(n525), .A2(n524), .ZN(n531) );
  INV_X1 U575 ( .A(G2104), .ZN(n526) );
  NAND2_X1 U576 ( .A1(G102), .A2(n882), .ZN(n529) );
  NAND2_X1 U577 ( .A1(n526), .A2(G2105), .ZN(n527) );
  XNOR2_X1 U578 ( .A(n527), .B(KEYINPUT65), .ZN(n879) );
  NAND2_X1 U579 ( .A1(G126), .A2(n879), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U581 ( .A1(G101), .A2(n882), .ZN(n533) );
  XOR2_X1 U582 ( .A(KEYINPUT66), .B(KEYINPUT23), .Z(n532) );
  XNOR2_X1 U583 ( .A(n533), .B(n532), .ZN(n535) );
  NAND2_X1 U584 ( .A1(n883), .A2(G137), .ZN(n534) );
  NAND2_X1 U585 ( .A1(n535), .A2(n534), .ZN(n539) );
  NAND2_X1 U586 ( .A1(G113), .A2(n878), .ZN(n537) );
  NAND2_X1 U587 ( .A1(G125), .A2(n879), .ZN(n536) );
  NAND2_X1 U588 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U589 ( .A1(G651), .A2(G543), .ZN(n642) );
  NAND2_X1 U590 ( .A1(G85), .A2(n642), .ZN(n541) );
  XOR2_X1 U591 ( .A(KEYINPUT0), .B(G543), .Z(n634) );
  INV_X1 U592 ( .A(G651), .ZN(n542) );
  NOR2_X1 U593 ( .A1(n634), .A2(n542), .ZN(n645) );
  NAND2_X1 U594 ( .A1(G72), .A2(n645), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n541), .A2(n540), .ZN(n547) );
  NOR2_X1 U596 ( .A1(G543), .A2(n542), .ZN(n543) );
  XOR2_X1 U597 ( .A(KEYINPUT1), .B(n543), .Z(n641) );
  NAND2_X1 U598 ( .A1(G60), .A2(n641), .ZN(n545) );
  NAND2_X1 U599 ( .A1(G47), .A2(n640), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n545), .A2(n544), .ZN(n546) );
  OR2_X1 U601 ( .A1(n547), .A2(n546), .ZN(G290) );
  AND2_X1 U602 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U603 ( .A1(n879), .A2(G123), .ZN(n548) );
  XNOR2_X1 U604 ( .A(n548), .B(KEYINPUT18), .ZN(n550) );
  NAND2_X1 U605 ( .A1(G135), .A2(n883), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n550), .A2(n549), .ZN(n555) );
  NAND2_X1 U607 ( .A1(G99), .A2(n882), .ZN(n552) );
  NAND2_X1 U608 ( .A1(G111), .A2(n878), .ZN(n551) );
  NAND2_X1 U609 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U610 ( .A(KEYINPUT76), .B(n553), .ZN(n554) );
  NOR2_X1 U611 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U612 ( .A(n556), .B(KEYINPUT77), .ZN(n1018) );
  XNOR2_X1 U613 ( .A(G2096), .B(n1018), .ZN(n557) );
  OR2_X1 U614 ( .A1(G2100), .A2(n557), .ZN(G156) );
  INV_X1 U615 ( .A(G132), .ZN(G219) );
  INV_X1 U616 ( .A(G82), .ZN(G220) );
  INV_X1 U617 ( .A(G120), .ZN(G236) );
  INV_X1 U618 ( .A(G69), .ZN(G235) );
  INV_X1 U619 ( .A(G108), .ZN(G238) );
  NAND2_X1 U620 ( .A1(G88), .A2(n642), .ZN(n559) );
  NAND2_X1 U621 ( .A1(G75), .A2(n645), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U623 ( .A1(G62), .A2(n641), .ZN(n561) );
  NAND2_X1 U624 ( .A1(G50), .A2(n640), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U626 ( .A1(n563), .A2(n562), .ZN(G166) );
  NAND2_X1 U627 ( .A1(G64), .A2(n641), .ZN(n565) );
  NAND2_X1 U628 ( .A1(G52), .A2(n640), .ZN(n564) );
  NAND2_X1 U629 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U630 ( .A(KEYINPUT68), .B(n566), .ZN(n571) );
  NAND2_X1 U631 ( .A1(G90), .A2(n642), .ZN(n568) );
  NAND2_X1 U632 ( .A1(G77), .A2(n645), .ZN(n567) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U634 ( .A(KEYINPUT9), .B(n569), .Z(n570) );
  NOR2_X1 U635 ( .A1(n571), .A2(n570), .ZN(G171) );
  NAND2_X1 U636 ( .A1(G63), .A2(n641), .ZN(n573) );
  NAND2_X1 U637 ( .A1(G51), .A2(n640), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(KEYINPUT6), .B(n574), .ZN(n580) );
  NAND2_X1 U640 ( .A1(n642), .A2(G89), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(KEYINPUT4), .ZN(n577) );
  NAND2_X1 U642 ( .A1(G76), .A2(n645), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U644 ( .A(n578), .B(KEYINPUT5), .Z(n579) );
  NOR2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(KEYINPUT7), .B(n581), .Z(n582) );
  XNOR2_X1 U647 ( .A(KEYINPUT74), .B(n582), .ZN(G168) );
  XOR2_X1 U648 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U649 ( .A1(G91), .A2(n642), .ZN(n584) );
  NAND2_X1 U650 ( .A1(G78), .A2(n645), .ZN(n583) );
  NAND2_X1 U651 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U652 ( .A1(G65), .A2(n641), .ZN(n585) );
  XNOR2_X1 U653 ( .A(KEYINPUT69), .B(n585), .ZN(n586) );
  NOR2_X1 U654 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U655 ( .A1(n640), .A2(G53), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n589), .A2(n588), .ZN(G299) );
  NAND2_X1 U657 ( .A1(G7), .A2(G661), .ZN(n590) );
  XNOR2_X1 U658 ( .A(n590), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U659 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n592) );
  INV_X1 U660 ( .A(G223), .ZN(n833) );
  NAND2_X1 U661 ( .A1(G567), .A2(n833), .ZN(n591) );
  XNOR2_X1 U662 ( .A(n592), .B(n591), .ZN(G234) );
  NAND2_X1 U663 ( .A1(n641), .A2(G56), .ZN(n593) );
  XNOR2_X1 U664 ( .A(KEYINPUT14), .B(n593), .ZN(n599) );
  NAND2_X1 U665 ( .A1(n642), .A2(G81), .ZN(n594) );
  XNOR2_X1 U666 ( .A(n594), .B(KEYINPUT12), .ZN(n596) );
  NAND2_X1 U667 ( .A1(G68), .A2(n645), .ZN(n595) );
  NAND2_X1 U668 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U669 ( .A(KEYINPUT13), .B(n597), .ZN(n598) );
  NAND2_X1 U670 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U671 ( .A(n600), .B(KEYINPUT71), .ZN(n602) );
  NAND2_X1 U672 ( .A1(n640), .A2(G43), .ZN(n601) );
  NAND2_X1 U673 ( .A1(n602), .A2(n601), .ZN(n964) );
  INV_X1 U674 ( .A(G860), .ZN(n616) );
  OR2_X1 U675 ( .A1(n964), .A2(n616), .ZN(n603) );
  XNOR2_X1 U676 ( .A(KEYINPUT72), .B(n603), .ZN(G153) );
  INV_X1 U677 ( .A(G171), .ZN(G301) );
  NAND2_X1 U678 ( .A1(G868), .A2(G301), .ZN(n613) );
  NAND2_X1 U679 ( .A1(G54), .A2(n640), .ZN(n610) );
  NAND2_X1 U680 ( .A1(G66), .A2(n641), .ZN(n605) );
  NAND2_X1 U681 ( .A1(G79), .A2(n645), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U683 ( .A1(G92), .A2(n642), .ZN(n606) );
  XNOR2_X1 U684 ( .A(KEYINPUT73), .B(n606), .ZN(n607) );
  NOR2_X1 U685 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U686 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U687 ( .A(n611), .B(KEYINPUT15), .ZN(n955) );
  OR2_X1 U688 ( .A1(n955), .A2(G868), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n613), .A2(n612), .ZN(G284) );
  NAND2_X1 U690 ( .A1(G868), .A2(G286), .ZN(n615) );
  INV_X1 U691 ( .A(G868), .ZN(n659) );
  NAND2_X1 U692 ( .A1(G299), .A2(n659), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n615), .A2(n614), .ZN(G297) );
  NAND2_X1 U694 ( .A1(n616), .A2(G559), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n617), .A2(n955), .ZN(n618) );
  XNOR2_X1 U696 ( .A(n618), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U697 ( .A1(G868), .A2(n964), .ZN(n619) );
  XOR2_X1 U698 ( .A(KEYINPUT75), .B(n619), .Z(n622) );
  NAND2_X1 U699 ( .A1(G868), .A2(n955), .ZN(n620) );
  NOR2_X1 U700 ( .A1(G559), .A2(n620), .ZN(n621) );
  NOR2_X1 U701 ( .A1(n622), .A2(n621), .ZN(G282) );
  NAND2_X1 U702 ( .A1(G61), .A2(n641), .ZN(n624) );
  NAND2_X1 U703 ( .A1(G86), .A2(n642), .ZN(n623) );
  NAND2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n645), .A2(G73), .ZN(n625) );
  XOR2_X1 U706 ( .A(KEYINPUT2), .B(n625), .Z(n626) );
  NOR2_X1 U707 ( .A1(n627), .A2(n626), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n640), .A2(G48), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(G305) );
  NAND2_X1 U710 ( .A1(G49), .A2(n640), .ZN(n631) );
  NAND2_X1 U711 ( .A1(G74), .A2(G651), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U713 ( .A(KEYINPUT80), .B(n632), .ZN(n633) );
  NOR2_X1 U714 ( .A1(n641), .A2(n633), .ZN(n636) );
  NAND2_X1 U715 ( .A1(n634), .A2(G87), .ZN(n635) );
  NAND2_X1 U716 ( .A1(n636), .A2(n635), .ZN(G288) );
  NAND2_X1 U717 ( .A1(G559), .A2(n955), .ZN(n637) );
  XNOR2_X1 U718 ( .A(n637), .B(n964), .ZN(n839) );
  XOR2_X1 U719 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n639) );
  XNOR2_X1 U720 ( .A(KEYINPUT19), .B(KEYINPUT81), .ZN(n638) );
  XNOR2_X1 U721 ( .A(n639), .B(n638), .ZN(n654) );
  NAND2_X1 U722 ( .A1(G55), .A2(n640), .ZN(n650) );
  NAND2_X1 U723 ( .A1(G67), .A2(n641), .ZN(n644) );
  NAND2_X1 U724 ( .A1(G93), .A2(n642), .ZN(n643) );
  NAND2_X1 U725 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U726 ( .A1(n645), .A2(G80), .ZN(n646) );
  XOR2_X1 U727 ( .A(KEYINPUT78), .B(n646), .Z(n647) );
  NOR2_X1 U728 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U729 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U730 ( .A(n651), .B(KEYINPUT79), .Z(n840) );
  XOR2_X1 U731 ( .A(n840), .B(G290), .Z(n652) );
  XNOR2_X1 U732 ( .A(n652), .B(G305), .ZN(n653) );
  XNOR2_X1 U733 ( .A(n654), .B(n653), .ZN(n656) );
  XNOR2_X1 U734 ( .A(G299), .B(G166), .ZN(n655) );
  XNOR2_X1 U735 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U736 ( .A(n657), .B(G288), .ZN(n905) );
  XNOR2_X1 U737 ( .A(n839), .B(n905), .ZN(n658) );
  NAND2_X1 U738 ( .A1(n658), .A2(G868), .ZN(n661) );
  NAND2_X1 U739 ( .A1(n659), .A2(n840), .ZN(n660) );
  NAND2_X1 U740 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n663), .ZN(n665) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(KEYINPUT84), .ZN(n664) );
  XNOR2_X1 U745 ( .A(n665), .B(n664), .ZN(n666) );
  NAND2_X1 U746 ( .A1(G2072), .A2(n666), .ZN(G158) );
  XNOR2_X1 U747 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U748 ( .A1(G235), .A2(G236), .ZN(n667) );
  XNOR2_X1 U749 ( .A(n667), .B(KEYINPUT85), .ZN(n668) );
  NOR2_X1 U750 ( .A1(G238), .A2(n668), .ZN(n669) );
  NAND2_X1 U751 ( .A1(G57), .A2(n669), .ZN(n837) );
  NAND2_X1 U752 ( .A1(G567), .A2(n837), .ZN(n674) );
  NOR2_X1 U753 ( .A1(G220), .A2(G219), .ZN(n670) );
  XOR2_X1 U754 ( .A(KEYINPUT22), .B(n670), .Z(n671) );
  NOR2_X1 U755 ( .A1(G218), .A2(n671), .ZN(n672) );
  NAND2_X1 U756 ( .A1(G96), .A2(n672), .ZN(n838) );
  NAND2_X1 U757 ( .A1(G2106), .A2(n838), .ZN(n673) );
  NAND2_X1 U758 ( .A1(n674), .A2(n673), .ZN(n842) );
  NAND2_X1 U759 ( .A1(G661), .A2(G483), .ZN(n675) );
  NOR2_X1 U760 ( .A1(n842), .A2(n675), .ZN(n836) );
  NAND2_X1 U761 ( .A1(G36), .A2(n836), .ZN(n676) );
  XNOR2_X1 U762 ( .A(n676), .B(KEYINPUT86), .ZN(G176) );
  INV_X1 U763 ( .A(G166), .ZN(G303) );
  NAND2_X1 U764 ( .A1(G40), .A2(G160), .ZN(n677) );
  XNOR2_X1 U765 ( .A(n677), .B(KEYINPUT88), .ZN(n710) );
  NOR2_X1 U766 ( .A1(G164), .A2(G1384), .ZN(n712) );
  NOR2_X1 U767 ( .A1(n710), .A2(n712), .ZN(n828) );
  XNOR2_X1 U768 ( .A(G2067), .B(KEYINPUT37), .ZN(n826) );
  NAND2_X1 U769 ( .A1(n878), .A2(G116), .ZN(n678) );
  XOR2_X1 U770 ( .A(KEYINPUT91), .B(n678), .Z(n680) );
  NAND2_X1 U771 ( .A1(n879), .A2(G128), .ZN(n679) );
  NAND2_X1 U772 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U773 ( .A(KEYINPUT35), .B(n681), .Z(n688) );
  XOR2_X1 U774 ( .A(KEYINPUT34), .B(KEYINPUT90), .Z(n686) );
  NAND2_X1 U775 ( .A1(n882), .A2(G104), .ZN(n682) );
  XOR2_X1 U776 ( .A(KEYINPUT89), .B(n682), .Z(n684) );
  NAND2_X1 U777 ( .A1(n883), .A2(G140), .ZN(n683) );
  NAND2_X1 U778 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U779 ( .A(n686), .B(n685), .Z(n687) );
  NOR2_X1 U780 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U781 ( .A(KEYINPUT36), .B(n689), .ZN(n900) );
  NOR2_X1 U782 ( .A1(n826), .A2(n900), .ZN(n690) );
  XNOR2_X1 U783 ( .A(n690), .B(KEYINPUT92), .ZN(n1013) );
  NAND2_X1 U784 ( .A1(n828), .A2(n1013), .ZN(n824) );
  NAND2_X1 U785 ( .A1(G95), .A2(n882), .ZN(n692) );
  NAND2_X1 U786 ( .A1(G131), .A2(n883), .ZN(n691) );
  NAND2_X1 U787 ( .A1(n692), .A2(n691), .ZN(n696) );
  NAND2_X1 U788 ( .A1(G107), .A2(n878), .ZN(n694) );
  NAND2_X1 U789 ( .A1(G119), .A2(n879), .ZN(n693) );
  NAND2_X1 U790 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U791 ( .A1(n696), .A2(n695), .ZN(n891) );
  INV_X1 U792 ( .A(G1991), .ZN(n817) );
  NOR2_X1 U793 ( .A1(n891), .A2(n817), .ZN(n708) );
  NAND2_X1 U794 ( .A1(G117), .A2(n878), .ZN(n698) );
  NAND2_X1 U795 ( .A1(G129), .A2(n879), .ZN(n697) );
  NAND2_X1 U796 ( .A1(n698), .A2(n697), .ZN(n701) );
  NAND2_X1 U797 ( .A1(n882), .A2(G105), .ZN(n699) );
  XOR2_X1 U798 ( .A(KEYINPUT38), .B(n699), .Z(n700) );
  NOR2_X1 U799 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U800 ( .A(KEYINPUT93), .B(n702), .Z(n704) );
  NAND2_X1 U801 ( .A1(n883), .A2(G141), .ZN(n703) );
  NAND2_X1 U802 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U803 ( .A(KEYINPUT94), .B(n705), .ZN(n893) );
  INV_X1 U804 ( .A(n893), .ZN(n706) );
  INV_X1 U805 ( .A(G1996), .ZN(n933) );
  NOR2_X1 U806 ( .A1(n706), .A2(n933), .ZN(n707) );
  NOR2_X1 U807 ( .A1(n708), .A2(n707), .ZN(n1017) );
  INV_X1 U808 ( .A(n1017), .ZN(n709) );
  NAND2_X1 U809 ( .A1(n709), .A2(n828), .ZN(n816) );
  NAND2_X1 U810 ( .A1(n824), .A2(n816), .ZN(n812) );
  INV_X1 U811 ( .A(n710), .ZN(n711) );
  NOR2_X1 U812 ( .A1(G2084), .A2(n765), .ZN(n713) );
  NAND2_X1 U813 ( .A1(G8), .A2(n713), .ZN(n764) );
  NAND2_X1 U814 ( .A1(G8), .A2(n765), .ZN(n804) );
  NOR2_X1 U815 ( .A1(G1966), .A2(n804), .ZN(n762) );
  NOR2_X1 U816 ( .A1(n762), .A2(n713), .ZN(n714) );
  NAND2_X1 U817 ( .A1(G8), .A2(n714), .ZN(n715) );
  XNOR2_X1 U818 ( .A(KEYINPUT30), .B(n715), .ZN(n716) );
  NOR2_X1 U819 ( .A1(G168), .A2(n716), .ZN(n723) );
  INV_X1 U820 ( .A(n765), .ZN(n717) );
  NOR2_X1 U821 ( .A1(n717), .A2(G1961), .ZN(n718) );
  XNOR2_X1 U822 ( .A(n718), .B(KEYINPUT95), .ZN(n721) );
  XNOR2_X1 U823 ( .A(KEYINPUT25), .B(G2078), .ZN(n935) );
  INV_X1 U824 ( .A(KEYINPUT96), .ZN(n719) );
  XNOR2_X1 U825 ( .A(n719), .B(n765), .ZN(n738) );
  NAND2_X1 U826 ( .A1(n935), .A2(n738), .ZN(n720) );
  NAND2_X1 U827 ( .A1(n721), .A2(n720), .ZN(n758) );
  NOR2_X1 U828 ( .A1(G171), .A2(n758), .ZN(n722) );
  NOR2_X1 U829 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U830 ( .A(KEYINPUT31), .B(n724), .Z(n770) );
  AND2_X1 U831 ( .A1(n738), .A2(G2072), .ZN(n726) );
  XOR2_X1 U832 ( .A(KEYINPUT97), .B(KEYINPUT27), .Z(n725) );
  XNOR2_X1 U833 ( .A(n726), .B(n725), .ZN(n748) );
  INV_X1 U834 ( .A(n738), .ZN(n727) );
  NAND2_X1 U835 ( .A1(n727), .A2(G1956), .ZN(n746) );
  NAND2_X1 U836 ( .A1(n748), .A2(n746), .ZN(n728) );
  NAND2_X1 U837 ( .A1(G299), .A2(n728), .ZN(n729) );
  XOR2_X1 U838 ( .A(KEYINPUT28), .B(n729), .Z(n754) );
  XOR2_X1 U839 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n730) );
  XNOR2_X1 U840 ( .A(n731), .B(n730), .ZN(n733) );
  NAND2_X1 U841 ( .A1(n765), .A2(G1341), .ZN(n732) );
  NAND2_X1 U842 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U843 ( .A1(n955), .A2(n736), .ZN(n735) );
  XNOR2_X1 U844 ( .A(n735), .B(KEYINPUT99), .ZN(n744) );
  NAND2_X1 U845 ( .A1(n955), .A2(n736), .ZN(n742) );
  NAND2_X1 U846 ( .A1(G1348), .A2(n765), .ZN(n737) );
  XNOR2_X1 U847 ( .A(n737), .B(KEYINPUT98), .ZN(n740) );
  NAND2_X1 U848 ( .A1(G2067), .A2(n738), .ZN(n739) );
  NAND2_X1 U849 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U850 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U851 ( .A1(n744), .A2(n743), .ZN(n750) );
  INV_X1 U852 ( .A(G299), .ZN(n745) );
  AND2_X1 U853 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U854 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U855 ( .A1(n750), .A2(n749), .ZN(n752) );
  NOR2_X1 U856 ( .A1(n754), .A2(n753), .ZN(n757) );
  XNOR2_X1 U857 ( .A(n757), .B(n756), .ZN(n760) );
  NAND2_X1 U858 ( .A1(G171), .A2(n758), .ZN(n759) );
  NAND2_X1 U859 ( .A1(n760), .A2(n759), .ZN(n772) );
  AND2_X1 U860 ( .A1(n770), .A2(n772), .ZN(n761) );
  NOR2_X1 U861 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U862 ( .A1(n764), .A2(n763), .ZN(n780) );
  NOR2_X1 U863 ( .A1(G1971), .A2(n804), .ZN(n767) );
  NOR2_X1 U864 ( .A1(G2090), .A2(n765), .ZN(n766) );
  NOR2_X1 U865 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U866 ( .A(n768), .B(KEYINPUT102), .ZN(n769) );
  NAND2_X1 U867 ( .A1(n769), .A2(G303), .ZN(n773) );
  AND2_X1 U868 ( .A1(n770), .A2(n773), .ZN(n771) );
  NAND2_X1 U869 ( .A1(n772), .A2(n771), .ZN(n776) );
  INV_X1 U870 ( .A(n773), .ZN(n774) );
  OR2_X1 U871 ( .A1(n774), .A2(G286), .ZN(n775) );
  AND2_X1 U872 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U873 ( .A1(n777), .A2(G8), .ZN(n778) );
  XNOR2_X1 U874 ( .A(KEYINPUT32), .B(n778), .ZN(n779) );
  NAND2_X1 U875 ( .A1(n780), .A2(n779), .ZN(n803) );
  NOR2_X1 U876 ( .A1(G1976), .A2(G288), .ZN(n781) );
  XOR2_X1 U877 ( .A(KEYINPUT103), .B(n781), .Z(n789) );
  NOR2_X1 U878 ( .A1(G1971), .A2(G303), .ZN(n782) );
  NOR2_X1 U879 ( .A1(n789), .A2(n782), .ZN(n784) );
  INV_X1 U880 ( .A(KEYINPUT33), .ZN(n783) );
  AND2_X1 U881 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U882 ( .A1(n803), .A2(n785), .ZN(n794) );
  INV_X1 U883 ( .A(n804), .ZN(n786) );
  NAND2_X1 U884 ( .A1(G1976), .A2(G288), .ZN(n953) );
  AND2_X1 U885 ( .A1(n786), .A2(n953), .ZN(n787) );
  NOR2_X1 U886 ( .A1(KEYINPUT33), .A2(n787), .ZN(n788) );
  XNOR2_X1 U887 ( .A(G1981), .B(G305), .ZN(n966) );
  NOR2_X1 U888 ( .A1(n788), .A2(n966), .ZN(n792) );
  INV_X1 U889 ( .A(n789), .ZN(n960) );
  NOR2_X1 U890 ( .A1(n804), .A2(n960), .ZN(n790) );
  NAND2_X1 U891 ( .A1(KEYINPUT33), .A2(n790), .ZN(n791) );
  AND2_X1 U892 ( .A1(n792), .A2(n791), .ZN(n793) );
  AND2_X1 U893 ( .A1(n794), .A2(n793), .ZN(n809) );
  NOR2_X1 U894 ( .A1(G2090), .A2(G303), .ZN(n795) );
  XNOR2_X1 U895 ( .A(KEYINPUT104), .B(n795), .ZN(n796) );
  NAND2_X1 U896 ( .A1(n796), .A2(G8), .ZN(n797) );
  XOR2_X1 U897 ( .A(KEYINPUT105), .B(n797), .Z(n801) );
  NOR2_X1 U898 ( .A1(G1981), .A2(G305), .ZN(n798) );
  XOR2_X1 U899 ( .A(n798), .B(KEYINPUT24), .Z(n799) );
  NOR2_X1 U900 ( .A1(n804), .A2(n799), .ZN(n805) );
  INV_X1 U901 ( .A(n805), .ZN(n800) );
  AND2_X1 U902 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U903 ( .A1(n803), .A2(n802), .ZN(n807) );
  OR2_X1 U904 ( .A1(n805), .A2(n804), .ZN(n806) );
  AND2_X1 U905 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U906 ( .A(n810), .B(KEYINPUT106), .ZN(n811) );
  NOR2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n814) );
  XNOR2_X1 U908 ( .A(G1986), .B(G290), .ZN(n959) );
  NAND2_X1 U909 ( .A1(n959), .A2(n828), .ZN(n813) );
  NAND2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n831) );
  NOR2_X1 U911 ( .A1(G1996), .A2(n893), .ZN(n815) );
  XOR2_X1 U912 ( .A(KEYINPUT107), .B(n815), .Z(n1008) );
  INV_X1 U913 ( .A(n816), .ZN(n820) );
  AND2_X1 U914 ( .A1(n817), .A2(n891), .ZN(n1015) );
  NOR2_X1 U915 ( .A1(G1986), .A2(G290), .ZN(n818) );
  NOR2_X1 U916 ( .A1(n1015), .A2(n818), .ZN(n819) );
  NOR2_X1 U917 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U918 ( .A(n821), .B(KEYINPUT108), .ZN(n822) );
  NOR2_X1 U919 ( .A1(n1008), .A2(n822), .ZN(n823) );
  XNOR2_X1 U920 ( .A(n823), .B(KEYINPUT39), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n900), .A2(n826), .ZN(n1019) );
  NAND2_X1 U923 ( .A1(n827), .A2(n1019), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U926 ( .A(KEYINPUT40), .B(n832), .ZN(G329) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U929 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U931 ( .A1(n836), .A2(n835), .ZN(G188) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  NOR2_X1 U934 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  NOR2_X1 U936 ( .A1(n839), .A2(G860), .ZN(n841) );
  XOR2_X1 U937 ( .A(n841), .B(n840), .Z(G145) );
  XNOR2_X1 U938 ( .A(KEYINPUT111), .B(n842), .ZN(G319) );
  XOR2_X1 U939 ( .A(G2100), .B(G2096), .Z(n844) );
  XNOR2_X1 U940 ( .A(KEYINPUT42), .B(G2678), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U942 ( .A(KEYINPUT43), .B(G2090), .Z(n846) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2072), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U945 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U946 ( .A(G2078), .B(G2084), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(G227) );
  XOR2_X1 U948 ( .A(G1976), .B(G1981), .Z(n852) );
  XNOR2_X1 U949 ( .A(G1966), .B(G1971), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U951 ( .A(n853), .B(G2474), .Z(n855) );
  XNOR2_X1 U952 ( .A(G1996), .B(G1991), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U954 ( .A(KEYINPUT41), .B(G1961), .Z(n857) );
  XNOR2_X1 U955 ( .A(G1986), .B(G1956), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n859), .B(n858), .ZN(G229) );
  NAND2_X1 U958 ( .A1(G100), .A2(n882), .ZN(n861) );
  NAND2_X1 U959 ( .A1(G112), .A2(n878), .ZN(n860) );
  NAND2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n867) );
  NAND2_X1 U961 ( .A1(G124), .A2(n879), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n862), .B(KEYINPUT44), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n863), .B(KEYINPUT112), .ZN(n865) );
  NAND2_X1 U964 ( .A1(G136), .A2(n883), .ZN(n864) );
  NAND2_X1 U965 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U966 ( .A1(n867), .A2(n866), .ZN(G162) );
  NAND2_X1 U967 ( .A1(G103), .A2(n882), .ZN(n869) );
  NAND2_X1 U968 ( .A1(G139), .A2(n883), .ZN(n868) );
  NAND2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n875) );
  NAND2_X1 U970 ( .A1(n879), .A2(G127), .ZN(n870) );
  XOR2_X1 U971 ( .A(KEYINPUT113), .B(n870), .Z(n872) );
  NAND2_X1 U972 ( .A1(n878), .A2(G115), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U974 ( .A(KEYINPUT47), .B(n873), .Z(n874) );
  NOR2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n1002) );
  XOR2_X1 U976 ( .A(KEYINPUT115), .B(KEYINPUT114), .Z(n877) );
  XNOR2_X1 U977 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n877), .B(n876), .ZN(n890) );
  NAND2_X1 U979 ( .A1(G118), .A2(n878), .ZN(n881) );
  NAND2_X1 U980 ( .A1(G130), .A2(n879), .ZN(n880) );
  NAND2_X1 U981 ( .A1(n881), .A2(n880), .ZN(n888) );
  NAND2_X1 U982 ( .A1(G106), .A2(n882), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G142), .A2(n883), .ZN(n884) );
  NAND2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U985 ( .A(n886), .B(KEYINPUT45), .Z(n887) );
  NOR2_X1 U986 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U987 ( .A(n890), .B(n889), .Z(n892) );
  XOR2_X1 U988 ( .A(n892), .B(n891), .Z(n895) );
  XNOR2_X1 U989 ( .A(G164), .B(n893), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U991 ( .A(n1018), .B(n896), .ZN(n898) );
  XNOR2_X1 U992 ( .A(G160), .B(G162), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U994 ( .A(n1002), .B(n899), .ZN(n901) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U996 ( .A1(G37), .A2(n902), .ZN(G395) );
  XNOR2_X1 U997 ( .A(G286), .B(KEYINPUT116), .ZN(n904) );
  XNOR2_X1 U998 ( .A(n955), .B(G171), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n907) );
  XOR2_X1 U1000 ( .A(n964), .B(n905), .Z(n906) );
  XNOR2_X1 U1001 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n908), .ZN(G397) );
  XNOR2_X1 U1003 ( .A(G2454), .B(G2443), .ZN(n918) );
  XOR2_X1 U1004 ( .A(G2430), .B(KEYINPUT110), .Z(n910) );
  XNOR2_X1 U1005 ( .A(G2446), .B(KEYINPUT109), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n910), .B(n909), .ZN(n914) );
  XOR2_X1 U1007 ( .A(G2451), .B(G2427), .Z(n912) );
  XNOR2_X1 U1008 ( .A(G1348), .B(G1341), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1010 ( .A(n914), .B(n913), .Z(n916) );
  XNOR2_X1 U1011 ( .A(G2435), .B(G2438), .ZN(n915) );
  XNOR2_X1 U1012 ( .A(n916), .B(n915), .ZN(n917) );
  XNOR2_X1 U1013 ( .A(n918), .B(n917), .ZN(n919) );
  NAND2_X1 U1014 ( .A1(n919), .A2(G14), .ZN(n925) );
  NAND2_X1 U1015 ( .A1(G319), .A2(n925), .ZN(n922) );
  NOR2_X1 U1016 ( .A1(G227), .A2(G229), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(KEYINPUT49), .B(n920), .ZN(n921) );
  NOR2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(n924) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(G57), .ZN(G237) );
  INV_X1 U1023 ( .A(n925), .ZN(G401) );
  XOR2_X1 U1024 ( .A(KEYINPUT124), .B(G29), .Z(n950) );
  XOR2_X1 U1025 ( .A(G34), .B(KEYINPUT123), .Z(n927) );
  XNOR2_X1 U1026 ( .A(G2084), .B(KEYINPUT54), .ZN(n926) );
  XNOR2_X1 U1027 ( .A(n927), .B(n926), .ZN(n947) );
  XOR2_X1 U1028 ( .A(G2090), .B(G35), .Z(n945) );
  XOR2_X1 U1029 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n942) );
  XNOR2_X1 U1030 ( .A(G1991), .B(G25), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(G2067), .B(G26), .ZN(n929) );
  XNOR2_X1 U1032 ( .A(G2072), .B(G33), .ZN(n928) );
  NOR2_X1 U1033 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1034 ( .A(KEYINPUT119), .B(n930), .ZN(n931) );
  NOR2_X1 U1035 ( .A1(n932), .A2(n931), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(G32), .B(n933), .ZN(n934) );
  NAND2_X1 U1037 ( .A1(n934), .A2(G28), .ZN(n938) );
  XOR2_X1 U1038 ( .A(G27), .B(n935), .Z(n936) );
  XNOR2_X1 U1039 ( .A(KEYINPUT120), .B(n936), .ZN(n937) );
  NOR2_X1 U1040 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1041 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1042 ( .A(n942), .B(n941), .ZN(n943) );
  XNOR2_X1 U1043 ( .A(n943), .B(KEYINPUT53), .ZN(n944) );
  NAND2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(KEYINPUT55), .B(n948), .ZN(n949) );
  NAND2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n1032) );
  XNOR2_X1 U1048 ( .A(G16), .B(KEYINPUT56), .ZN(n974) );
  XNOR2_X1 U1049 ( .A(G299), .B(G1956), .ZN(n952) );
  XNOR2_X1 U1050 ( .A(G301), .B(G1961), .ZN(n951) );
  NOR2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n954) );
  NAND2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n963) );
  XNOR2_X1 U1053 ( .A(G166), .B(G1971), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(n955), .B(G1348), .ZN(n956) );
  NAND2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n961) );
  NAND2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n972) );
  XNOR2_X1 U1059 ( .A(n964), .B(G1341), .ZN(n970) );
  XOR2_X1 U1060 ( .A(G168), .B(G1966), .Z(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1062 ( .A(KEYINPUT57), .B(n967), .Z(n968) );
  XNOR2_X1 U1063 ( .A(KEYINPUT125), .B(n968), .ZN(n969) );
  NOR2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n999) );
  INV_X1 U1067 ( .A(G16), .ZN(n997) );
  XNOR2_X1 U1068 ( .A(G1971), .B(G22), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(G23), .B(G1976), .ZN(n975) );
  NOR2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n978) );
  XOR2_X1 U1071 ( .A(G1986), .B(G24), .Z(n977) );
  NAND2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n980) );
  XOR2_X1 U1073 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n979) );
  XNOR2_X1 U1074 ( .A(n980), .B(n979), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(G1966), .B(G21), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(G1961), .B(G5), .ZN(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n994) );
  XOR2_X1 U1079 ( .A(G1348), .B(KEYINPUT59), .Z(n985) );
  XNOR2_X1 U1080 ( .A(G4), .B(n985), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(G20), .B(G1956), .ZN(n986) );
  NOR2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(G1341), .B(G19), .ZN(n989) );
  XNOR2_X1 U1084 ( .A(G1981), .B(G6), .ZN(n988) );
  NOR2_X1 U1085 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1086 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1087 ( .A(KEYINPUT60), .B(n992), .ZN(n993) );
  NOR2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1089 ( .A(KEYINPUT61), .B(n995), .ZN(n996) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1092 ( .A(KEYINPUT127), .B(n1000), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1001), .A2(G11), .ZN(n1030) );
  XNOR2_X1 U1094 ( .A(G2072), .B(n1002), .ZN(n1004) );
  XNOR2_X1 U1095 ( .A(G164), .B(G2078), .ZN(n1003) );
  NAND2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1097 ( .A(n1005), .B(KEYINPUT117), .ZN(n1006) );
  XNOR2_X1 U1098 ( .A(n1006), .B(KEYINPUT50), .ZN(n1011) );
  XOR2_X1 U1099 ( .A(G2090), .B(G162), .Z(n1007) );
  NOR2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1101 ( .A(KEYINPUT51), .B(n1009), .Z(n1010) );
  NAND2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1023) );
  XOR2_X1 U1104 ( .A(G160), .B(G2084), .Z(n1014) );
  NOR2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(KEYINPUT118), .B(n1024), .ZN(n1025) );
  XNOR2_X1 U1111 ( .A(n1025), .B(KEYINPUT52), .ZN(n1026) );
  NOR2_X1 U1112 ( .A1(KEYINPUT55), .A2(n1026), .ZN(n1028) );
  INV_X1 U1113 ( .A(G29), .ZN(n1027) );
  NOR2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1117 ( .A(KEYINPUT62), .B(n1033), .Z(G311) );
  INV_X1 U1118 ( .A(G311), .ZN(G150) );
endmodule

