

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582;

  XNOR2_X2 U320 ( .A(n390), .B(KEYINPUT41), .ZN(n547) );
  NOR2_X1 U321 ( .A1(n384), .A2(n552), .ZN(n385) );
  NOR2_X1 U322 ( .A1(n525), .A2(n544), .ZN(n530) );
  XNOR2_X1 U323 ( .A(n431), .B(KEYINPUT55), .ZN(n432) );
  XNOR2_X1 U324 ( .A(n472), .B(n471), .ZN(n501) );
  XNOR2_X1 U325 ( .A(n411), .B(n410), .ZN(n520) );
  XOR2_X1 U326 ( .A(n396), .B(n395), .Z(n288) );
  XNOR2_X1 U327 ( .A(n412), .B(KEYINPUT116), .ZN(n413) );
  INV_X1 U328 ( .A(n400), .ZN(n401) );
  XNOR2_X1 U329 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U330 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U331 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U332 ( .A(n404), .B(n403), .ZN(n406) );
  XNOR2_X1 U333 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U334 ( .A(n433), .B(n432), .ZN(n448) );
  XNOR2_X1 U335 ( .A(n364), .B(n363), .ZN(n390) );
  AND2_X1 U336 ( .A1(n448), .A2(n523), .ZN(n559) );
  XOR2_X1 U337 ( .A(n447), .B(n446), .Z(n523) );
  XNOR2_X1 U338 ( .A(n449), .B(G190GAT), .ZN(n450) );
  XNOR2_X1 U339 ( .A(n475), .B(KEYINPUT97), .ZN(n476) );
  XNOR2_X1 U340 ( .A(n451), .B(n450), .ZN(G1351GAT) );
  XNOR2_X1 U341 ( .A(n477), .B(n476), .ZN(G1328GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT3), .B(G162GAT), .Z(n290) );
  XNOR2_X1 U343 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n289) );
  XNOR2_X1 U344 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U345 ( .A(G141GAT), .B(n291), .Z(n420) );
  XOR2_X1 U346 ( .A(KEYINPUT83), .B(KEYINPUT85), .Z(n293) );
  XNOR2_X1 U347 ( .A(G85GAT), .B(KEYINPUT84), .ZN(n292) );
  XNOR2_X1 U348 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U349 ( .A(n294), .B(KEYINPUT5), .Z(n296) );
  XOR2_X1 U350 ( .A(G29GAT), .B(G134GAT), .Z(n377) );
  XNOR2_X1 U351 ( .A(G1GAT), .B(n377), .ZN(n295) );
  XNOR2_X1 U352 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U353 ( .A(n420), .B(n297), .ZN(n307) );
  XOR2_X1 U354 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n299) );
  NAND2_X1 U355 ( .A1(G225GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U356 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U357 ( .A(n300), .B(KEYINPUT6), .Z(n305) );
  XOR2_X1 U358 ( .A(G127GAT), .B(KEYINPUT0), .Z(n302) );
  XNOR2_X1 U359 ( .A(G113GAT), .B(KEYINPUT80), .ZN(n301) );
  XNOR2_X1 U360 ( .A(n302), .B(n301), .ZN(n436) );
  XNOR2_X1 U361 ( .A(G120GAT), .B(G148GAT), .ZN(n303) );
  XNOR2_X1 U362 ( .A(n303), .B(G57GAT), .ZN(n358) );
  XNOR2_X1 U363 ( .A(n436), .B(n358), .ZN(n304) );
  XNOR2_X1 U364 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U365 ( .A(n307), .B(n306), .Z(n464) );
  XOR2_X1 U366 ( .A(KEYINPUT86), .B(n464), .Z(n518) );
  XOR2_X1 U367 ( .A(KEYINPUT14), .B(G64GAT), .Z(n309) );
  XNOR2_X1 U368 ( .A(G211GAT), .B(G57GAT), .ZN(n308) );
  XNOR2_X1 U369 ( .A(n309), .B(n308), .ZN(n325) );
  XOR2_X1 U370 ( .A(G8GAT), .B(KEYINPUT77), .Z(n400) );
  XOR2_X1 U371 ( .A(G78GAT), .B(G155GAT), .Z(n311) );
  XNOR2_X1 U372 ( .A(G183GAT), .B(G127GAT), .ZN(n310) );
  XNOR2_X1 U373 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U374 ( .A(n400), .B(n312), .Z(n314) );
  NAND2_X1 U375 ( .A1(G231GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U376 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U377 ( .A(KEYINPUT12), .B(KEYINPUT79), .Z(n316) );
  XNOR2_X1 U378 ( .A(KEYINPUT78), .B(KEYINPUT15), .ZN(n315) );
  XNOR2_X1 U379 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U380 ( .A(n318), .B(n317), .Z(n323) );
  XOR2_X1 U381 ( .A(KEYINPUT69), .B(G1GAT), .Z(n320) );
  XNOR2_X1 U382 ( .A(G15GAT), .B(G22GAT), .ZN(n319) );
  XNOR2_X1 U383 ( .A(n320), .B(n319), .ZN(n331) );
  XNOR2_X1 U384 ( .A(G71GAT), .B(KEYINPUT71), .ZN(n321) );
  XNOR2_X1 U385 ( .A(n321), .B(KEYINPUT13), .ZN(n346) );
  XNOR2_X1 U386 ( .A(n331), .B(n346), .ZN(n322) );
  XNOR2_X1 U387 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U388 ( .A(n325), .B(n324), .ZN(n560) );
  XOR2_X1 U389 ( .A(KEYINPUT70), .B(KEYINPUT66), .Z(n327) );
  XNOR2_X1 U390 ( .A(G197GAT), .B(G8GAT), .ZN(n326) );
  XNOR2_X1 U391 ( .A(n327), .B(n326), .ZN(n343) );
  XNOR2_X1 U392 ( .A(KEYINPUT67), .B(KEYINPUT29), .ZN(n328) );
  XNOR2_X1 U393 ( .A(n328), .B(KEYINPUT68), .ZN(n329) );
  XOR2_X1 U394 ( .A(n329), .B(KEYINPUT30), .Z(n333) );
  XNOR2_X1 U395 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n330) );
  XNOR2_X1 U396 ( .A(n330), .B(KEYINPUT8), .ZN(n378) );
  XNOR2_X1 U397 ( .A(n378), .B(n331), .ZN(n332) );
  XNOR2_X1 U398 ( .A(n333), .B(n332), .ZN(n341) );
  XOR2_X1 U399 ( .A(G141GAT), .B(G113GAT), .Z(n335) );
  XNOR2_X1 U400 ( .A(G169GAT), .B(G50GAT), .ZN(n334) );
  XNOR2_X1 U401 ( .A(n335), .B(n334), .ZN(n337) );
  XOR2_X1 U402 ( .A(G29GAT), .B(G36GAT), .Z(n336) );
  XNOR2_X1 U403 ( .A(n337), .B(n336), .ZN(n339) );
  NAND2_X1 U404 ( .A1(G229GAT), .A2(G233GAT), .ZN(n338) );
  XOR2_X1 U405 ( .A(n343), .B(n342), .Z(n565) );
  INV_X1 U406 ( .A(n565), .ZN(n557) );
  INV_X1 U407 ( .A(n346), .ZN(n344) );
  XOR2_X1 U408 ( .A(G99GAT), .B(G85GAT), .Z(n375) );
  NAND2_X1 U409 ( .A1(n344), .A2(n375), .ZN(n348) );
  INV_X1 U410 ( .A(n375), .ZN(n345) );
  NAND2_X1 U411 ( .A1(n346), .A2(n345), .ZN(n347) );
  NAND2_X1 U412 ( .A1(n348), .A2(n347), .ZN(n350) );
  NAND2_X1 U413 ( .A1(G230GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U414 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U415 ( .A(n351), .B(KEYINPUT33), .ZN(n352) );
  INV_X1 U416 ( .A(n352), .ZN(n356) );
  XOR2_X1 U417 ( .A(G78GAT), .B(G204GAT), .Z(n354) );
  XNOR2_X1 U418 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n353) );
  XNOR2_X1 U419 ( .A(n354), .B(n353), .ZN(n426) );
  XNOR2_X1 U420 ( .A(n426), .B(KEYINPUT72), .ZN(n355) );
  XNOR2_X1 U421 ( .A(n356), .B(n355), .ZN(n364) );
  XNOR2_X1 U422 ( .A(G176GAT), .B(G92GAT), .ZN(n357) );
  XNOR2_X1 U423 ( .A(n357), .B(G64GAT), .ZN(n395) );
  XOR2_X1 U424 ( .A(n358), .B(n395), .Z(n362) );
  XOR2_X1 U425 ( .A(KEYINPUT31), .B(KEYINPUT73), .Z(n360) );
  XNOR2_X1 U426 ( .A(KEYINPUT32), .B(KEYINPUT75), .ZN(n359) );
  XNOR2_X1 U427 ( .A(n360), .B(n359), .ZN(n361) );
  AND2_X1 U428 ( .A1(n557), .A2(n547), .ZN(n365) );
  XNOR2_X1 U429 ( .A(n365), .B(KEYINPUT46), .ZN(n366) );
  NOR2_X1 U430 ( .A1(n560), .A2(n366), .ZN(n367) );
  XNOR2_X1 U431 ( .A(n367), .B(KEYINPUT111), .ZN(n384) );
  XOR2_X1 U432 ( .A(KEYINPUT9), .B(G92GAT), .Z(n369) );
  XNOR2_X1 U433 ( .A(G162GAT), .B(G106GAT), .ZN(n368) );
  XNOR2_X1 U434 ( .A(n369), .B(n368), .ZN(n382) );
  XOR2_X1 U435 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n371) );
  NAND2_X1 U436 ( .A1(G232GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U437 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U438 ( .A(n372), .B(KEYINPUT76), .Z(n374) );
  XOR2_X1 U439 ( .A(G50GAT), .B(G218GAT), .Z(n422) );
  XOR2_X1 U440 ( .A(G36GAT), .B(G190GAT), .Z(n396) );
  XNOR2_X1 U441 ( .A(n422), .B(n396), .ZN(n373) );
  XNOR2_X1 U442 ( .A(n374), .B(n373), .ZN(n376) );
  XOR2_X1 U443 ( .A(n376), .B(n375), .Z(n380) );
  XNOR2_X1 U444 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U445 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n382), .B(n381), .ZN(n386) );
  INV_X1 U447 ( .A(n386), .ZN(n383) );
  INV_X1 U448 ( .A(n383), .ZN(n552) );
  XNOR2_X1 U449 ( .A(n385), .B(KEYINPUT47), .ZN(n393) );
  XOR2_X1 U450 ( .A(n386), .B(KEYINPUT98), .Z(n387) );
  XNOR2_X1 U451 ( .A(n387), .B(KEYINPUT36), .ZN(n580) );
  INV_X1 U452 ( .A(n560), .ZN(n577) );
  NOR2_X1 U453 ( .A1(n580), .A2(n577), .ZN(n388) );
  XOR2_X1 U454 ( .A(KEYINPUT45), .B(n388), .Z(n389) );
  NOR2_X1 U455 ( .A1(n557), .A2(n389), .ZN(n391) );
  BUF_X1 U456 ( .A(n390), .Z(n573) );
  NAND2_X1 U457 ( .A1(n391), .A2(n573), .ZN(n392) );
  NAND2_X1 U458 ( .A1(n393), .A2(n392), .ZN(n394) );
  XNOR2_X1 U459 ( .A(n394), .B(KEYINPUT48), .ZN(n542) );
  NAND2_X1 U460 ( .A1(G226GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n288), .B(n397), .ZN(n398) );
  XOR2_X1 U462 ( .A(n398), .B(KEYINPUT87), .Z(n404) );
  XNOR2_X1 U463 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n399) );
  XNOR2_X1 U464 ( .A(n399), .B(G211GAT), .ZN(n421) );
  XNOR2_X1 U465 ( .A(n421), .B(KEYINPUT88), .ZN(n402) );
  XNOR2_X1 U466 ( .A(G204GAT), .B(G218GAT), .ZN(n405) );
  XNOR2_X1 U467 ( .A(n406), .B(n405), .ZN(n411) );
  XOR2_X1 U468 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n408) );
  XNOR2_X1 U469 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n407) );
  XNOR2_X1 U470 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U471 ( .A(G169GAT), .B(n409), .Z(n447) );
  INV_X1 U472 ( .A(n447), .ZN(n410) );
  NAND2_X1 U473 ( .A1(n542), .A2(n520), .ZN(n414) );
  XOR2_X1 U474 ( .A(KEYINPUT117), .B(KEYINPUT54), .Z(n412) );
  XNOR2_X1 U475 ( .A(n414), .B(n413), .ZN(n415) );
  NOR2_X1 U476 ( .A1(n518), .A2(n415), .ZN(n416) );
  XNOR2_X1 U477 ( .A(n416), .B(KEYINPUT64), .ZN(n563) );
  XOR2_X1 U478 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n418) );
  XNOR2_X1 U479 ( .A(G22GAT), .B(G148GAT), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U481 ( .A(n420), .B(n419), .ZN(n430) );
  XOR2_X1 U482 ( .A(n422), .B(n421), .Z(n424) );
  NAND2_X1 U483 ( .A1(G228GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U485 ( .A(n425), .B(KEYINPUT82), .Z(n428) );
  XNOR2_X1 U486 ( .A(n426), .B(KEYINPUT22), .ZN(n427) );
  XNOR2_X1 U487 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U488 ( .A(n430), .B(n429), .ZN(n458) );
  NAND2_X1 U489 ( .A1(n563), .A2(n458), .ZN(n433) );
  XOR2_X1 U490 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n431) );
  XOR2_X1 U491 ( .A(G99GAT), .B(G43GAT), .Z(n435) );
  NAND2_X1 U492 ( .A1(G227GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n437) );
  XOR2_X1 U494 ( .A(n437), .B(n436), .Z(n445) );
  XOR2_X1 U495 ( .A(KEYINPUT20), .B(KEYINPUT81), .Z(n439) );
  XNOR2_X1 U496 ( .A(G134GAT), .B(G190GAT), .ZN(n438) );
  XNOR2_X1 U497 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U498 ( .A(G120GAT), .B(G71GAT), .Z(n441) );
  XNOR2_X1 U499 ( .A(G15GAT), .B(G176GAT), .ZN(n440) );
  XNOR2_X1 U500 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U501 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U502 ( .A(n445), .B(n444), .ZN(n446) );
  NAND2_X1 U503 ( .A1(n559), .A2(n552), .ZN(n451) );
  XOR2_X1 U504 ( .A(KEYINPUT121), .B(KEYINPUT58), .Z(n449) );
  XNOR2_X1 U505 ( .A(n458), .B(KEYINPUT65), .ZN(n452) );
  XNOR2_X1 U506 ( .A(n452), .B(KEYINPUT28), .ZN(n525) );
  XNOR2_X1 U507 ( .A(n520), .B(KEYINPUT27), .ZN(n457) );
  NAND2_X1 U508 ( .A1(n457), .A2(n518), .ZN(n453) );
  XOR2_X1 U509 ( .A(KEYINPUT89), .B(n453), .Z(n544) );
  INV_X1 U510 ( .A(n523), .ZN(n532) );
  NAND2_X1 U511 ( .A1(n530), .A2(n532), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n454), .B(KEYINPUT90), .ZN(n467) );
  NOR2_X1 U513 ( .A1(n523), .A2(n458), .ZN(n455) );
  XOR2_X1 U514 ( .A(KEYINPUT26), .B(n455), .Z(n456) );
  XNOR2_X1 U515 ( .A(KEYINPUT91), .B(n456), .ZN(n562) );
  NAND2_X1 U516 ( .A1(n457), .A2(n562), .ZN(n463) );
  NAND2_X1 U517 ( .A1(n520), .A2(n523), .ZN(n459) );
  NAND2_X1 U518 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U519 ( .A(n460), .B(KEYINPUT92), .ZN(n461) );
  XOR2_X1 U520 ( .A(KEYINPUT25), .B(n461), .Z(n462) );
  NAND2_X1 U521 ( .A1(n463), .A2(n462), .ZN(n465) );
  NAND2_X1 U522 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U523 ( .A1(n467), .A2(n466), .ZN(n483) );
  NAND2_X1 U524 ( .A1(n577), .A2(n483), .ZN(n468) );
  NOR2_X1 U525 ( .A1(n580), .A2(n468), .ZN(n469) );
  XNOR2_X1 U526 ( .A(KEYINPUT37), .B(n469), .ZN(n517) );
  NAND2_X1 U527 ( .A1(n573), .A2(n557), .ZN(n485) );
  NOR2_X1 U528 ( .A1(n517), .A2(n485), .ZN(n472) );
  XOR2_X1 U529 ( .A(KEYINPUT100), .B(KEYINPUT38), .Z(n470) );
  XNOR2_X1 U530 ( .A(KEYINPUT99), .B(n470), .ZN(n471) );
  NAND2_X1 U531 ( .A1(n518), .A2(n501), .ZN(n477) );
  XOR2_X1 U532 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n474) );
  XNOR2_X1 U533 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n474), .B(n473), .ZN(n475) );
  NAND2_X1 U535 ( .A1(n559), .A2(n547), .ZN(n481) );
  XOR2_X1 U536 ( .A(G176GAT), .B(KEYINPUT56), .Z(n479) );
  XNOR2_X1 U537 ( .A(KEYINPUT57), .B(KEYINPUT120), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(G1349GAT) );
  NOR2_X1 U540 ( .A1(n577), .A2(n552), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(KEYINPUT16), .ZN(n484) );
  NAND2_X1 U542 ( .A1(n484), .A2(n483), .ZN(n506) );
  NOR2_X1 U543 ( .A1(n485), .A2(n506), .ZN(n486) );
  XOR2_X1 U544 ( .A(KEYINPUT93), .B(n486), .Z(n495) );
  NAND2_X1 U545 ( .A1(n518), .A2(n495), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n487), .B(KEYINPUT34), .ZN(n488) );
  XNOR2_X1 U547 ( .A(G1GAT), .B(n488), .ZN(G1324GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n490) );
  NAND2_X1 U549 ( .A1(n495), .A2(n520), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U551 ( .A(G8GAT), .B(n491), .ZN(G1325GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT35), .B(KEYINPUT96), .Z(n493) );
  NAND2_X1 U553 ( .A1(n495), .A2(n523), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G15GAT), .B(n494), .ZN(G1326GAT) );
  NAND2_X1 U556 ( .A1(n495), .A2(n525), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n496), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U558 ( .A(G36GAT), .B(KEYINPUT103), .Z(n498) );
  NAND2_X1 U559 ( .A1(n501), .A2(n520), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(G1329GAT) );
  NAND2_X1 U561 ( .A1(n501), .A2(n523), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n499), .B(KEYINPUT40), .ZN(n500) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n500), .ZN(G1330GAT) );
  NAND2_X1 U564 ( .A1(n501), .A2(n525), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n502), .B(KEYINPUT104), .ZN(n503) );
  XNOR2_X1 U566 ( .A(G50GAT), .B(n503), .ZN(G1331GAT) );
  XNOR2_X1 U567 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n504), .B(KEYINPUT106), .ZN(n505) );
  XOR2_X1 U569 ( .A(KEYINPUT105), .B(n505), .Z(n508) );
  NAND2_X1 U570 ( .A1(n565), .A2(n547), .ZN(n516) );
  NOR2_X1 U571 ( .A1(n506), .A2(n516), .ZN(n512) );
  NAND2_X1 U572 ( .A1(n512), .A2(n518), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(G1332GAT) );
  XOR2_X1 U574 ( .A(G64GAT), .B(KEYINPUT107), .Z(n510) );
  NAND2_X1 U575 ( .A1(n512), .A2(n520), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n512), .A2(n523), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n511), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U580 ( .A1(n512), .A2(n525), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(n515), .ZN(G1335GAT) );
  NOR2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n526) );
  NAND2_X1 U584 ( .A1(n526), .A2(n518), .ZN(n519) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(n519), .ZN(G1336GAT) );
  XOR2_X1 U586 ( .A(G92GAT), .B(KEYINPUT109), .Z(n522) );
  NAND2_X1 U587 ( .A1(n526), .A2(n520), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n526), .A2(n523), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n524), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n528) );
  NAND2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U594 ( .A(G106GAT), .B(n529), .Z(G1339GAT) );
  NAND2_X1 U595 ( .A1(n542), .A2(n530), .ZN(n531) );
  NOR2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n557), .A2(n539), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n533), .B(KEYINPUT112), .ZN(n534) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n534), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n536) );
  NAND2_X1 U601 ( .A1(n539), .A2(n547), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  NAND2_X1 U603 ( .A1(n560), .A2(n539), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n537), .B(KEYINPUT50), .ZN(n538) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U607 ( .A1(n539), .A2(n552), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  NAND2_X1 U609 ( .A1(n542), .A2(n562), .ZN(n543) );
  NOR2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U611 ( .A(KEYINPUT113), .B(n545), .Z(n553) );
  NAND2_X1 U612 ( .A1(n557), .A2(n553), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n546), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n549) );
  NAND2_X1 U615 ( .A1(n553), .A2(n547), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(n550), .ZN(G1345GAT) );
  NAND2_X1 U618 ( .A1(n560), .A2(n553), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n551), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n555) );
  NAND2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(G162GAT), .B(n556), .ZN(G1347GAT) );
  NAND2_X1 U624 ( .A1(n559), .A2(n557), .ZN(n558) );
  XNOR2_X1 U625 ( .A(G169GAT), .B(n558), .ZN(G1348GAT) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U629 ( .A(KEYINPUT122), .B(n564), .ZN(n579) );
  NOR2_X1 U630 ( .A1(n579), .A2(n565), .ZN(n572) );
  XOR2_X1 U631 ( .A(KEYINPUT123), .B(KEYINPUT125), .Z(n567) );
  XNOR2_X1 U632 ( .A(KEYINPUT59), .B(KEYINPUT60), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(n568), .B(KEYINPUT126), .Z(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  XNOR2_X1 U638 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n575) );
  NOR2_X1 U639 ( .A1(n573), .A2(n579), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U641 ( .A(G204GAT), .B(n576), .Z(G1353GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n579), .ZN(n578) );
  XOR2_X1 U643 ( .A(G211GAT), .B(n578), .Z(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(KEYINPUT62), .B(n581), .Z(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

