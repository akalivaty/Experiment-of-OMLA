//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1023,
    new_n1024, new_n1025, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT67), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT1), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT65), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT65), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(G143), .B(G146), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n193), .A2(new_n194), .A3(G128), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(new_n190), .A3(new_n192), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n194), .B1(new_n198), .B2(G128), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n188), .B1(new_n195), .B2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n193), .A2(new_n194), .A3(G128), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(new_n197), .ZN(new_n204));
  OAI211_X1 g018(.A(KEYINPUT67), .B(new_n201), .C1(new_n204), .C2(new_n194), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n200), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT11), .ZN(new_n207));
  INV_X1    g021(.A(G134), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(G137), .ZN(new_n209));
  INV_X1    g023(.A(G137), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT11), .A3(G134), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n208), .A2(G137), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n209), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n215));
  OR2_X1    g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n215), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n210), .A2(G134), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n216), .A2(new_n217), .B1(G131), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n206), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n209), .A2(new_n213), .A3(new_n211), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G131), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n214), .A2(new_n215), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n214), .A2(new_n215), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n194), .A2(KEYINPUT0), .A3(G128), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT0), .B(G128), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n194), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT2), .A2(G113), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT66), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(KEYINPUT2), .A3(G113), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT2), .ZN(new_n237));
  INV_X1    g051(.A(G113), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G116), .B(G119), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n233), .A2(new_n235), .B1(new_n237), .B2(new_n238), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n241), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n243), .A2(KEYINPUT68), .A3(new_n245), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n221), .A2(new_n231), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n206), .A2(new_n220), .B1(new_n226), .B2(new_n230), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(KEYINPUT69), .A3(new_n250), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n201), .B1(new_n204), .B2(new_n194), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n219), .A2(G131), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n257), .B(new_n258), .C1(new_n224), .C2(new_n225), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT30), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n231), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n261), .B1(new_n254), .B2(new_n260), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n246), .ZN(new_n263));
  NOR2_X1   g077(.A1(G237), .A2(G953), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G210), .ZN(new_n265));
  XOR2_X1   g079(.A(new_n265), .B(KEYINPUT27), .Z(new_n266));
  XNOR2_X1  g080(.A(new_n266), .B(KEYINPUT26), .ZN(new_n267));
  INV_X1    g081(.A(G101), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n267), .B(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n256), .A2(new_n263), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT31), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n253), .A2(new_n255), .B1(new_n262), .B2(new_n246), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(KEYINPUT31), .A3(new_n269), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT28), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n251), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n231), .A2(new_n259), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n277), .A2(new_n246), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n278), .B1(new_n253), .B2(new_n255), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n276), .B1(new_n279), .B2(new_n275), .ZN(new_n280));
  INV_X1    g094(.A(new_n269), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n272), .A2(new_n274), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(G472), .A2(G902), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n187), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT31), .B1(new_n273), .B2(new_n269), .ZN(new_n286));
  AND4_X1   g100(.A1(KEYINPUT31), .A2(new_n256), .A3(new_n263), .A4(new_n269), .ZN(new_n287));
  INV_X1    g101(.A(new_n276), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n277), .A2(new_n246), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n254), .A2(KEYINPUT69), .A3(new_n250), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT69), .B1(new_n254), .B2(new_n250), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n288), .B1(new_n292), .B2(KEYINPUT28), .ZN(new_n293));
  OAI22_X1  g107(.A1(new_n286), .A2(new_n287), .B1(new_n293), .B2(new_n269), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(KEYINPUT32), .A3(new_n283), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n285), .A2(new_n295), .A3(KEYINPUT70), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT70), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n297), .B(new_n187), .C1(new_n282), .C2(new_n284), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT71), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n300), .B1(new_n273), .B2(new_n269), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n256), .A2(new_n263), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(KEYINPUT71), .A3(new_n281), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n276), .B(new_n269), .C1(new_n279), .C2(new_n275), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n301), .A2(new_n303), .A3(new_n304), .A4(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n256), .B1(new_n254), .B2(new_n250), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n288), .B1(new_n307), .B2(KEYINPUT28), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n281), .A2(new_n305), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G902), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n306), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G472), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n299), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G217), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n315), .B1(G234), .B2(new_n311), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT25), .ZN(new_n318));
  INV_X1    g132(.A(G953), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(G221), .A3(G234), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(KEYINPUT22), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n321), .B(G137), .ZN(new_n322));
  INV_X1    g136(.A(G140), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G125), .ZN(new_n324));
  INV_X1    g138(.A(G125), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G140), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(KEYINPUT75), .A3(KEYINPUT16), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT16), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n323), .A3(G125), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n324), .A2(new_n326), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n331), .B1(new_n332), .B2(new_n329), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n328), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n196), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n328), .A2(new_n333), .A3(G146), .A4(new_n330), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(G119), .B(G128), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT72), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n338), .B(new_n339), .ZN(new_n340));
  XOR2_X1   g154(.A(KEYINPUT24), .B(G110), .Z(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  OR2_X1    g159(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n346), .A2(G119), .A3(new_n202), .A4(new_n343), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(G110), .A3(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(KEYINPUT74), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n337), .A2(new_n342), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT76), .B1(new_n327), .B2(new_n196), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n327), .A2(KEYINPUT76), .A3(new_n196), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n340), .A2(new_n341), .ZN(new_n353));
  AOI21_X1  g167(.A(G110), .B1(new_n345), .B2(new_n347), .ZN(new_n354));
  OAI221_X1 g168(.A(new_n336), .B1(new_n351), .B2(new_n352), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n322), .B1(new_n350), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n350), .A2(new_n355), .A3(new_n322), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n318), .B1(new_n359), .B2(G902), .ZN(new_n360));
  INV_X1    g174(.A(new_n358), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(new_n356), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(KEYINPUT25), .A3(new_n311), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n317), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n316), .A2(G902), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n364), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(G234), .A2(G237), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n367), .A2(G952), .A3(new_n319), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n367), .A2(G902), .A3(G953), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  XOR2_X1   g185(.A(KEYINPUT21), .B(G898), .Z(new_n372));
  OAI21_X1  g186(.A(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G475), .ZN(new_n374));
  OAI22_X1  g188(.A1(new_n352), .A2(new_n351), .B1(new_n196), .B2(new_n327), .ZN(new_n375));
  AOI21_X1  g189(.A(G143), .B1(new_n264), .B2(G214), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n264), .A2(G143), .A3(G214), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT18), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n377), .B(new_n378), .C1(new_n379), .C2(new_n212), .ZN(new_n380));
  INV_X1    g194(.A(new_n378), .ZN(new_n381));
  OAI21_X1  g195(.A(G131), .B1(new_n381), .B2(new_n376), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n375), .B(new_n380), .C1(new_n379), .C2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT17), .ZN(new_n384));
  OR2_X1    g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n377), .A2(new_n212), .A3(new_n378), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n382), .A2(new_n386), .A3(new_n384), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n335), .A2(new_n385), .A3(new_n336), .A4(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G113), .B(G122), .ZN(new_n389));
  INV_X1    g203(.A(G104), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n389), .B(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n383), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n327), .B(KEYINPUT19), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n196), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n382), .A2(new_n386), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n336), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n391), .B1(new_n383), .B2(new_n397), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n374), .B(new_n311), .C1(new_n393), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT20), .ZN(new_n400));
  INV_X1    g214(.A(new_n398), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n392), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT20), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n402), .A2(new_n403), .A3(new_n374), .A4(new_n311), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n391), .B1(new_n383), .B2(new_n388), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n311), .B1(new_n393), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT92), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI211_X1 g223(.A(KEYINPUT92), .B(new_n311), .C1(new_n393), .C2(new_n406), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(G475), .A3(new_n410), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n405), .A2(new_n411), .ZN(new_n412));
  XOR2_X1   g226(.A(KEYINPUT9), .B(G234), .Z(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(G217), .A3(new_n319), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G143), .ZN(new_n416));
  AOI21_X1  g230(.A(KEYINPUT13), .B1(new_n416), .B2(G128), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(G128), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT94), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT94), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n202), .A2(G143), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n202), .A2(G143), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n420), .B(new_n421), .C1(new_n422), .C2(KEYINPUT13), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(KEYINPUT13), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n419), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G134), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT95), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n422), .A2(new_n418), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n208), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT93), .ZN(new_n430));
  INV_X1    g244(.A(G116), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G122), .ZN(new_n432));
  INV_X1    g246(.A(G122), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G116), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n430), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n434), .A3(new_n430), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(G107), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G107), .ZN(new_n439));
  INV_X1    g253(.A(new_n437), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n439), .B1(new_n440), .B2(new_n435), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT95), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n425), .A2(new_n443), .A3(G134), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n427), .A2(new_n429), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n432), .A2(KEYINPUT14), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT96), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT96), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n432), .A2(new_n448), .A3(KEYINPUT14), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(new_n449), .A3(new_n434), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n432), .A2(KEYINPUT14), .ZN(new_n451));
  OAI21_X1  g265(.A(G107), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n428), .B(new_n208), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n453), .A3(new_n441), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n415), .B1(new_n445), .B2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT98), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n445), .A2(new_n454), .A3(new_n415), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT97), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT97), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n445), .A2(new_n459), .A3(new_n454), .A4(new_n415), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(G902), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT99), .ZN(new_n463));
  INV_X1    g277(.A(G478), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(KEYINPUT15), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n462), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n455), .A2(KEYINPUT98), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT98), .ZN(new_n469));
  AOI211_X1 g283(.A(new_n469), .B(new_n415), .C1(new_n445), .C2(new_n454), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n461), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(new_n463), .A3(new_n311), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n465), .ZN(new_n473));
  AND4_X1   g287(.A1(new_n373), .A2(new_n412), .A3(new_n467), .A4(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(G221), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(new_n413), .B2(new_n311), .ZN(new_n476));
  XOR2_X1   g290(.A(new_n476), .B(KEYINPUT77), .Z(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(G214), .B1(G237), .B2(G902), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n390), .A2(G107), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n439), .A2(G104), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n268), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT3), .B1(new_n390), .B2(G107), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT3), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n439), .A3(G104), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n486), .A2(new_n488), .A3(new_n483), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT78), .B(G101), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n489), .A2(KEYINPUT79), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT79), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n486), .A2(new_n488), .A3(new_n483), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n493), .B1(new_n494), .B2(new_n490), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n485), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n202), .B1(new_n497), .B2(KEYINPUT80), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT80), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n197), .A2(new_n499), .A3(KEYINPUT1), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n194), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n496), .B1(new_n195), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT10), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n492), .A2(new_n495), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n489), .A2(new_n268), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(KEYINPUT4), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT4), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n229), .B1(new_n508), .B2(new_n505), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n502), .A2(new_n503), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n226), .ZN(new_n511));
  AOI211_X1 g325(.A(new_n503), .B(new_n485), .C1(new_n492), .C2(new_n495), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT81), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n513), .A3(new_n206), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n513), .B1(new_n512), .B2(new_n206), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n510), .B(new_n511), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(G110), .B(G140), .ZN(new_n518));
  INV_X1    g332(.A(G227), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(G953), .ZN(new_n520));
  XOR2_X1   g334(.A(new_n518), .B(new_n520), .Z(new_n521));
  INV_X1    g335(.A(new_n485), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n504), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n195), .A2(new_n199), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n511), .B1(new_n525), .B2(new_n502), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT12), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(KEYINPUT82), .A3(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n501), .A2(new_n195), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n523), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n496), .A2(new_n257), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n226), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n517), .A2(new_n521), .A3(new_n528), .A4(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT83), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n521), .ZN(new_n538));
  INV_X1    g352(.A(new_n517), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n512), .A2(new_n206), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT81), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n514), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n511), .B1(new_n542), .B2(new_n510), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n538), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n533), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n526), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n527), .A2(KEYINPUT82), .ZN(new_n547));
  AOI211_X1 g361(.A(new_n511), .B(new_n547), .C1(new_n525), .C2(new_n502), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n549), .A2(KEYINPUT83), .A3(new_n517), .A4(new_n521), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n537), .A2(new_n544), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G469), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n552), .A3(new_n311), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n521), .B1(new_n539), .B2(new_n543), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n549), .A2(new_n517), .A3(new_n538), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(G469), .B1(new_n556), .B2(G902), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n482), .B1(new_n553), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n229), .A2(G125), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT85), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT85), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n229), .A2(new_n561), .A3(G125), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n524), .A2(new_n325), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT87), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT86), .B(G224), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n319), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT87), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n560), .A2(new_n563), .A3(new_n569), .A4(new_n562), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n565), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n568), .B1(new_n565), .B2(new_n570), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT6), .ZN(new_n575));
  XOR2_X1   g389(.A(G110), .B(G122), .Z(new_n576));
  NAND3_X1  g390(.A1(new_n494), .A2(new_n508), .A3(G101), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n244), .A2(new_n241), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n236), .A2(new_n239), .A3(new_n241), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n508), .B1(new_n492), .B2(new_n495), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n580), .B1(new_n581), .B2(new_n506), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n431), .A2(G119), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT5), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n238), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(G119), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(G116), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n431), .A2(G119), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(new_n588), .A3(KEYINPUT5), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n244), .A2(new_n241), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT79), .B1(new_n489), .B2(new_n491), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n494), .A2(new_n493), .A3(new_n490), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n522), .B(new_n590), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT84), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n582), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n580), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n507), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT84), .B1(new_n598), .B2(new_n593), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n576), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n582), .A2(new_n594), .A3(new_n576), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n575), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n576), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n595), .B1(new_n582), .B2(new_n594), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n598), .A2(KEYINPUT84), .A3(new_n593), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n607), .A2(KEYINPUT6), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n574), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n567), .A2(KEYINPUT7), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n564), .B(new_n610), .ZN(new_n611));
  OR2_X1    g425(.A1(new_n589), .A2(KEYINPUT89), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n589), .A2(KEYINPUT89), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n585), .A3(new_n613), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n496), .A2(new_n245), .A3(new_n614), .ZN(new_n615));
  OR3_X1    g429(.A1(new_n496), .A2(KEYINPUT90), .A3(new_n590), .ZN(new_n616));
  OAI21_X1  g430(.A(KEYINPUT90), .B1(new_n496), .B2(new_n590), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT88), .B(KEYINPUT8), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n576), .B(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n611), .B(new_n602), .C1(new_n618), .C2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n311), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(G210), .B1(G237), .B2(G902), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(KEYINPUT91), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n609), .A2(new_n624), .A3(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(KEYINPUT6), .B1(new_n607), .B2(new_n601), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n600), .A2(new_n575), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n573), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n626), .B1(new_n631), .B2(new_n623), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n474), .A2(new_n558), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n314), .A2(new_n366), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(new_n490), .ZN(G3));
  AOI21_X1  g450(.A(new_n478), .B1(new_n553), .B2(new_n557), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n366), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(G472), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n294), .B2(new_n311), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT100), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n644), .B1(new_n282), .B2(new_n284), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n643), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n457), .B1(new_n455), .B2(KEYINPUT102), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n445), .A2(new_n648), .A3(new_n454), .A4(new_n415), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT33), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT33), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n461), .B(new_n652), .C1(new_n468), .C2(new_n470), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n654), .A2(G478), .A3(new_n311), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n471), .A2(new_n311), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n464), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n405), .A2(new_n411), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n373), .A2(new_n479), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n625), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n625), .A2(new_n662), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n609), .A2(new_n624), .A3(new_n663), .A4(new_n664), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n662), .B(new_n625), .C1(new_n631), .C2(new_n623), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n660), .A2(new_n661), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n640), .A2(new_n646), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT34), .B(G104), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G6));
  INV_X1    g485(.A(KEYINPUT103), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n411), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n409), .A2(KEYINPUT103), .A3(G475), .A4(new_n410), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n673), .A2(new_n405), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n661), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n675), .A2(new_n676), .A3(new_n666), .A4(new_n665), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n473), .A2(new_n467), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n640), .A2(new_n680), .A3(new_n646), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT35), .B(G107), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G9));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n684));
  INV_X1    g498(.A(new_n322), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(KEYINPUT36), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n350), .A2(new_n688), .A3(new_n355), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n688), .B1(new_n350), .B2(new_n355), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n687), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n350), .A2(new_n355), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT104), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n686), .A3(new_n689), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n365), .ZN(new_n697));
  OAI21_X1  g511(.A(KEYINPUT105), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n692), .A2(new_n695), .A3(new_n699), .A4(new_n365), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n684), .B1(new_n701), .B2(new_n364), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n360), .A2(new_n363), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n316), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n704), .A2(KEYINPUT106), .A3(new_n698), .A4(new_n700), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n634), .A2(new_n646), .A3(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(new_n707), .B(KEYINPUT37), .Z(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G110), .ZN(G12));
  INV_X1    g523(.A(G900), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n370), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n369), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n675), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n679), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n665), .A2(new_n666), .A3(new_n479), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n638), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n314), .A2(new_n706), .A3(new_n714), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G128), .ZN(G30));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n307), .A2(new_n269), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(G902), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n302), .A2(new_n269), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n641), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n299), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n633), .B(KEYINPUT38), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n412), .B1(new_n473), .B2(new_n467), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n701), .A2(new_n364), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n480), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n725), .A2(new_n726), .A3(new_n727), .A4(new_n730), .ZN(new_n731));
  XOR2_X1   g545(.A(new_n712), .B(KEYINPUT39), .Z(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n637), .A2(new_n733), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n734), .A2(KEYINPUT108), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(KEYINPUT108), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n719), .A2(new_n731), .B1(new_n737), .B2(KEYINPUT40), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n738), .B1(KEYINPUT40), .B2(new_n737), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n731), .A2(new_n719), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n416), .ZN(G45));
  INV_X1    g556(.A(new_n712), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n660), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n314), .A2(new_n706), .A3(new_n716), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G146), .ZN(G48));
  NAND2_X1  g560(.A1(new_n551), .A2(new_n311), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(G469), .ZN(new_n748));
  INV_X1    g562(.A(new_n476), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n749), .A3(new_n553), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n314), .A2(new_n366), .A3(new_n668), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(KEYINPUT41), .B(G113), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(G15));
  NAND4_X1  g568(.A1(new_n314), .A2(new_n366), .A3(new_n680), .A4(new_n751), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G116), .ZN(G18));
  NOR2_X1   g570(.A1(new_n750), .A2(new_n715), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n314), .A2(new_n474), .A3(new_n706), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT109), .ZN(new_n759));
  AOI22_X1  g573(.A1(new_n299), .A2(new_n313), .B1(new_n702), .B2(new_n705), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n760), .A2(new_n761), .A3(new_n474), .A4(new_n757), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G119), .ZN(G21));
  XNOR2_X1  g578(.A(new_n283), .B(KEYINPUT110), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n308), .A2(new_n269), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n272), .A2(new_n274), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n639), .A2(new_n769), .A3(new_n642), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n678), .A2(new_n659), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n715), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n770), .A2(new_n373), .A3(new_n751), .A4(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G122), .ZN(G24));
  NOR3_X1   g588(.A1(new_n769), .A2(new_n728), .A3(new_n642), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n757), .A2(new_n744), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G125), .ZN(G27));
  AOI22_X1  g591(.A1(new_n296), .A2(new_n298), .B1(G472), .B2(new_n312), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n628), .A2(new_n632), .A3(new_n479), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n553), .A2(new_n557), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(new_n749), .A3(new_n780), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n778), .A2(new_n639), .A3(new_n781), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n660), .A2(KEYINPUT42), .A3(new_n743), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n779), .A2(new_n749), .A3(new_n780), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n313), .A2(new_n285), .A3(new_n295), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(new_n366), .A3(new_n744), .A4(new_n785), .ZN(new_n786));
  AOI22_X1  g600(.A1(new_n782), .A2(new_n783), .B1(new_n786), .B2(KEYINPUT42), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT111), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(new_n212), .ZN(G33));
  NAND4_X1  g603(.A1(new_n314), .A2(new_n366), .A3(new_n714), .A4(new_n784), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G134), .ZN(G36));
  OAI21_X1  g605(.A(new_n510), .B1(new_n515), .B2(new_n516), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n226), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n538), .B1(new_n793), .B2(new_n517), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n517), .A2(new_n538), .A3(new_n528), .A4(new_n534), .ZN(new_n795));
  OAI21_X1  g609(.A(KEYINPUT45), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n554), .A2(new_n797), .A3(new_n555), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n796), .A2(new_n798), .A3(G469), .ZN(new_n799));
  NAND2_X1  g613(.A1(G469), .A2(G902), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n799), .A2(KEYINPUT46), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT46), .B1(new_n799), .B2(new_n800), .ZN(new_n802));
  INV_X1    g616(.A(new_n553), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n804), .A2(new_n476), .A3(new_n732), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n658), .A2(new_n412), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT43), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(KEYINPUT112), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n659), .B1(new_n655), .B2(new_n657), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n809), .B1(new_n810), .B2(KEYINPUT43), .ZN(new_n811));
  AOI211_X1 g625(.A(new_n464), .B(G902), .C1(new_n651), .C2(new_n653), .ZN(new_n812));
  INV_X1    g626(.A(new_n657), .ZN(new_n813));
  OAI211_X1 g627(.A(KEYINPUT43), .B(new_n412), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n810), .A2(KEYINPUT113), .A3(KEYINPUT43), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n808), .A2(new_n811), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n818), .A2(new_n646), .A3(new_n728), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT112), .B1(new_n806), .B2(new_n807), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n810), .A2(new_n809), .A3(KEYINPUT43), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n814), .A2(new_n815), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT113), .B1(new_n810), .B2(KEYINPUT43), .ZN(new_n823));
  OAI22_X1  g637(.A1(new_n820), .A2(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n646), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(KEYINPUT44), .A3(new_n825), .A4(new_n729), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n779), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n827), .A2(KEYINPUT114), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(KEYINPUT114), .ZN(new_n829));
  OAI221_X1 g643(.A(new_n805), .B1(KEYINPUT44), .B2(new_n819), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(G137), .ZN(G39));
  NOR3_X1   g645(.A1(new_n804), .A2(KEYINPUT47), .A3(new_n476), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT47), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n799), .A2(new_n800), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT46), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n799), .A2(KEYINPUT46), .A3(new_n800), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n836), .A2(new_n553), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n833), .B1(new_n838), .B2(new_n749), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n832), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n314), .A2(new_n366), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n744), .A3(new_n779), .A4(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(G140), .ZN(G42));
  NAND2_X1  g657(.A1(new_n780), .A2(new_n728), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n299), .B2(new_n724), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n715), .A2(new_n771), .A3(new_n476), .A4(new_n743), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT115), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n723), .B1(new_n296), .B2(new_n298), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n665), .A2(new_n666), .A3(new_n479), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n749), .A3(new_n712), .A4(new_n727), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT115), .ZN(new_n851));
  NOR4_X1   g665(.A1(new_n848), .A2(new_n850), .A3(new_n851), .A4(new_n844), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n717), .A2(new_n745), .A3(new_n776), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT52), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n717), .A2(new_n745), .A3(new_n776), .ZN(new_n856));
  INV_X1    g670(.A(new_n844), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n725), .A2(new_n846), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n851), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n845), .A2(KEYINPUT115), .A3(new_n846), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT52), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n856), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n855), .A2(new_n863), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n752), .A2(new_n755), .A3(new_n773), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n678), .A2(new_n412), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n661), .B1(new_n660), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n640), .A2(new_n646), .A3(new_n633), .A4(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n635), .A2(new_n868), .A3(new_n707), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n763), .A2(new_n865), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n784), .A2(new_n744), .A3(new_n775), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n706), .A2(new_n679), .A3(new_n637), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n628), .A2(new_n632), .A3(new_n479), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n713), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n314), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n787), .A2(new_n790), .A3(new_n872), .A4(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n864), .A2(KEYINPUT53), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n855), .A2(new_n863), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n786), .A2(KEYINPUT42), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n314), .A2(new_n366), .A3(new_n784), .A4(new_n783), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n882), .A2(new_n883), .A3(new_n790), .A4(new_n876), .ZN(new_n884));
  INV_X1    g698(.A(new_n872), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n869), .B1(new_n762), .B2(new_n759), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(new_n887), .A3(new_n865), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n880), .B1(new_n881), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT116), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n879), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  OAI211_X1 g705(.A(KEYINPUT116), .B(new_n880), .C1(new_n881), .C2(new_n888), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(KEYINPUT54), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n717), .A2(new_n776), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT52), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n864), .A2(KEYINPUT53), .A3(new_n878), .A4(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n896), .A2(new_n897), .A3(new_n889), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT117), .B1(new_n832), .B2(new_n839), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT47), .B1(new_n804), .B2(new_n476), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT117), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n838), .A2(new_n833), .A3(new_n749), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n748), .A2(new_n478), .A3(new_n553), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n899), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT118), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n769), .A2(new_n642), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n366), .ZN(new_n908));
  NOR4_X1   g722(.A1(new_n818), .A2(new_n369), .A3(new_n908), .A4(new_n874), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n905), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n906), .B1(new_n905), .B2(new_n909), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n818), .A2(new_n369), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n750), .A2(new_n874), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n913), .A2(KEYINPUT119), .A3(new_n775), .A4(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n824), .A2(new_n368), .A3(new_n775), .A4(new_n914), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT119), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n639), .A2(new_n369), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n848), .A2(new_n914), .A3(new_n412), .A4(new_n920), .ZN(new_n921));
  OR3_X1    g735(.A1(new_n921), .A2(KEYINPUT120), .A3(new_n658), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT120), .B1(new_n921), .B2(new_n658), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR4_X1   g738(.A1(new_n818), .A2(new_n369), .A3(new_n908), .A4(new_n750), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n726), .A2(new_n479), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT50), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n824), .A2(new_n368), .A3(new_n751), .A4(new_n770), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT50), .ZN(new_n929));
  INV_X1    g743(.A(new_n926), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n919), .B(new_n924), .C1(new_n927), .C2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT121), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n925), .A2(KEYINPUT50), .A3(new_n926), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n929), .B1(new_n928), .B2(new_n930), .ZN(new_n935));
  AOI22_X1  g749(.A1(new_n934), .A2(new_n935), .B1(new_n922), .B2(new_n923), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT121), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n936), .A2(new_n937), .A3(new_n919), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n912), .A2(new_n933), .A3(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT51), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(G952), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n848), .A2(new_n914), .A3(new_n920), .ZN(new_n943));
  INV_X1    g757(.A(new_n660), .ZN(new_n944));
  AOI211_X1 g758(.A(new_n942), .B(G953), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n785), .A2(new_n366), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n913), .A2(new_n946), .A3(new_n914), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n947), .A2(KEYINPUT48), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n947), .A2(KEYINPUT48), .ZN(new_n949));
  OAI221_X1 g763(.A(new_n945), .B1(new_n715), .B2(new_n928), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n904), .B1(new_n832), .B2(new_n839), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n940), .B1(new_n951), .B2(new_n909), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n936), .A2(new_n919), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT122), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n936), .A2(new_n952), .A3(KEYINPUT122), .A4(new_n919), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n950), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n893), .A2(new_n898), .A3(new_n941), .A4(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT123), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n942), .A2(new_n319), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n941), .A2(new_n957), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n962), .A2(KEYINPUT123), .A3(new_n893), .A4(new_n898), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n960), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n748), .A2(new_n553), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n965), .A2(KEYINPUT49), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(KEYINPUT49), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n966), .A2(new_n967), .A3(new_n639), .ZN(new_n968));
  INV_X1    g782(.A(new_n726), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n806), .A2(new_n482), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n968), .A2(new_n969), .A3(new_n848), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n964), .A2(new_n971), .ZN(G75));
  NAND3_X1  g786(.A1(new_n629), .A2(new_n630), .A3(new_n573), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n609), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT55), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT124), .ZN(new_n977));
  INV_X1    g791(.A(G210), .ZN(new_n978));
  AOI211_X1 g792(.A(new_n978), .B(new_n311), .C1(new_n896), .C2(new_n889), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n977), .B1(new_n979), .B2(KEYINPUT56), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n896), .A2(new_n889), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n981), .A2(G210), .A3(G902), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT56), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n982), .A2(KEYINPUT124), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n976), .B1(new_n980), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n319), .A2(G952), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n982), .A2(new_n983), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n975), .B1(new_n987), .B2(new_n977), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n985), .A2(new_n986), .A3(new_n988), .ZN(G51));
  INV_X1    g803(.A(new_n898), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n897), .B1(new_n896), .B2(new_n889), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n800), .B(KEYINPUT57), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n551), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n311), .B1(new_n896), .B2(new_n889), .ZN(new_n995));
  INV_X1    g809(.A(new_n799), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n986), .B1(new_n994), .B2(new_n997), .ZN(G54));
  NAND3_X1  g812(.A1(new_n995), .A2(KEYINPUT58), .A3(G475), .ZN(new_n999));
  INV_X1    g813(.A(new_n402), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n999), .A2(new_n1000), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n1001), .A2(new_n1002), .A3(new_n986), .ZN(G60));
  NAND2_X1  g817(.A1(G478), .A2(G902), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT59), .Z(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n654), .B(new_n1006), .C1(new_n990), .C2(new_n991), .ZN(new_n1007));
  INV_X1    g821(.A(new_n986), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1005), .B1(new_n893), .B2(new_n898), .ZN(new_n1009));
  OAI211_X1 g823(.A(new_n1007), .B(new_n1008), .C1(new_n1009), .C2(new_n654), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(G63));
  NAND2_X1  g825(.A1(G217), .A2(G902), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT125), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1013), .B(KEYINPUT60), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n981), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1008), .B1(new_n1015), .B2(new_n696), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT61), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n362), .B(KEYINPUT126), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1018), .B1(new_n981), .B2(new_n1014), .ZN(new_n1019));
  OR3_X1    g833(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1017), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(new_n1021), .ZN(G66));
  AOI21_X1  g836(.A(new_n319), .B1(new_n372), .B2(new_n566), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1023), .B1(new_n871), .B2(new_n319), .ZN(new_n1024));
  OAI211_X1 g838(.A(new_n629), .B(new_n630), .C1(G898), .C2(new_n319), .ZN(new_n1025));
  XOR2_X1   g839(.A(new_n1024), .B(new_n1025), .Z(G69));
  XOR2_X1   g840(.A(new_n262), .B(new_n394), .Z(new_n1027));
  OAI21_X1  g841(.A(G953), .B1(new_n1027), .B2(new_n519), .ZN(new_n1028));
  AOI211_X1 g842(.A(new_n710), .B(new_n1028), .C1(new_n519), .C2(new_n1027), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT62), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1030), .B1(new_n741), .B2(new_n854), .ZN(new_n1031));
  OAI211_X1 g845(.A(KEYINPUT62), .B(new_n856), .C1(new_n739), .C2(new_n740), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n734), .A2(new_n874), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n660), .A2(new_n866), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n314), .A2(new_n1034), .A3(new_n366), .A4(new_n1035), .ZN(new_n1036));
  NAND4_X1  g850(.A1(new_n1033), .A2(new_n830), .A3(new_n842), .A4(new_n1036), .ZN(new_n1037));
  AOI21_X1  g851(.A(G953), .B1(new_n1037), .B2(new_n1027), .ZN(new_n1038));
  AND2_X1   g852(.A1(new_n946), .A2(new_n772), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1039), .A2(new_n805), .ZN(new_n1040));
  AND3_X1   g854(.A1(new_n787), .A2(new_n1040), .A3(new_n790), .ZN(new_n1041));
  NAND4_X1  g855(.A1(new_n830), .A2(new_n842), .A3(new_n1041), .A4(new_n856), .ZN(new_n1042));
  OR2_X1    g856(.A1(new_n1042), .A2(new_n1027), .ZN(new_n1043));
  AOI21_X1  g857(.A(new_n1029), .B1(new_n1038), .B2(new_n1043), .ZN(G72));
  NAND2_X1  g858(.A1(G472), .A2(G902), .ZN(new_n1045));
  XOR2_X1   g859(.A(new_n1045), .B(KEYINPUT63), .Z(new_n1046));
  OAI21_X1  g860(.A(new_n1046), .B1(new_n1037), .B2(new_n871), .ZN(new_n1047));
  INV_X1    g861(.A(new_n722), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n986), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1046), .B1(new_n1042), .B2(new_n871), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1050), .A2(KEYINPUT127), .ZN(new_n1051));
  INV_X1    g865(.A(KEYINPUT127), .ZN(new_n1052));
  OAI211_X1 g866(.A(new_n1052), .B(new_n1046), .C1(new_n1042), .C2(new_n871), .ZN(new_n1053));
  NAND4_X1  g867(.A1(new_n1051), .A2(new_n281), .A3(new_n273), .A4(new_n1053), .ZN(new_n1054));
  NAND3_X1  g868(.A1(new_n301), .A2(new_n303), .A3(new_n270), .ZN(new_n1055));
  NAND4_X1  g869(.A1(new_n891), .A2(new_n892), .A3(new_n1046), .A4(new_n1055), .ZN(new_n1056));
  AND3_X1   g870(.A1(new_n1049), .A2(new_n1054), .A3(new_n1056), .ZN(G57));
endmodule


