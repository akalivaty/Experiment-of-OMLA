//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT0), .ZN(new_n206));
  XNOR2_X1  g0006(.A(KEYINPUT66), .B(G244), .ZN(new_n207));
  INV_X1    g0007(.A(G77), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G116), .A2(G270), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n203), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT64), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g0018(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT65), .Z(new_n226));
  OAI221_X1 g0026(.A(new_n206), .B1(KEYINPUT1), .B2(new_n215), .C1(new_n224), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n215), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n231), .B(new_n232), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(new_n241), .B(KEYINPUT68), .Z(new_n242));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NOR2_X1   g0046(.A1(G20), .A2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G150), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT8), .B(G58), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n222), .A2(G33), .ZN(new_n250));
  NOR3_X1   g0050(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n251));
  OAI221_X1 g0051(.A(new_n248), .B1(new_n249), .B2(new_n250), .C1(new_n251), .C2(new_n222), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n218), .A2(new_n219), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G50), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n252), .A2(new_n254), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n254), .A2(new_n258), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n260), .B(G50), .C1(G1), .C2(new_n222), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OR2_X1    g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(G222), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n266), .A2(G223), .A3(G1698), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n268), .B(new_n269), .C1(new_n208), .C2(new_n266), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  AND3_X1   g0071(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n272));
  AOI21_X1  g0072(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  INV_X1    g0077(.A(G45), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(G1), .A2(G13), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n256), .A2(new_n279), .B1(new_n280), .B2(new_n271), .ZN(new_n281));
  INV_X1    g0081(.A(G274), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n282), .B1(new_n280), .B2(new_n271), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n281), .A2(G226), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n276), .A2(new_n286), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n263), .A2(KEYINPUT9), .B1(new_n287), .B2(G200), .ZN(new_n288));
  INV_X1    g0088(.A(new_n287), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT9), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n289), .A2(G190), .B1(new_n262), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT10), .ZN(new_n293));
  INV_X1    g0093(.A(G169), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n263), .B1(new_n294), .B2(new_n287), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n295), .B1(G179), .B2(new_n287), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n283), .A2(new_n285), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n280), .A2(new_n271), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n284), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n298), .B1(new_n300), .B2(new_n207), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n230), .A2(G1698), .ZN(new_n302));
  INV_X1    g0102(.A(G238), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(new_n267), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n266), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G107), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(new_n266), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT69), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n274), .B1(new_n307), .B2(new_n308), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n301), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G179), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n254), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT15), .B(G87), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT70), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(new_n316), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n319), .A2(new_n250), .ZN(new_n320));
  INV_X1    g0120(.A(new_n249), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n321), .A2(new_n247), .B1(G20), .B2(G77), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n314), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  XOR2_X1   g0123(.A(new_n257), .B(KEYINPUT71), .Z(new_n324));
  NOR2_X1   g0124(.A1(new_n324), .A2(new_n254), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n208), .B1(new_n256), .B2(G20), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n257), .B(KEYINPUT71), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(G77), .B2(new_n328), .ZN(new_n329));
  OAI221_X1 g0129(.A(new_n313), .B1(G169), .B2(new_n311), .C1(new_n323), .C2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n323), .A2(new_n329), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n311), .A2(G190), .ZN(new_n332));
  INV_X1    g0132(.A(G200), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n331), .B(new_n332), .C1(new_n333), .C2(new_n311), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n297), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT16), .ZN(new_n337));
  INV_X1    g0137(.A(G68), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n264), .A2(new_n222), .A3(new_n265), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT7), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AND2_X1   g0141(.A1(KEYINPUT3), .A2(G33), .ZN(new_n342));
  NOR2_X1   g0142(.A1(KEYINPUT3), .A2(G33), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(KEYINPUT7), .A3(new_n222), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n338), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G58), .A2(G68), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT77), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G58), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n338), .ZN(new_n351));
  NAND3_X1  g0151(.A1(KEYINPUT77), .A2(G58), .A3(G68), .ZN(new_n352));
  AND3_X1   g0152(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G159), .ZN(new_n354));
  INV_X1    g0154(.A(new_n247), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n353), .A2(new_n222), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n337), .B1(new_n346), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT7), .B1(new_n344), .B2(new_n222), .ZN(new_n358));
  NOR4_X1   g0158(.A1(new_n342), .A2(new_n343), .A3(new_n340), .A4(G20), .ZN(new_n359));
  OAI21_X1  g0159(.A(G68), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n349), .B(new_n352), .C1(G58), .C2(G68), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n361), .A2(G20), .B1(G159), .B2(new_n247), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(new_n362), .A3(KEYINPUT16), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n357), .A2(new_n363), .A3(new_n254), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n249), .B1(new_n256), .B2(G20), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n260), .A2(new_n365), .B1(new_n258), .B2(new_n249), .ZN(new_n366));
  NAND2_X1  g0166(.A1(G33), .A2(G87), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT78), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n367), .B(new_n368), .ZN(new_n369));
  OR2_X1    g0169(.A1(G223), .A2(G1698), .ZN(new_n370));
  INV_X1    g0170(.A(G226), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G1698), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n370), .B(new_n372), .C1(new_n342), .C2(new_n343), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n275), .ZN(new_n375));
  INV_X1    g0175(.A(G190), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n281), .A2(G232), .B1(new_n283), .B2(new_n285), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n274), .B1(new_n369), .B2(new_n373), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n299), .A2(G232), .A3(new_n284), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n298), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n333), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n364), .A2(new_n366), .A3(new_n383), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n384), .B(KEYINPUT17), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n375), .A2(new_n312), .A3(new_n377), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n294), .B1(new_n379), .B2(new_n381), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(new_n364), .B2(new_n366), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT18), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI211_X1 g0191(.A(KEYINPUT18), .B(new_n388), .C1(new_n364), .C2(new_n366), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT79), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT79), .ZN(new_n394));
  INV_X1    g0194(.A(new_n366), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n360), .A2(new_n362), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n314), .B1(new_n396), .B2(new_n337), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n395), .B1(new_n397), .B2(new_n363), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT18), .B1(new_n398), .B2(new_n388), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n389), .A2(new_n390), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n394), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n385), .B1(new_n393), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(G226), .A2(G1698), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(new_n230), .B2(G1698), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n266), .ZN(new_n405));
  INV_X1    g0205(.A(G33), .ZN(new_n406));
  INV_X1    g0206(.A(G97), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n408), .A2(new_n275), .B1(G238), .B2(new_n281), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT73), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT72), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n298), .B(new_n411), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT13), .A4(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT13), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT73), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n410), .A2(KEYINPUT13), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n298), .B(KEYINPUT72), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n404), .A2(new_n266), .B1(G33), .B2(G97), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n418), .A2(new_n274), .B1(new_n303), .B2(new_n300), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n415), .B(new_n416), .C1(new_n417), .C2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n413), .A2(new_n420), .A3(G169), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT14), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n409), .A2(KEYINPUT74), .A3(KEYINPUT13), .A4(new_n412), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT74), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n417), .A2(new_n419), .B1(new_n424), .B2(new_n414), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(G179), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT14), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n413), .A2(new_n420), .A3(new_n428), .A4(G169), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n422), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT11), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n338), .A2(G20), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n250), .B2(new_n208), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT75), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(new_n247), .B2(G50), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n247), .A2(new_n434), .A3(G50), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n433), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n431), .B1(new_n438), .B2(new_n314), .ZN(new_n439));
  INV_X1    g0239(.A(new_n437), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(new_n435), .ZN(new_n441));
  OAI211_X1 g0241(.A(KEYINPUT11), .B(new_n254), .C1(new_n441), .C2(new_n433), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT76), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n439), .A2(KEYINPUT76), .A3(new_n442), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n338), .B1(new_n256), .B2(G20), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT12), .B1(new_n328), .B2(G68), .ZN(new_n448));
  INV_X1    g0248(.A(G13), .ZN(new_n449));
  OR4_X1    g0249(.A1(KEYINPUT12), .A2(new_n432), .A3(G1), .A4(new_n449), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n325), .A2(new_n447), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n445), .A2(new_n446), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n430), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n376), .B1(new_n423), .B2(new_n425), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(new_n452), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n413), .A2(new_n420), .A3(G200), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n336), .A2(new_n402), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n306), .A2(KEYINPUT6), .A3(G97), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n407), .A2(new_n306), .ZN(new_n461));
  NOR2_X1   g0261(.A1(G97), .A2(G107), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n460), .B1(new_n463), .B2(KEYINPUT6), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n464), .A2(G20), .B1(G77), .B2(new_n247), .ZN(new_n465));
  OAI21_X1  g0265(.A(G107), .B1(new_n358), .B2(new_n359), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n314), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n258), .A2(new_n407), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n406), .A2(G1), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n254), .A2(new_n258), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n468), .B1(new_n471), .B2(new_n407), .ZN(new_n472));
  OR2_X1    g0272(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT4), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(G1698), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n475), .B(G244), .C1(new_n343), .C2(new_n342), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G283), .ZN(new_n477));
  INV_X1    g0277(.A(G244), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n478), .B1(new_n264), .B2(new_n265), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n476), .B(new_n477), .C1(new_n479), .C2(KEYINPUT4), .ZN(new_n480));
  OAI21_X1  g0280(.A(G250), .B1(new_n342), .B2(new_n343), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n267), .B1(new_n481), .B2(KEYINPUT4), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT80), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G250), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n484), .B1(new_n264), .B2(new_n265), .ZN(new_n485));
  OAI21_X1  g0285(.A(G1698), .B1(new_n485), .B2(new_n474), .ZN(new_n486));
  OAI21_X1  g0286(.A(G244), .B1(new_n342), .B2(new_n343), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n487), .A2(new_n474), .B1(G33), .B2(G283), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT80), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n486), .A2(new_n488), .A3(new_n489), .A4(new_n476), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n483), .A2(new_n275), .A3(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n256), .B(G45), .C1(new_n277), .C2(KEYINPUT5), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT5), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(G41), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n299), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(G257), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT82), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n278), .A2(G1), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n277), .A2(KEYINPUT5), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n493), .A2(G41), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT82), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n501), .A2(new_n502), .A3(G257), .A4(new_n299), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT81), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n492), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n498), .A2(KEYINPUT81), .A3(new_n500), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n283), .A2(new_n499), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n497), .A2(new_n503), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n491), .A2(new_n312), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n497), .A2(new_n503), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n505), .A2(new_n506), .A3(new_n283), .A4(new_n499), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n486), .A2(new_n488), .A3(new_n476), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n274), .B1(new_n515), .B2(KEYINPUT80), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n514), .B1(new_n516), .B2(new_n490), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n473), .B(new_n511), .C1(new_n517), .C2(G169), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n266), .A2(new_n222), .A3(G68), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT19), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n222), .B1(new_n406), .B2(new_n407), .ZN(new_n521));
  INV_X1    g0321(.A(G87), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n462), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n520), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n250), .A2(KEYINPUT19), .A3(new_n407), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n519), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n314), .B1(new_n526), .B2(KEYINPUT85), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT85), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n519), .B(new_n528), .C1(new_n524), .C2(new_n525), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n328), .B1(new_n318), .B2(new_n317), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT86), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n471), .B2(new_n319), .ZN(new_n534));
  INV_X1    g0334(.A(new_n319), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n535), .A2(KEYINPUT86), .A3(new_n470), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n530), .A2(new_n532), .A3(new_n534), .A4(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n498), .A2(new_n282), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n484), .B1(new_n278), .B2(G1), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(new_n299), .A3(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(G238), .B(new_n267), .C1(new_n342), .C2(new_n343), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G116), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(G244), .B(G1698), .C1(new_n342), .C2(new_n343), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT83), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n266), .A2(KEYINPUT83), .A3(G244), .A4(G1698), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n543), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n275), .B1(new_n548), .B2(KEYINPUT84), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT84), .ZN(new_n550));
  AOI211_X1 g0350(.A(new_n550), .B(new_n543), .C1(new_n546), .C2(new_n547), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n312), .B(new_n540), .C1(new_n549), .C2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n540), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n541), .A2(new_n542), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT83), .B1(new_n479), .B2(G1698), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n544), .A2(new_n545), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n274), .B1(new_n557), .B2(new_n550), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n548), .A2(KEYINPUT84), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n553), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n537), .B(new_n552), .C1(new_n560), .C2(G169), .ZN(new_n561));
  OAI211_X1 g0361(.A(G190), .B(new_n540), .C1(new_n549), .C2(new_n551), .ZN(new_n562));
  NOR4_X1   g0362(.A1(new_n254), .A2(new_n258), .A3(new_n522), .A4(new_n469), .ZN(new_n563));
  AOI211_X1 g0363(.A(new_n531), .B(new_n563), .C1(new_n527), .C2(new_n529), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n562), .B(new_n564), .C1(new_n560), .C2(new_n333), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n491), .A2(G190), .A3(new_n510), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n467), .A2(new_n472), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n566), .B(new_n567), .C1(new_n517), .C2(new_n333), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n518), .A2(new_n561), .A3(new_n565), .A4(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n266), .A2(G257), .A3(G1698), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n266), .A2(G250), .A3(new_n267), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G33), .A2(G294), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n495), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n573), .A2(new_n275), .B1(G264), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n513), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n294), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n312), .A3(new_n513), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT24), .ZN(new_n579));
  OAI21_X1  g0379(.A(KEYINPUT23), .B1(new_n222), .B2(G107), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT23), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n581), .A2(new_n306), .A3(G20), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n222), .A2(G33), .A3(G116), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT89), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT89), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n580), .A2(new_n582), .A3(new_n583), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n222), .B(G87), .C1(new_n342), .C2(new_n343), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT22), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT22), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n266), .A2(new_n591), .A3(new_n222), .A4(G87), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n579), .B1(new_n588), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n588), .A2(new_n593), .A3(new_n579), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n314), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT25), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n257), .B2(G107), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n258), .A2(KEYINPUT25), .A3(new_n306), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n470), .A2(G107), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n577), .B(new_n578), .C1(new_n597), .C2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n501), .A2(G270), .A3(new_n299), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n513), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(G264), .B(G1698), .C1(new_n342), .C2(new_n343), .ZN(new_n607));
  OAI211_X1 g0407(.A(G257), .B(new_n267), .C1(new_n342), .C2(new_n343), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n264), .A2(G303), .A3(new_n265), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT87), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n275), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n611), .B1(new_n610), .B2(new_n275), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n606), .B(G179), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n614), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n605), .B1(new_n616), .B2(new_n612), .ZN(new_n617));
  NAND2_X1  g0417(.A1(KEYINPUT21), .A2(G169), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n615), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(G116), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n469), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n328), .A2(new_n314), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT88), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(G20), .B1(G33), .B2(G283), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n406), .A2(G97), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n625), .A2(new_n626), .B1(G20), .B2(new_n620), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n254), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT20), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n627), .A2(new_n254), .A3(KEYINPUT20), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n324), .A2(new_n620), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n328), .A2(KEYINPUT88), .A3(new_n314), .A4(new_n621), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n624), .A2(new_n632), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n619), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n606), .B1(new_n613), .B2(new_n614), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n637), .A2(new_n635), .A3(G169), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT21), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n603), .A2(new_n636), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n635), .B1(G200), .B2(new_n637), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n642), .B1(new_n376), .B2(new_n637), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n576), .A2(G200), .ZN(new_n644));
  INV_X1    g0444(.A(new_n596), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n254), .B1(new_n645), .B2(new_n594), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n575), .A2(G190), .A3(new_n513), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n644), .A2(new_n646), .A3(new_n601), .A4(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n569), .A2(new_n641), .A3(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n459), .A2(new_n650), .ZN(G372));
  INV_X1    g0451(.A(new_n385), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n311), .A2(G169), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n331), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n457), .A2(new_n313), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n652), .B1(new_n655), .B2(new_n453), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT90), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n391), .B2(new_n392), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n399), .A2(KEYINPUT90), .A3(new_n400), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n293), .B1(new_n656), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n296), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT91), .ZN(new_n663));
  INV_X1    g0463(.A(new_n561), .ZN(new_n664));
  AND4_X1   g0464(.A1(new_n518), .A2(new_n561), .A3(new_n565), .A4(new_n568), .ZN(new_n665));
  AND4_X1   g0465(.A1(new_n646), .A2(new_n644), .A3(new_n601), .A4(new_n647), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n619), .A2(new_n635), .B1(new_n638), .B2(new_n639), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n666), .B1(new_n667), .B2(new_n603), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n664), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT26), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n561), .A2(new_n565), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(new_n671), .B2(new_n518), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n491), .A2(new_n312), .A3(new_n510), .ZN(new_n673));
  AOI21_X1  g0473(.A(G169), .B1(new_n491), .B2(new_n510), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n673), .A2(new_n674), .A3(new_n567), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n675), .A2(KEYINPUT26), .A3(new_n561), .A4(new_n565), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n669), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n459), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n663), .A2(new_n679), .ZN(G369));
  NOR2_X1   g0480(.A1(new_n449), .A2(G1), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n222), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n681), .A2(new_n684), .A3(new_n222), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(G213), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT92), .ZN(new_n687));
  XOR2_X1   g0487(.A(KEYINPUT93), .B(G343), .Z(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n635), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n667), .B(new_n690), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n691), .A2(new_n643), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G330), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n603), .A2(new_n689), .ZN(new_n694));
  INV_X1    g0494(.A(new_n603), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n689), .B1(new_n597), .B2(new_n602), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n695), .B1(new_n648), .B2(new_n696), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n693), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n694), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n667), .A2(new_n689), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n603), .B2(new_n689), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n698), .A2(new_n702), .ZN(G399));
  NOR2_X1   g0503(.A1(new_n523), .A2(G116), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT94), .Z(new_n705));
  INV_X1    g0505(.A(new_n204), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n705), .A2(new_n256), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n225), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n708), .B1(new_n709), .B2(new_n707), .ZN(new_n710));
  XOR2_X1   g0510(.A(new_n710), .B(KEYINPUT28), .Z(new_n711));
  INV_X1    g0511(.A(new_n689), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n641), .A2(new_n648), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT98), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n713), .A2(new_n569), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(KEYINPUT98), .B1(new_n665), .B2(new_n668), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n561), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n676), .A2(KEYINPUT97), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT97), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n718), .B1(new_n677), .B2(new_n719), .ZN(new_n720));
  OAI211_X1 g0520(.A(KEYINPUT29), .B(new_n712), .C1(new_n717), .C2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n678), .A2(new_n712), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT29), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n637), .A2(new_n576), .A3(new_n312), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n725), .A2(new_n560), .A3(new_n517), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n540), .B(new_n575), .C1(new_n549), .C2(new_n551), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT96), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n491), .A2(new_n510), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n615), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n557), .A2(new_n550), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(new_n559), .A3(new_n275), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n733), .A2(KEYINPUT96), .A3(new_n540), .A4(new_n575), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n729), .A2(new_n731), .A3(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT30), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n726), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n729), .A2(new_n731), .A3(new_n734), .A4(KEYINPUT30), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n712), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g0539(.A(KEYINPUT95), .B(KEYINPUT31), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n641), .A2(new_n649), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(new_n665), .A3(new_n712), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n742), .B(new_n744), .C1(KEYINPUT31), .C2(new_n739), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n721), .A2(new_n724), .B1(G330), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n711), .B1(new_n746), .B2(G1), .ZN(G364));
  INV_X1    g0547(.A(new_n707), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n449), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n256), .B1(new_n749), .B2(G45), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n748), .A2(KEYINPUT99), .A3(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT99), .ZN(new_n752));
  INV_X1    g0552(.A(new_n750), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n752), .B1(new_n707), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n693), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n692), .A2(G330), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G13), .A2(G33), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G20), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n692), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n221), .B1(G20), .B2(new_n294), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR4_X1   g0565(.A1(new_n222), .A2(new_n333), .A3(G179), .A4(G190), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n306), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n222), .A2(new_n312), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G190), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR4_X1   g0572(.A1(new_n222), .A2(new_n376), .A3(new_n333), .A4(G179), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n772), .A2(new_n338), .B1(new_n522), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n770), .A2(new_n376), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n768), .B(new_n775), .C1(G50), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n376), .A2(G200), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n222), .B1(new_n778), .B2(new_n312), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT101), .Z(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G97), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G190), .A2(G200), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n782), .A2(G20), .A3(new_n312), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n354), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT32), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n769), .A2(new_n782), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n266), .B1(new_n786), .B2(new_n208), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n769), .A2(new_n778), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n787), .B1(G58), .B2(new_n789), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n777), .A2(new_n781), .A3(new_n785), .A4(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G322), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G311), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n344), .B1(new_n786), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n783), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n793), .B(new_n795), .C1(G329), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n766), .A2(G283), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT33), .B(G317), .ZN(new_n799));
  INV_X1    g0599(.A(new_n779), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n771), .A2(new_n799), .B1(new_n800), .B2(G294), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n776), .A2(G326), .B1(G303), .B2(new_n773), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n797), .A2(new_n798), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n765), .B1(new_n791), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n706), .A2(new_n344), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n805), .A2(G355), .B1(new_n620), .B2(new_n706), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n245), .A2(new_n278), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n706), .A2(new_n266), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n226), .B2(G45), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n806), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT100), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n764), .A2(new_n761), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  NOR3_X1   g0616(.A1(new_n804), .A2(new_n816), .A3(new_n755), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n758), .B1(new_n763), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(G396));
  INV_X1    g0619(.A(new_n786), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G143), .A2(new_n789), .B1(new_n820), .B2(G159), .ZN(new_n821));
  INV_X1    g0621(.A(G150), .ZN(new_n822));
  INV_X1    g0622(.A(G137), .ZN(new_n823));
  INV_X1    g0623(.A(new_n776), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n821), .B1(new_n772), .B2(new_n822), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  XOR2_X1   g0625(.A(KEYINPUT102), .B(KEYINPUT34), .Z(new_n826));
  XNOR2_X1  g0626(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n767), .A2(new_n338), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n344), .B(new_n828), .C1(G132), .C2(new_n796), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n800), .A2(G58), .B1(new_n773), .B2(G50), .ZN(new_n830));
  AND3_X1   g0630(.A1(new_n827), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G294), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n788), .A2(new_n832), .B1(new_n786), .B2(new_n620), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n266), .B(new_n833), .C1(G311), .C2(new_n796), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n776), .A2(G303), .B1(G87), .B2(new_n766), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n771), .A2(G283), .B1(G107), .B2(new_n773), .ZN(new_n836));
  AND4_X1   g0636(.A1(new_n781), .A2(new_n834), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n764), .B1(new_n831), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n764), .A2(new_n759), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n755), .B1(new_n839), .B2(new_n208), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n330), .A2(new_n689), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n689), .B1(new_n323), .B2(new_n329), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n334), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n841), .B1(new_n330), .B2(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n838), .B(new_n840), .C1(new_n844), .C2(new_n760), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n843), .A2(new_n330), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n654), .A2(new_n313), .A3(new_n712), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n722), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n335), .A2(new_n712), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n672), .A2(new_n676), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n561), .B1(new_n713), .B2(new_n569), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n745), .A2(G330), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n755), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n855), .A2(new_n856), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n845), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT103), .ZN(G384));
  OR2_X1    g0661(.A1(new_n464), .A2(KEYINPUT35), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n464), .A2(KEYINPUT35), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n862), .A2(G116), .A3(new_n223), .A4(new_n863), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n864), .B(KEYINPUT36), .Z(new_n865));
  NAND4_X1  g0665(.A1(new_n709), .A2(G77), .A3(new_n349), .A4(new_n352), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n255), .A2(G68), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n256), .B(G13), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT91), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n662), .B(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n721), .A2(new_n459), .A3(new_n724), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(KEYINPUT105), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT105), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n721), .A2(new_n459), .A3(new_n874), .A4(new_n724), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT39), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n687), .B1(new_n364), .B2(new_n366), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n402), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n364), .A2(new_n366), .ZN(new_n880));
  INV_X1    g0680(.A(new_n388), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n687), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n882), .A2(new_n884), .A3(new_n885), .A4(new_n384), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT104), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n384), .B1(new_n398), .B2(new_n687), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT37), .B1(new_n888), .B2(new_n389), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g0690(.A(KEYINPUT104), .B(KEYINPUT37), .C1(new_n888), .C2(new_n389), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n879), .A2(KEYINPUT38), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n658), .A2(new_n659), .A3(new_n385), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n878), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n884), .A2(KEYINPUT90), .A3(new_n384), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n364), .A2(new_n366), .A3(new_n383), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n897), .A2(new_n878), .ZN(new_n898));
  AOI22_X1  g0698(.A1(KEYINPUT37), .A2(new_n896), .B1(new_n898), .B2(new_n882), .ZN(new_n899));
  NOR4_X1   g0699(.A1(new_n888), .A2(KEYINPUT90), .A3(new_n885), .A4(new_n389), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n895), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n877), .B1(new_n893), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n430), .A2(new_n452), .A3(new_n712), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n890), .A2(new_n891), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT79), .B1(new_n391), .B2(new_n392), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n399), .A2(new_n394), .A3(new_n400), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n884), .B1(new_n910), .B2(new_n385), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n906), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n879), .A2(KEYINPUT38), .A3(new_n892), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(KEYINPUT39), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n903), .A2(new_n905), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n452), .A2(new_n689), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n453), .A2(new_n457), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n916), .B1(new_n453), .B2(new_n457), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n854), .B2(new_n847), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n912), .A2(new_n913), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n920), .A2(new_n921), .B1(new_n660), .B2(new_n687), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n915), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n876), .B(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(G330), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n402), .A2(new_n878), .B1(new_n890), .B2(new_n891), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n902), .B1(KEYINPUT38), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n916), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n458), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n453), .A2(new_n457), .A3(new_n916), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n848), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n744), .B1(new_n739), .B2(new_n741), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n739), .A2(KEYINPUT31), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT40), .B1(new_n927), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n844), .B1(new_n917), .B2(new_n918), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n735), .A2(new_n736), .ZN(new_n937));
  INV_X1    g0737(.A(new_n726), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n937), .A2(new_n738), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n689), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n940), .A2(new_n740), .B1(new_n650), .B2(new_n712), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n739), .A2(KEYINPUT31), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n936), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT40), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n921), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n935), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n941), .A2(new_n942), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n459), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n925), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n948), .B2(new_n946), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n924), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n256), .B2(new_n749), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n924), .A2(new_n950), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n869), .B1(new_n952), .B2(new_n953), .ZN(G367));
  OAI211_X1 g0754(.A(new_n518), .B(new_n568), .C1(new_n567), .C2(new_n712), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n675), .A2(new_n689), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n699), .A2(new_n700), .A3(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT42), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n518), .B1(new_n955), .B2(new_n603), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n958), .A2(KEYINPUT42), .B1(new_n712), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n712), .A2(new_n564), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n664), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n671), .B2(new_n962), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n959), .A2(new_n961), .B1(KEYINPUT43), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n965), .B(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n698), .A2(new_n957), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n967), .B(new_n968), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n707), .B(KEYINPUT41), .Z(new_n970));
  XNOR2_X1  g0770(.A(new_n699), .B(new_n700), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(new_n693), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT108), .Z(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n693), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT107), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n976), .A2(new_n746), .ZN(new_n977));
  INV_X1    g0777(.A(new_n957), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n702), .A2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT44), .Z(new_n980));
  NOR2_X1   g0780(.A1(new_n702), .A2(new_n978), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT45), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n980), .A2(KEYINPUT106), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n698), .ZN(new_n984));
  AND3_X1   g0784(.A1(new_n980), .A2(new_n984), .A3(new_n982), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n984), .B1(new_n980), .B2(new_n982), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n977), .B(new_n983), .C1(new_n987), .C2(KEYINPUT106), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n970), .B1(new_n988), .B2(new_n746), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n969), .B1(new_n989), .B2(new_n753), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n815), .B1(new_n236), .B2(new_n808), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n535), .A2(new_n706), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n755), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(G303), .ZN(new_n994));
  INV_X1    g0794(.A(G283), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n788), .A2(new_n994), .B1(new_n786), .B2(new_n995), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n266), .B(new_n996), .C1(G317), .C2(new_n796), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n773), .A2(G116), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT46), .ZN(new_n999));
  AOI22_X1  g0799(.A1(G311), .A2(new_n776), .B1(new_n800), .B2(G107), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n767), .A2(new_n407), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(G294), .B2(new_n771), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n771), .A2(G159), .B1(new_n820), .B2(G50), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT109), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n780), .A2(G68), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n266), .B1(new_n783), .B2(new_n823), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G150), .B2(new_n789), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n773), .A2(G58), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n767), .A2(new_n208), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G143), .B2(new_n776), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1006), .A2(new_n1008), .A3(new_n1009), .A4(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1003), .B1(new_n1005), .B2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT47), .Z(new_n1014));
  OAI221_X1 g0814(.A(new_n993), .B1(new_n1014), .B2(new_n765), .C1(new_n762), .C2(new_n964), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n990), .A2(new_n1015), .ZN(G387));
  NOR2_X1   g0816(.A1(new_n977), .A2(new_n748), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n746), .B2(new_n976), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n761), .B1(new_n697), .B2(new_n694), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n755), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n705), .A2(new_n805), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(G107), .B2(new_n204), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n808), .ZN(new_n1023));
  AOI211_X1 g0823(.A(G45), .B(new_n705), .C1(G68), .C2(G77), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n321), .A2(new_n255), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT50), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1023), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT110), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n233), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n1028), .A2(new_n1029), .B1(new_n1031), .B2(G45), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1022), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1020), .B1(new_n1033), .B2(new_n815), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n786), .A2(new_n338), .B1(new_n783), .B2(new_n822), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n344), .B(new_n1035), .C1(G50), .C2(new_n789), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n780), .A2(new_n535), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1001), .B1(G77), .B2(new_n773), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G159), .A2(new_n776), .B1(new_n771), .B2(new_n321), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n266), .B1(new_n796), .B2(G326), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G303), .A2(new_n820), .B1(new_n789), .B2(G317), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n772), .B2(new_n794), .C1(new_n792), .C2(new_n824), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT48), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n800), .A2(G283), .B1(new_n773), .B2(G294), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT49), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT111), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1041), .B1(new_n620), .B2(new_n767), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1049), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1052), .A2(KEYINPUT111), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1040), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1034), .B1(new_n1054), .B2(new_n764), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n976), .A2(new_n753), .B1(new_n1019), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1018), .A2(new_n1056), .ZN(G393));
  NAND2_X1  g0857(.A1(new_n987), .A2(new_n753), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n814), .B1(new_n407), .B2(new_n204), .C1(new_n241), .C2(new_n1023), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n1020), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n774), .A2(new_n338), .B1(new_n767), .B2(new_n522), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n771), .B2(G50), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n780), .A2(G77), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n820), .A2(new_n321), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n344), .B1(new_n796), .B2(G143), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n776), .A2(G150), .B1(new_n789), .B2(G159), .ZN(new_n1067));
  XOR2_X1   g0867(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n1068));
  XNOR2_X1  g0868(.A(new_n1067), .B(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n776), .A2(G317), .B1(new_n789), .B2(G311), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT52), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n768), .B1(G116), .B2(new_n800), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n344), .B1(new_n786), .B2(new_n832), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(G322), .B2(new_n796), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n771), .A2(G303), .B1(G283), .B2(new_n773), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n1066), .A2(new_n1069), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1060), .B1(new_n1077), .B2(new_n764), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n957), .B2(new_n762), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1058), .A2(new_n1079), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n988), .A2(new_n707), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n977), .A2(new_n987), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(G390));
  XNOR2_X1  g0884(.A(new_n904), .B(KEYINPUT113), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n927), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n718), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n852), .B2(KEYINPUT97), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n714), .B1(new_n713), .B2(new_n569), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n665), .A2(KEYINPUT98), .A3(new_n668), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n664), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n689), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n841), .B1(new_n1092), .B2(new_n846), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1086), .B1(new_n1093), .B2(new_n919), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n903), .A2(new_n914), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT114), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n920), .B2(new_n905), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n929), .A2(new_n930), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n850), .B1(new_n669), .B2(new_n677), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1098), .B1(new_n1099), .B2(new_n841), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1100), .A2(KEYINPUT114), .A3(new_n904), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1095), .A2(new_n1097), .A3(new_n1101), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n745), .A2(G330), .A3(new_n844), .A4(new_n1098), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1094), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1100), .A2(new_n904), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1096), .A2(new_n1105), .B1(new_n903), .B2(new_n914), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n712), .B(new_n846), .C1(new_n717), .C2(new_n720), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n847), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n1098), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1106), .A2(new_n1101), .B1(new_n1109), .B2(new_n1086), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n925), .B1(new_n941), .B2(new_n942), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n931), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1104), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n745), .A2(G330), .A3(new_n844), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1114), .A2(new_n919), .B1(new_n1111), .B2(new_n931), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1099), .A2(new_n841), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1103), .A2(new_n847), .A3(new_n1107), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1098), .B1(new_n1111), .B2(new_n844), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1115), .A2(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n459), .A2(new_n1111), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1119), .A2(new_n873), .A3(new_n875), .A4(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n748), .B1(new_n1113), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n1113), .B2(new_n1121), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1113), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1095), .A2(new_n759), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n788), .A2(new_n620), .B1(new_n783), .B2(new_n832), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n266), .B(new_n1126), .C1(G97), .C2(new_n820), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n828), .B1(G87), .B2(new_n773), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n771), .A2(G107), .B1(new_n776), .B2(G283), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1127), .A2(new_n1063), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n780), .A2(G159), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n776), .A2(G128), .B1(G50), .B2(new_n766), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1131), .B(new_n1132), .C1(new_n823), .C2(new_n772), .ZN(new_n1133));
  OR3_X1    g0933(.A1(new_n774), .A2(KEYINPUT53), .A3(new_n822), .ZN(new_n1134));
  OAI21_X1  g0934(.A(KEYINPUT53), .B1(new_n774), .B2(new_n822), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n344), .B1(new_n796), .B2(G125), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT54), .B(G143), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(G132), .A2(new_n789), .B1(new_n820), .B2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .A4(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1130), .B1(new_n1133), .B2(new_n1140), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1141), .A2(new_n764), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n755), .B(new_n1142), .C1(new_n249), .C2(new_n839), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1124), .A2(new_n753), .B1(new_n1125), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1123), .A2(new_n1144), .ZN(G378));
  INV_X1    g0945(.A(KEYINPUT118), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n872), .A2(KEYINPUT105), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1147), .A2(new_n663), .A3(new_n875), .A4(new_n1120), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n1113), .B2(new_n1121), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n883), .A2(new_n262), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n297), .B(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1152), .B(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n925), .B1(new_n935), .B2(new_n945), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1156), .A2(new_n923), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n923), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1155), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n946), .A2(G330), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n915), .A2(new_n922), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1156), .A2(new_n923), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n1154), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1159), .A2(new_n1164), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1150), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1146), .B1(new_n1166), .B2(KEYINPUT57), .ZN(new_n1167));
  AOI21_X1  g0967(.A(KEYINPUT57), .B1(new_n1150), .B2(new_n1165), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(KEYINPUT118), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1150), .A2(new_n1165), .A3(KEYINPUT57), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1167), .A2(new_n707), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1165), .A2(new_n753), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n266), .A2(G41), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n255), .B1(G33), .B2(G41), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1173), .B1(new_n995), .B2(new_n783), .C1(new_n306), .C2(new_n788), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n535), .B2(new_n820), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n773), .A2(G77), .B1(new_n766), .B2(G58), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n771), .A2(G97), .B1(new_n776), .B2(G116), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1177), .A2(new_n1006), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT58), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1175), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n1181), .B2(new_n1180), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G128), .A2(new_n789), .B1(new_n773), .B2(new_n1138), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT115), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n780), .A2(G150), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n771), .A2(G132), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n776), .A2(G125), .B1(new_n820), .B2(G137), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT116), .Z(new_n1190));
  OR2_X1    g0990(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1191));
  AOI211_X1 g0991(.A(G33), .B(G41), .C1(new_n796), .C2(G124), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n354), .B2(new_n767), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1190), .B2(KEYINPUT59), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1183), .B1(new_n1191), .B2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1195), .A2(new_n765), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT117), .Z(new_n1197));
  AOI21_X1  g0997(.A(new_n755), .B1(new_n839), .B2(new_n255), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(new_n1155), .C2(new_n760), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1172), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1171), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(KEYINPUT119), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT119), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1171), .A2(new_n1204), .A3(new_n1201), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(G375));
  NAND2_X1  g1007(.A1(new_n919), .A2(new_n759), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n788), .A2(new_n995), .B1(new_n783), .B2(new_n994), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n266), .B(new_n1209), .C1(G107), .C2(new_n820), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1010), .B1(G294), .B2(new_n776), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n771), .A2(G116), .B1(G97), .B2(new_n773), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1210), .A2(new_n1037), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n780), .A2(G50), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n788), .A2(new_n823), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n266), .B1(new_n786), .B2(new_n822), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(G128), .C2(new_n796), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n771), .A2(new_n1138), .B1(G58), .B2(new_n766), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n776), .A2(G132), .B1(G159), .B2(new_n773), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1214), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n765), .B1(new_n1213), .B2(new_n1220), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n755), .B(new_n1221), .C1(new_n338), .C2(new_n839), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1119), .A2(new_n753), .B1(new_n1208), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n970), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1121), .A2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1149), .A2(new_n1119), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1223), .B1(new_n1225), .B2(new_n1226), .ZN(G381));
  INV_X1    g1027(.A(G378), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1083), .A2(new_n990), .A3(new_n1015), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NOR4_X1   g1030(.A1(G393), .A2(G396), .A3(G384), .A4(G381), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1206), .A2(new_n1228), .A3(new_n1230), .A4(new_n1231), .ZN(G407));
  AOI21_X1  g1032(.A(G378), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n688), .A2(G213), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT120), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1233), .A2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1236), .A2(G407), .A3(G213), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT121), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT121), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1236), .A2(G407), .A3(new_n1239), .A4(G213), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(G409));
  NAND2_X1  g1041(.A1(G387), .A2(G390), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1229), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(G393), .B(new_n818), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1244), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1246), .A2(new_n1229), .A3(new_n1242), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1234), .ZN(new_n1249));
  INV_X1    g1049(.A(G384), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1119), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1251), .A2(KEYINPUT60), .A3(new_n1148), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT122), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1251), .A2(KEYINPUT122), .A3(KEYINPUT60), .A4(new_n1148), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n707), .B1(new_n1251), .B2(new_n1148), .ZN(new_n1257));
  AOI21_X1  g1057(.A(KEYINPUT60), .B1(new_n1251), .B2(new_n1148), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1250), .B1(new_n1260), .B2(new_n1223), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1223), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n1262), .B(G384), .C1(new_n1256), .C2(new_n1259), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n707), .B(new_n1170), .C1(new_n1168), .C2(KEYINPUT118), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1146), .B(KEYINPUT57), .C1(new_n1150), .C2(new_n1165), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G378), .B(new_n1201), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1166), .A2(new_n1224), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1228), .B1(new_n1268), .B2(new_n1200), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n1249), .B(new_n1264), .C1(new_n1267), .C2(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1270), .A2(KEYINPUT62), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1235), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT126), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1272), .A2(KEYINPUT126), .A3(new_n1273), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1264), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1279), .A2(KEYINPUT62), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1271), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n1258), .B(new_n1257), .C1(new_n1254), .C2(new_n1255), .ZN(new_n1282));
  OAI21_X1  g1082(.A(G384), .B1(new_n1282), .B2(new_n1262), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1260), .A2(new_n1250), .A3(new_n1223), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1235), .A2(G2897), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1249), .A2(G2897), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1287), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT125), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1286), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1289), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1276), .A2(new_n1277), .A3(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT61), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1248), .B1(new_n1281), .B2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1278), .A2(KEYINPUT63), .A3(new_n1279), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT123), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1298), .B1(new_n1270), .B2(KEYINPUT63), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT63), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1272), .A2(new_n1234), .ZN(new_n1301));
  OAI211_X1 g1101(.A(KEYINPUT123), .B(new_n1300), .C1(new_n1301), .C2(new_n1264), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1301), .A2(KEYINPUT124), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT124), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1272), .A2(new_n1305), .A3(new_n1234), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1304), .A2(new_n1292), .A3(new_n1306), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1245), .A2(new_n1294), .A3(new_n1247), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1297), .A2(new_n1303), .A3(new_n1307), .A4(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1296), .A2(new_n1309), .ZN(G405));
  NAND2_X1  g1110(.A1(new_n1202), .A2(G378), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1264), .B1(new_n1233), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1205), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1204), .B1(new_n1171), .B2(new_n1201), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1228), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1316), .A2(new_n1279), .A3(new_n1311), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT127), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1245), .A2(new_n1318), .A3(new_n1247), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1313), .A2(new_n1317), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1248), .A2(KEYINPUT127), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1321), .A2(new_n1313), .A3(new_n1317), .A4(new_n1319), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(G402));
endmodule


