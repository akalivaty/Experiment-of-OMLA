//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 1 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT67), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G237), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(KEYINPUT86), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G214), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n196), .B1(KEYINPUT86), .B2(new_n193), .ZN(new_n197));
  AND4_X1   g011(.A1(new_n187), .A2(new_n192), .A3(new_n195), .A4(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(G953), .B1(new_n189), .B2(new_n191), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n195), .B1(new_n199), .B2(new_n197), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT18), .A3(G131), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n192), .A2(new_n187), .A3(new_n197), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(new_n194), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n199), .A2(new_n195), .A3(new_n197), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT18), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G125), .B(G140), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n210), .B(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n202), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(G113), .B(G122), .ZN(new_n214));
  INV_X1    g028(.A(G104), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n214), .B(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(G131), .B1(new_n204), .B2(new_n205), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n204), .A2(G131), .A3(new_n205), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT87), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT87), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n204), .A2(new_n221), .A3(G131), .A4(new_n205), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n218), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n210), .A2(KEYINPUT16), .ZN(new_n224));
  INV_X1    g038(.A(G125), .ZN(new_n225));
  OR3_X1    g039(.A1(new_n225), .A2(KEYINPUT16), .A3(G140), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(G146), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT75), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT75), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n224), .A2(new_n229), .A3(new_n226), .A4(G146), .ZN(new_n230));
  XOR2_X1   g044(.A(new_n210), .B(KEYINPUT19), .Z(new_n231));
  OAI211_X1 g045(.A(new_n228), .B(new_n230), .C1(new_n231), .C2(G146), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n213), .B(new_n217), .C1(new_n223), .C2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(G475), .A2(G902), .ZN(new_n234));
  INV_X1    g048(.A(new_n213), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n220), .A2(KEYINPUT17), .A3(new_n222), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT88), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n220), .A2(KEYINPUT88), .A3(KEYINPUT17), .A4(new_n222), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT17), .ZN(new_n240));
  INV_X1    g054(.A(new_n218), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n221), .B1(new_n201), .B2(G131), .ZN(new_n242));
  INV_X1    g056(.A(new_n222), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n240), .B(new_n241), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n238), .A2(new_n239), .B1(new_n244), .B2(KEYINPUT89), .ZN(new_n245));
  INV_X1    g059(.A(new_n227), .ZN(new_n246));
  AOI21_X1  g060(.A(G146), .B1(new_n224), .B2(new_n226), .ZN(new_n247));
  OR2_X1    g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI211_X1 g062(.A(KEYINPUT17), .B(new_n218), .C1(new_n220), .C2(new_n222), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT89), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n235), .B1(new_n245), .B2(new_n251), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n233), .B(new_n234), .C1(new_n252), .C2(new_n217), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT90), .B1(new_n253), .B2(KEYINPUT20), .ZN(new_n254));
  INV_X1    g068(.A(new_n233), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n238), .A2(new_n239), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n244), .A2(KEYINPUT89), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n223), .A2(new_n250), .A3(new_n240), .ZN(new_n258));
  INV_X1    g072(.A(new_n248), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n256), .A2(new_n257), .A3(new_n258), .A4(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n213), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n255), .B1(new_n261), .B2(new_n216), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT90), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT20), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n262), .A2(new_n263), .A3(new_n264), .A4(new_n234), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n253), .A2(KEYINPUT20), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n254), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  OR2_X1    g081(.A1(new_n216), .A2(KEYINPUT91), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n261), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G902), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n261), .B2(new_n268), .ZN(new_n271));
  OAI21_X1  g085(.A(G475), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G478), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(KEYINPUT15), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G128), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT13), .B1(new_n276), .B2(G143), .ZN(new_n277));
  INV_X1    g091(.A(G134), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(G128), .B(G143), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G122), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G116), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT92), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n283), .B(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G107), .ZN(new_n286));
  INV_X1    g100(.A(G116), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G122), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n285), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n286), .B1(new_n285), .B2(new_n288), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n281), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n285), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n288), .B(KEYINPUT14), .ZN(new_n294));
  OAI21_X1  g108(.A(G107), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n280), .B(new_n278), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n289), .A3(new_n296), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  XOR2_X1   g112(.A(KEYINPUT72), .B(G217), .Z(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT9), .B(G234), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n299), .A2(G953), .A3(new_n300), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n298), .A2(new_n301), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n270), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT93), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT93), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n306), .B(new_n270), .C1(new_n302), .C2(new_n303), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n275), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G952), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(G953), .ZN(new_n310));
  INV_X1    g124(.A(G234), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(new_n188), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  AOI211_X1 g127(.A(new_n270), .B(new_n187), .C1(G234), .C2(G237), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT21), .B(G898), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n274), .B1(new_n304), .B2(KEYINPUT93), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n308), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n267), .A2(new_n272), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT94), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT94), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n267), .A2(new_n321), .A3(new_n272), .A4(new_n318), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n299), .B1(G234), .B2(new_n270), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT25), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n210), .A2(new_n211), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n276), .A2(KEYINPUT23), .A3(G119), .ZN(new_n328));
  INV_X1    g142(.A(G119), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G128), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n329), .A2(G128), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n328), .B(new_n330), .C1(new_n331), .C2(KEYINPUT23), .ZN(new_n332));
  XOR2_X1   g146(.A(KEYINPUT74), .B(G110), .Z(new_n333));
  XOR2_X1   g147(.A(KEYINPUT24), .B(G110), .Z(new_n334));
  XNOR2_X1  g148(.A(G119), .B(G128), .ZN(new_n335));
  OAI22_X1  g149(.A1(new_n332), .A2(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n228), .A2(new_n230), .A3(new_n327), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n332), .A2(G110), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(KEYINPUT73), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n334), .A2(new_n335), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n340), .B1(new_n246), .B2(new_n247), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n337), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT22), .B(G137), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n343), .B(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(KEYINPUT76), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n337), .B(new_n345), .C1(new_n339), .C2(new_n341), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n326), .B1(new_n349), .B2(G902), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n347), .A2(KEYINPUT25), .A3(new_n270), .A4(new_n348), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n325), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NOR3_X1   g166(.A1(new_n349), .A2(G902), .A3(new_n324), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(G472), .A2(G902), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n329), .A2(G116), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n287), .A2(G119), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT2), .B(G113), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n359), .A2(new_n361), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT30), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT11), .B1(new_n278), .B2(G137), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT11), .ZN(new_n368));
  INV_X1    g182(.A(G137), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n369), .A3(G134), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT66), .B1(new_n369), .B2(G134), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT66), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n278), .A3(G137), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n371), .A2(new_n208), .A3(new_n372), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n211), .A2(G143), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n193), .A2(G146), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n376), .B(new_n377), .C1(KEYINPUT1), .C2(new_n276), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n377), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n376), .A2(KEYINPUT1), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(G128), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n278), .A2(G137), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n369), .A2(G134), .ZN(new_n383));
  OAI21_X1  g197(.A(G131), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n375), .A2(new_n378), .A3(new_n381), .A4(new_n384), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n367), .A2(new_n370), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n372), .A2(new_n374), .ZN(new_n387));
  OAI21_X1  g201(.A(G131), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n388), .A2(new_n375), .ZN(new_n389));
  AND2_X1   g203(.A1(KEYINPUT0), .A2(G128), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(new_n376), .B2(new_n377), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT0), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n276), .A3(KEYINPUT64), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT64), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n394), .B1(KEYINPUT0), .B2(G128), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT65), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n376), .A2(new_n377), .A3(new_n390), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n391), .A2(new_n396), .A3(KEYINPUT65), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n366), .B(new_n385), .C1(new_n389), .C2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n388), .A2(new_n375), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n401), .A2(new_n400), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(new_n399), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n366), .B1(new_n407), .B2(new_n385), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n365), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n199), .A2(G210), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n410), .B(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT26), .B(G101), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n365), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n415), .B(new_n385), .C1(new_n389), .C2(new_n402), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n409), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT69), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n409), .A2(KEYINPUT69), .A3(new_n414), .A4(new_n416), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n419), .A2(KEYINPUT31), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT31), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n409), .A2(new_n422), .A3(new_n414), .A4(new_n416), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n401), .A2(new_n400), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT65), .B1(new_n391), .B2(new_n396), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n375), .A2(new_n384), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n381), .A2(new_n378), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n426), .A2(new_n405), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(KEYINPUT28), .B1(new_n430), .B2(new_n415), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n431), .A2(KEYINPUT70), .ZN(new_n432));
  INV_X1    g246(.A(new_n416), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n415), .B1(new_n407), .B2(new_n385), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT28), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n431), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n432), .B1(new_n437), .B2(KEYINPUT70), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n423), .B1(new_n438), .B2(new_n414), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n356), .B1(new_n421), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT32), .ZN(new_n441));
  INV_X1    g255(.A(new_n356), .ZN(new_n442));
  INV_X1    g256(.A(new_n423), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT28), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n385), .B1(new_n389), .B2(new_n402), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n365), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n444), .B1(new_n446), .B2(new_n416), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT70), .B1(new_n447), .B2(new_n431), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT70), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n436), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n414), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n443), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n419), .A2(KEYINPUT31), .A3(new_n420), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n442), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT32), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n441), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G472), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n446), .A2(new_n416), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n431), .B1(new_n460), .B2(KEYINPUT28), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n414), .B(new_n450), .C1(new_n461), .C2(new_n449), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT71), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n448), .A2(KEYINPUT71), .A3(new_n414), .A4(new_n450), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n409), .A2(new_n416), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT29), .B1(new_n466), .B2(new_n452), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n464), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n448), .A2(KEYINPUT29), .A3(new_n414), .A4(new_n450), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n469), .A2(new_n270), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n459), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n355), .B1(new_n458), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT80), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT79), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT3), .B1(new_n215), .B2(G107), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT3), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(new_n286), .A3(G104), .ZN(new_n478));
  INV_X1    g292(.A(G101), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n215), .A2(G107), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n476), .A2(new_n478), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n215), .A2(G107), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n286), .A2(G104), .ZN(new_n483));
  OAI21_X1  g297(.A(G101), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n428), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n381), .A2(new_n378), .A3(new_n481), .A4(new_n484), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(KEYINPUT12), .A3(new_n405), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(KEYINPUT12), .B1(new_n488), .B2(new_n405), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n475), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n488), .A2(new_n405), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT12), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(KEYINPUT79), .A3(new_n489), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT77), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT4), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n476), .A2(new_n478), .A3(KEYINPUT77), .A4(new_n480), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n500), .A2(new_n501), .A3(G101), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT78), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n479), .B1(new_n498), .B2(new_n499), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT78), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n505), .A2(new_n506), .A3(new_n501), .A4(new_n502), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n481), .A2(KEYINPUT4), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n509), .B1(new_n505), .B2(new_n502), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n402), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g326(.A1(new_n487), .A2(KEYINPUT10), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n487), .A2(KEYINPUT10), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n512), .A2(new_n515), .A3(new_n389), .ZN(new_n516));
  XNOR2_X1  g330(.A(G110), .B(G140), .ZN(new_n517));
  INV_X1    g331(.A(G227), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(G953), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n517), .B(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n474), .B1(new_n497), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n508), .A2(new_n511), .B1(new_n514), .B2(new_n513), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n520), .B1(new_n524), .B2(new_n389), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n525), .A2(KEYINPUT80), .A3(new_n492), .A4(new_n496), .ZN(new_n526));
  INV_X1    g340(.A(new_n516), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n524), .A2(new_n389), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n520), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n523), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G469), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n270), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n531), .A2(new_n270), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n495), .A2(new_n489), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n521), .B1(new_n516), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(new_n522), .B2(new_n528), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n532), .B(new_n534), .C1(new_n531), .C2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(G221), .B1(new_n300), .B2(G902), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(G210), .B1(G237), .B2(G902), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(G224), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(G953), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT82), .ZN(new_n546));
  OAI21_X1  g360(.A(G125), .B1(new_n424), .B2(new_n425), .ZN(new_n547));
  AOI21_X1  g361(.A(G125), .B1(new_n381), .B2(new_n378), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n546), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT82), .B1(new_n402), .B2(G125), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n545), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n547), .A2(new_n546), .ZN(new_n553));
  INV_X1    g367(.A(new_n545), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n548), .B1(new_n402), .B2(G125), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n553), .B(new_n554), .C1(new_n555), .C2(new_n546), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n357), .A2(new_n358), .A3(KEYINPUT5), .ZN(new_n558));
  OAI21_X1  g372(.A(G113), .B1(new_n357), .B2(KEYINPUT5), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n363), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n560), .A2(new_n485), .ZN(new_n561));
  XNOR2_X1  g375(.A(G110), .B(G122), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n510), .A2(new_n415), .ZN(new_n564));
  AOI211_X1 g378(.A(new_n561), .B(new_n563), .C1(new_n508), .C2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT6), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n561), .B1(new_n508), .B2(new_n564), .ZN(new_n567));
  XOR2_X1   g381(.A(new_n562), .B(KEYINPUT81), .Z(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  OAI22_X1  g383(.A1(new_n565), .A2(new_n566), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n508), .A2(new_n564), .ZN(new_n571));
  INV_X1    g385(.A(new_n561), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(KEYINPUT6), .A3(new_n568), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n557), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n571), .A2(new_n572), .A3(new_n562), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n554), .A2(KEYINPUT7), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n550), .B2(new_n551), .ZN(new_n578));
  INV_X1    g392(.A(new_n577), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n553), .B(new_n579), .C1(new_n555), .C2(new_n546), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT84), .ZN(new_n581));
  INV_X1    g395(.A(new_n485), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n581), .B1(new_n582), .B2(KEYINPUT83), .ZN(new_n583));
  INV_X1    g397(.A(new_n560), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n562), .B(KEYINPUT8), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n560), .B1(KEYINPUT84), .B2(new_n485), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n585), .B(new_n586), .C1(new_n583), .C2(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n576), .A2(new_n578), .A3(new_n580), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n270), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n543), .B1(new_n575), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n552), .A2(new_n556), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n576), .A2(KEYINPUT6), .B1(new_n573), .B2(new_n568), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n567), .A2(new_n566), .A3(new_n569), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n589), .A2(new_n270), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(new_n596), .A3(new_n542), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n591), .A2(new_n597), .A3(KEYINPUT85), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n542), .B1(new_n595), .B2(new_n596), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT85), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(G214), .B1(G237), .B2(G902), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n598), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n541), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n323), .A2(new_n473), .A3(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT95), .B(G101), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G3));
  NAND2_X1  g421(.A1(new_n451), .A2(new_n452), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n454), .A2(new_n608), .A3(new_n423), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n459), .B1(new_n609), .B2(new_n270), .ZN(new_n610));
  NOR4_X1   g424(.A1(new_n541), .A2(new_n455), .A3(new_n355), .A4(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n302), .A2(new_n303), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n273), .A2(G902), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n616));
  INV_X1    g430(.A(new_n304), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n616), .B1(new_n617), .B2(G478), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n304), .A2(KEYINPUT96), .A3(new_n273), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n614), .A2(new_n615), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n316), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n575), .A2(new_n590), .A3(new_n543), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n621), .B(new_n602), .C1(new_n622), .C2(new_n599), .ZN(new_n623));
  AOI211_X1 g437(.A(new_n620), .B(new_n623), .C1(new_n267), .C2(new_n272), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n611), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT34), .B(G104), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  NOR2_X1   g441(.A1(new_n308), .A2(new_n317), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n262), .A2(new_n264), .A3(new_n234), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n266), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n629), .A2(new_n631), .A3(new_n272), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n623), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n611), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT35), .B(G107), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G9));
  NOR2_X1   g450(.A1(new_n610), .A2(new_n455), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n350), .A2(new_n351), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n324), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n346), .A2(KEYINPUT36), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(new_n342), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n324), .A2(G902), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n637), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT97), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n637), .A2(KEYINPUT97), .A3(new_n644), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n323), .A2(new_n604), .A3(new_n647), .A4(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT37), .B(G110), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT98), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n649), .B(new_n651), .ZN(G12));
  AOI21_X1  g466(.A(new_n471), .B1(new_n441), .B2(new_n457), .ZN(new_n653));
  INV_X1    g467(.A(new_n644), .ZN(new_n654));
  INV_X1    g468(.A(new_n602), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n591), .B2(new_n597), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n539), .A2(new_n540), .A3(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n653), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(G900), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n314), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n312), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n632), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G128), .ZN(G30));
  XNOR2_X1  g479(.A(new_n661), .B(KEYINPUT39), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n541), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT40), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n598), .A2(new_n601), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(KEYINPUT38), .Z(new_n671));
  NAND2_X1  g485(.A1(new_n267), .A2(new_n272), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n628), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n419), .A2(new_n420), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n414), .B1(new_n416), .B2(new_n446), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n270), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(G472), .ZN(new_n678));
  AOI211_X1 g492(.A(new_n655), .B(new_n644), .C1(new_n458), .C2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n669), .A2(new_n671), .A3(new_n674), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G143), .ZN(G45));
  INV_X1    g495(.A(new_n620), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n672), .A2(new_n682), .A3(new_n661), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT99), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n620), .B1(new_n267), .B2(new_n272), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT99), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n685), .A2(new_n686), .A3(new_n661), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n684), .A2(new_n658), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT100), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n684), .A2(new_n658), .A3(KEYINPUT100), .A4(new_n687), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G146), .ZN(G48));
  NAND2_X1  g507(.A1(new_n530), .A2(new_n270), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(G469), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n532), .ZN(new_n696));
  INV_X1    g510(.A(new_n540), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n473), .A2(new_n624), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT41), .B(G113), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G15));
  NAND3_X1  g515(.A1(new_n473), .A2(new_n633), .A3(new_n698), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G116), .ZN(G18));
  NAND4_X1  g517(.A1(new_n656), .A2(new_n695), .A3(new_n540), .A4(new_n532), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n653), .A2(new_n654), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n323), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G119), .ZN(G21));
  XNOR2_X1  g521(.A(new_n356), .B(KEYINPUT101), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n609), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT102), .ZN(new_n710));
  INV_X1    g524(.A(new_n353), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n639), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT102), .B1(new_n352), .B2(new_n353), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(G902), .B1(new_n453), .B2(new_n454), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n709), .B(new_n714), .C1(new_n715), .C2(new_n459), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT103), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n609), .A2(new_n270), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(G472), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n720), .A2(KEYINPUT103), .A3(new_n714), .A4(new_n709), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n656), .ZN(new_n723));
  AOI211_X1 g537(.A(new_n628), .B(new_n723), .C1(new_n267), .C2(new_n272), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n696), .A2(new_n316), .A3(new_n697), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n722), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  INV_X1    g541(.A(new_n704), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n720), .A2(new_n644), .A3(new_n709), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n684), .A2(new_n687), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G125), .ZN(G27));
  INV_X1    g545(.A(KEYINPUT42), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n684), .A2(new_n687), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT104), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n670), .B2(new_n602), .ZN(new_n735));
  AOI211_X1 g549(.A(KEYINPUT104), .B(new_n655), .C1(new_n598), .C2(new_n601), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n735), .A2(new_n736), .A3(new_n541), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n473), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n732), .B1(new_n733), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n714), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n653), .A2(new_n740), .A3(new_n732), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n684), .A2(new_n741), .A3(new_n737), .A4(new_n687), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g557(.A(KEYINPUT105), .B(G131), .Z(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(G33));
  NAND2_X1  g559(.A1(new_n670), .A2(new_n602), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT104), .ZN(new_n747));
  INV_X1    g561(.A(new_n541), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n670), .A2(new_n734), .A3(new_n602), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n440), .A2(KEYINPUT32), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n455), .A2(new_n456), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n472), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n354), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n663), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G134), .ZN(G36));
  NAND2_X1  g571(.A1(new_n673), .A2(new_n682), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT106), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n759), .A2(KEYINPUT43), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(KEYINPUT43), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n762), .B1(new_n758), .B2(new_n761), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n637), .A2(new_n654), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n763), .A2(KEYINPUT44), .A3(new_n764), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n522), .A2(new_n528), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(new_n536), .ZN(new_n770));
  OAI21_X1  g584(.A(G469), .B1(new_n770), .B2(KEYINPUT45), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT45), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n538), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n534), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT46), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n532), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n777), .B1(new_n774), .B2(new_n775), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n697), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n735), .A2(new_n736), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n779), .A2(new_n780), .A3(new_n666), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n767), .A2(new_n768), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G137), .ZN(G39));
  XNOR2_X1  g597(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n779), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n779), .A2(new_n784), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n780), .A2(new_n653), .A3(new_n355), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n733), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(G140), .Z(G42));
  NAND3_X1  g605(.A1(new_n714), .A2(new_n602), .A3(new_n540), .ZN(new_n792));
  AOI211_X1 g606(.A(new_n792), .B(new_n758), .C1(KEYINPUT49), .C2(new_n696), .ZN(new_n793));
  XOR2_X1   g607(.A(new_n793), .B(KEYINPUT108), .Z(new_n794));
  NAND2_X1  g608(.A1(new_n458), .A2(new_n678), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n696), .A2(KEYINPUT49), .ZN(new_n796));
  OR4_X1    g610(.A1(new_n671), .A2(new_n794), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n539), .A2(new_n540), .A3(new_n654), .A4(new_n661), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n799), .A2(KEYINPUT111), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n799), .A2(KEYINPUT111), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n795), .B(new_n724), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n730), .A2(new_n664), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n692), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n798), .B1(new_n804), .B2(KEYINPUT112), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n804), .A2(KEYINPUT112), .A3(new_n798), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AND4_X1   g622(.A1(new_n686), .A2(new_n672), .A3(new_n682), .A4(new_n661), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n686), .B1(new_n685), .B2(new_n661), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n729), .A3(new_n737), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT110), .ZN(new_n813));
  AND4_X1   g627(.A1(new_n272), .A2(new_n631), .A3(new_n628), .A4(new_n661), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n753), .A2(new_n644), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n813), .B1(new_n815), .B2(new_n750), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n653), .A2(new_n654), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n737), .A2(KEYINPUT110), .A3(new_n817), .A4(new_n814), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n812), .A2(new_n819), .A3(new_n756), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n603), .A2(new_n316), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n611), .A2(new_n673), .A3(new_n629), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n649), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n611), .A2(new_n822), .A3(new_n685), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n605), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n824), .B1(KEYINPUT109), .B2(new_n826), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n473), .B(new_n698), .C1(new_n624), .C2(new_n633), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n706), .A2(new_n828), .A3(new_n726), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n739), .B2(new_n742), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT109), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n605), .A2(new_n831), .A3(new_n825), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n821), .A2(new_n827), .A3(new_n830), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(KEYINPUT53), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n706), .A2(new_n828), .A3(new_n726), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT42), .B1(new_n811), .B2(new_n755), .ZN(new_n836));
  INV_X1    g650(.A(new_n742), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(new_n820), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n826), .A2(KEYINPUT109), .ZN(new_n840));
  INV_X1    g654(.A(new_n824), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n840), .A2(new_n841), .A3(new_n832), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n692), .A2(new_n803), .A3(KEYINPUT52), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT52), .B1(new_n692), .B2(new_n803), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n839), .B(new_n842), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n808), .A2(new_n834), .B1(new_n845), .B2(KEYINPUT53), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT54), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n829), .B(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n850), .B1(new_n739), .B2(new_n742), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n849), .A2(new_n821), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n808), .A2(new_n842), .A3(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT52), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n804), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n692), .A2(new_n803), .A3(KEYINPUT52), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n816), .A2(new_n818), .B1(new_n755), .B2(new_n663), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n743), .A2(new_n859), .A3(new_n812), .A4(new_n835), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n840), .A2(new_n841), .A3(new_n832), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI211_X1 g676(.A(new_n854), .B(KEYINPUT53), .C1(new_n858), .C2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT114), .B1(new_n845), .B2(new_n850), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n853), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n847), .B1(KEYINPUT54), .B2(new_n865), .ZN(new_n866));
  XOR2_X1   g680(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n867));
  AND3_X1   g681(.A1(new_n763), .A2(new_n313), .A3(new_n722), .ZN(new_n868));
  NOR4_X1   g682(.A1(new_n671), .A2(new_n602), .A3(new_n697), .A4(new_n696), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT50), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n780), .A2(new_n698), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n763), .A2(new_n313), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n729), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n355), .A2(new_n312), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n872), .A2(new_n458), .A3(new_n678), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n673), .A2(new_n620), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n871), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n868), .A2(new_n780), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n696), .A2(new_n540), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n787), .B2(KEYINPUT117), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(KEYINPUT117), .B2(new_n787), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n867), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n787), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n880), .B1(new_n886), .B2(new_n881), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n879), .A2(KEYINPUT51), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n653), .A2(new_n740), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n873), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT48), .ZN(new_n891));
  INV_X1    g705(.A(new_n685), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n310), .B1(new_n876), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n893), .B1(new_n868), .B2(new_n728), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n888), .A2(new_n891), .A3(new_n894), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n866), .A2(new_n885), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(G952), .A2(G953), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n797), .B1(new_n896), .B2(new_n897), .ZN(G75));
  NAND2_X1  g712(.A1(new_n309), .A2(G953), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT119), .Z(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n865), .A2(G210), .A3(G902), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT56), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n593), .A2(new_n594), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n557), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n595), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT55), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n901), .B1(new_n904), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT118), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n902), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n865), .A2(KEYINPUT118), .A3(G210), .A4(G902), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n908), .A2(KEYINPUT56), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n909), .A2(new_n914), .ZN(G51));
  XNOR2_X1  g729(.A(new_n533), .B(KEYINPUT57), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n843), .A2(new_n844), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n850), .B1(new_n918), .B2(new_n833), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n854), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n845), .A2(KEYINPUT114), .A3(new_n850), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n917), .B1(new_n922), .B2(new_n853), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n842), .A2(new_n849), .A3(new_n821), .A4(new_n851), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n807), .B2(new_n806), .ZN(new_n925));
  AOI211_X1 g739(.A(KEYINPUT54), .B(new_n925), .C1(new_n920), .C2(new_n921), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n916), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n530), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n865), .A2(G902), .ZN(new_n929));
  OR3_X1    g743(.A1(new_n929), .A2(new_n773), .A3(new_n771), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n901), .B1(new_n928), .B2(new_n930), .ZN(G54));
  INV_X1    g745(.A(new_n262), .ZN(new_n932));
  NAND2_X1  g746(.A1(KEYINPUT58), .A2(G475), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n932), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n900), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n929), .A2(new_n932), .A3(new_n933), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(G60));
  NOR2_X1   g751(.A1(new_n923), .A2(new_n926), .ZN(new_n938));
  XNOR2_X1  g752(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n939));
  NAND2_X1  g753(.A1(G478), .A2(G902), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n614), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n900), .B1(new_n938), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n614), .B1(new_n866), .B2(new_n941), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(G63));
  NAND2_X1  g759(.A1(G217), .A2(G902), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT60), .Z(new_n947));
  NAND2_X1  g761(.A1(new_n865), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n349), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n865), .A2(new_n641), .A3(new_n947), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n949), .A2(KEYINPUT61), .A3(new_n900), .A4(new_n950), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n949), .A2(new_n900), .A3(new_n950), .ZN(new_n952));
  XOR2_X1   g766(.A(KEYINPUT121), .B(KEYINPUT61), .Z(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(G66));
  OAI21_X1  g768(.A(G953), .B1(new_n315), .B2(new_n544), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n861), .A2(new_n829), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n955), .B1(new_n956), .B2(G953), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n905), .B1(G898), .B2(new_n187), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT122), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n957), .B(new_n959), .ZN(G69));
  AND2_X1   g774(.A1(new_n730), .A2(new_n664), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n692), .A2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n680), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n964), .A2(KEYINPUT62), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(KEYINPUT62), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n685), .B1(new_n673), .B2(new_n629), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n738), .A2(new_n667), .A3(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n790), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n965), .A2(new_n782), .A3(new_n966), .A4(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n187), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n404), .A2(new_n408), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n231), .B(KEYINPUT123), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n187), .A2(G900), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT125), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n889), .A2(new_n724), .A3(new_n779), .A4(new_n666), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n756), .B(new_n978), .C1(new_n789), .C2(new_n733), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n980), .A2(new_n743), .A3(new_n782), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n977), .B1(new_n981), .B2(new_n962), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n979), .B1(new_n739), .B2(new_n742), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n983), .A2(KEYINPUT125), .A3(new_n782), .A4(new_n963), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n976), .B1(new_n985), .B2(new_n187), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n975), .B1(new_n986), .B2(new_n974), .ZN(new_n987));
  OAI21_X1  g801(.A(G953), .B1(new_n518), .B2(new_n659), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT124), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n987), .B(new_n989), .ZN(G72));
  NAND3_X1  g804(.A1(new_n982), .A2(new_n956), .A3(new_n984), .ZN(new_n991));
  XOR2_X1   g805(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n992));
  NOR2_X1   g806(.A1(new_n459), .A2(new_n270), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n992), .B(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n466), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n995), .A2(new_n452), .A3(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n956), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n994), .B1(new_n970), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n999), .A2(new_n414), .A3(new_n466), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n997), .A2(new_n1000), .A3(new_n900), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n996), .A2(new_n414), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n846), .B(new_n994), .C1(new_n1002), .C2(new_n675), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT127), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OR2_X1    g819(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1001), .B1(new_n1005), .B2(new_n1006), .ZN(G57));
endmodule


