//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n860, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983, new_n984, new_n985;
  INV_X1    g000(.A(G169gat), .ZN(new_n202));
  INV_X1    g001(.A(G176gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT23), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(KEYINPUT25), .ZN(new_n210));
  INV_X1    g009(.A(G183gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(KEYINPUT24), .ZN(new_n212));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n212), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n210), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n214), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n215), .B(KEYINPUT65), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n209), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT25), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n217), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT27), .B(G183gat), .ZN(new_n223));
  INV_X1    g022(.A(G190gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n204), .A2(KEYINPUT26), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT67), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n204), .A2(KEYINPUT26), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n204), .A2(KEYINPUT67), .A3(KEYINPUT26), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .A4(new_n207), .ZN(new_n233));
  INV_X1    g032(.A(new_n213), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n234), .B1(new_n225), .B2(new_n226), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n227), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n222), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G113gat), .B(G120gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n239), .A2(KEYINPUT1), .ZN(new_n240));
  XOR2_X1   g039(.A(G127gat), .B(G134gat), .Z(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n238), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n242), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(new_n222), .B2(new_n237), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G227gat), .ZN(new_n247));
  INV_X1    g046(.A(G233gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT69), .B(KEYINPUT34), .Z(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n247), .A2(new_n248), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT64), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(KEYINPUT34), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n246), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G71gat), .B(G99gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT68), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(G15gat), .ZN(new_n259));
  INV_X1    g058(.A(G43gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n253), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n262), .B1(new_n243), .B2(new_n245), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n261), .B1(new_n263), .B2(KEYINPUT33), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT32), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n264), .A2(new_n266), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n256), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n269), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n249), .A2(new_n250), .B1(new_n246), .B2(new_n254), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(new_n272), .A3(new_n267), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT3), .ZN(new_n276));
  XNOR2_X1  g075(.A(G211gat), .B(G218gat), .ZN(new_n277));
  XOR2_X1   g076(.A(G197gat), .B(G204gat), .Z(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT70), .B(G218gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G211gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT22), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n278), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n277), .B1(new_n282), .B2(KEYINPUT86), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n283), .A2(KEYINPUT86), .A3(new_n282), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT29), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n283), .B1(KEYINPUT86), .B2(new_n282), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n276), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT2), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT83), .B(G155gat), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n289), .B1(new_n290), .B2(G162gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT84), .ZN(new_n292));
  INV_X1    g091(.A(G148gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G141gat), .ZN(new_n294));
  OR2_X1    g093(.A1(new_n294), .A2(KEYINPUT82), .ZN(new_n295));
  XNOR2_X1  g094(.A(G155gat), .B(G162gat), .ZN(new_n296));
  INV_X1    g095(.A(G141gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G148gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n298), .A2(new_n294), .A3(KEYINPUT82), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n295), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n292), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G155gat), .ZN(new_n303));
  INV_X1    g102(.A(G162gat), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT2), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT81), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n305), .A2(new_n306), .B1(new_n298), .B2(new_n294), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(new_n306), .B2(new_n305), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n296), .A2(KEYINPUT80), .ZN(new_n309));
  OR2_X1    g108(.A1(new_n296), .A2(KEYINPUT80), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n302), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n288), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n302), .A2(new_n276), .A3(new_n311), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT85), .ZN(new_n315));
  OR2_X1    g114(.A1(new_n291), .A2(KEYINPUT84), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n291), .A2(KEYINPUT84), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n300), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT85), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(new_n321), .A3(new_n276), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT29), .B1(new_n315), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n280), .A2(new_n281), .ZN(new_n324));
  INV_X1    g123(.A(new_n278), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT72), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n277), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT71), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT72), .B1(new_n282), .B2(KEYINPUT71), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n330), .B1(new_n331), .B2(new_n277), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n313), .B1(new_n323), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G228gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n335), .A2(new_n248), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n285), .B(new_n330), .C1(new_n331), .C2(new_n277), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n340), .A2(new_n276), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT87), .B1(new_n341), .B2(new_n320), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n276), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT87), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(new_n344), .A3(new_n312), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n342), .A2(new_n345), .A3(new_n336), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT73), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n347), .ZN(new_n348));
  OAI211_X1 g147(.A(KEYINPUT73), .B(new_n330), .C1(new_n331), .C2(new_n277), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n321), .B1(new_n320), .B2(new_n276), .ZN(new_n351));
  NOR4_X1   g150(.A1(new_n318), .A2(new_n319), .A3(KEYINPUT85), .A4(KEYINPUT3), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n285), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n350), .B1(new_n353), .B2(KEYINPUT88), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT88), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n323), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n346), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(G22gat), .B1(new_n339), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G22gat), .ZN(new_n359));
  INV_X1    g158(.A(new_n350), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(new_n323), .B2(new_n355), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n353), .A2(KEYINPUT88), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n359), .B(new_n338), .C1(new_n363), .C2(new_n346), .ZN(new_n364));
  XNOR2_X1  g163(.A(G78gat), .B(G106gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT31), .B(G50gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n358), .A2(new_n364), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n367), .B1(new_n358), .B2(new_n364), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n275), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G226gat), .A2(G233gat), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n371), .B(KEYINPUT74), .Z(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(new_n222), .B2(new_n237), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n218), .A2(new_n219), .ZN(new_n375));
  INV_X1    g174(.A(new_n209), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n377), .A2(KEYINPUT25), .B1(new_n210), .B2(new_n216), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT29), .B1(new_n378), .B2(new_n236), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n374), .B1(new_n379), .B2(new_n373), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT75), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n360), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n372), .B1(new_n378), .B2(new_n236), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n285), .B1(new_n222), .B2(new_n237), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n383), .B1(new_n372), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n333), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n381), .B1(new_n360), .B2(new_n380), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT76), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT75), .B1(new_n385), .B2(new_n350), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT76), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n390), .A2(new_n391), .A3(new_n382), .A4(new_n386), .ZN(new_n392));
  XOR2_X1   g191(.A(G8gat), .B(G36gat), .Z(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT77), .ZN(new_n394));
  XNOR2_X1  g193(.A(G64gat), .B(G92gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(KEYINPUT78), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n389), .A2(new_n392), .A3(new_n398), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n390), .A2(new_n386), .A3(new_n382), .A4(new_n396), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT30), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT79), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G1gat), .B(G29gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(KEYINPUT0), .ZN(new_n407));
  XNOR2_X1  g206(.A(G57gat), .B(G85gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(G225gat), .A2(G233gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n318), .A2(new_n244), .A3(new_n319), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n242), .B1(new_n302), .B2(new_n311), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT5), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n315), .A2(new_n322), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n242), .B1(new_n312), .B2(KEYINPUT3), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT4), .B1(new_n312), .B2(new_n244), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT4), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n413), .A2(new_n420), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n417), .A2(new_n418), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n416), .B1(new_n422), .B2(new_n411), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT5), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n418), .B1(new_n351), .B2(new_n352), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n421), .A2(new_n419), .ZN(new_n426));
  AND4_X1   g225(.A1(new_n424), .A2(new_n425), .A3(new_n411), .A4(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n410), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429));
  INV_X1    g228(.A(new_n416), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n425), .A2(new_n426), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n430), .B1(new_n431), .B2(new_n412), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n422), .A2(new_n424), .A3(new_n411), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n409), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n428), .A2(new_n429), .A3(new_n434), .ZN(new_n435));
  OAI211_X1 g234(.A(KEYINPUT6), .B(new_n410), .C1(new_n423), .C2(new_n427), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT30), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n400), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n399), .A2(new_n402), .A3(KEYINPUT79), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n405), .A2(new_n437), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT35), .B1(new_n370), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n358), .A2(new_n364), .ZN(new_n443));
  INV_X1    g242(.A(new_n367), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n358), .A2(new_n364), .A3(new_n367), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n274), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT35), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n399), .A2(new_n402), .A3(new_n448), .A4(new_n439), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT90), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n436), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n409), .B1(new_n432), .B2(new_n433), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(KEYINPUT90), .A3(KEYINPUT6), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n449), .B1(new_n454), .B2(new_n435), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n447), .A2(new_n455), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n270), .A2(new_n273), .A3(KEYINPUT36), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT36), .B1(new_n270), .B2(new_n273), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n368), .A2(new_n369), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n459), .B1(new_n441), .B2(new_n460), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n389), .A2(KEYINPUT37), .A3(new_n392), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT37), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n390), .A2(new_n463), .A3(new_n382), .A4(new_n386), .ZN(new_n464));
  INV_X1    g263(.A(new_n396), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT38), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n463), .B1(new_n385), .B2(new_n360), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n380), .A2(new_n333), .ZN(new_n469));
  AOI211_X1 g268(.A(KEYINPUT38), .B(new_n397), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n401), .B1(new_n464), .B2(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n467), .A2(new_n454), .A3(new_n435), .A4(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT39), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT89), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(new_n431), .B2(new_n412), .ZN(new_n475));
  AOI211_X1 g274(.A(KEYINPUT89), .B(new_n411), .C1(new_n425), .C2(new_n426), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT89), .B1(new_n422), .B2(new_n411), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n431), .A2(new_n474), .A3(new_n412), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n413), .A2(new_n414), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n473), .B1(new_n480), .B2(new_n411), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n477), .A2(new_n409), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT40), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n399), .A2(new_n402), .A3(new_n439), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n477), .A2(new_n482), .A3(KEYINPUT40), .A4(new_n409), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n485), .A2(new_n428), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n445), .A2(new_n446), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n472), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n442), .A2(new_n456), .B1(new_n461), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(G1gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT16), .ZN(new_n493));
  INV_X1    g292(.A(G15gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(G22gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n359), .A2(G15gat), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n493), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(G1gat), .B1(new_n495), .B2(new_n496), .ZN(new_n498));
  OAI21_X1  g297(.A(G8gat), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n495), .A2(new_n496), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n492), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n493), .A2(new_n495), .A3(new_n496), .ZN(new_n502));
  INV_X1    g301(.A(G8gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT93), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT93), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n499), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT15), .B1(new_n260), .B2(G50gat), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n510), .B1(new_n260), .B2(G50gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT15), .ZN(new_n512));
  INV_X1    g311(.A(G50gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT92), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT92), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(G50gat), .ZN(new_n516));
  AOI21_X1  g315(.A(G43gat), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT91), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(new_n260), .B2(G50gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n513), .A2(KEYINPUT91), .A3(G43gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n512), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT14), .B(G29gat), .ZN(new_n523));
  INV_X1    g322(.A(G36gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(G29gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n526), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n511), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n528), .A2(new_n511), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT17), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n528), .A2(new_n511), .ZN(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT92), .B(G50gat), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n519), .B(new_n520), .C1(new_n534), .C2(G43gat), .ZN(new_n535));
  AOI22_X1  g334(.A1(new_n535), .A2(new_n512), .B1(new_n525), .B2(new_n527), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n532), .B(new_n533), .C1(new_n536), .C2(new_n511), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n509), .A2(new_n531), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G229gat), .A2(G233gat), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n529), .A2(new_n530), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n505), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n509), .A2(new_n531), .A3(KEYINPUT94), .A4(new_n537), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n540), .A2(new_n541), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT18), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n542), .B(new_n505), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n541), .B(KEYINPUT13), .Z(new_n548));
  AOI22_X1  g347(.A1(new_n545), .A2(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n544), .A2(new_n543), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n550), .A2(KEYINPUT18), .A3(new_n541), .A4(new_n540), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G113gat), .B(G141gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(G197gat), .ZN(new_n554));
  XOR2_X1   g353(.A(KEYINPUT11), .B(G169gat), .Z(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT12), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n549), .A2(new_n557), .A3(new_n551), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n491), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G71gat), .A2(G78gat), .ZN(new_n564));
  INV_X1    g363(.A(G71gat), .ZN(new_n565));
  INV_X1    g364(.A(G78gat), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT9), .ZN(new_n567));
  INV_X1    g366(.A(G64gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n568), .A2(G57gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n564), .A2(new_n567), .B1(new_n569), .B2(KEYINPUT95), .ZN(new_n570));
  INV_X1    g369(.A(G57gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(G64gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n568), .A2(G57gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT95), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n573), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT9), .ZN(new_n577));
  AND2_X1   g376(.A1(G71gat), .A2(G78gat), .ZN(new_n578));
  NOR2_X1   g377(.A1(G71gat), .A2(G78gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n570), .A2(new_n575), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n581), .A2(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n582), .B(new_n583), .Z(new_n584));
  XOR2_X1   g383(.A(G127gat), .B(G155gat), .Z(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT96), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n584), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G183gat), .B(G211gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n505), .B1(KEYINPUT21), .B2(new_n581), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n589), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT8), .ZN(new_n596));
  NAND2_X1  g395(.A1(G85gat), .A2(G92gat), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT7), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(G85gat), .ZN(new_n600));
  INV_X1    g399(.A(G92gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n596), .A2(new_n599), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G99gat), .B(G106gat), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n607), .A2(KEYINPUT98), .ZN(new_n608));
  AND3_X1   g407(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI22_X1  g410(.A1(KEYINPUT8), .A2(new_n595), .B1(new_n600), .B2(new_n601), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(new_n605), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n607), .A2(KEYINPUT98), .A3(new_n613), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n531), .A2(new_n537), .A3(new_n608), .A4(new_n614), .ZN(new_n615));
  AND3_X1   g414(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n608), .A2(new_n614), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n616), .B1(new_n542), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G190gat), .B(G218gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n615), .A2(new_n618), .A3(new_n620), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n622), .A2(KEYINPUT97), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT99), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(G134gat), .B(G162gat), .Z(new_n627));
  AOI21_X1  g426(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n626), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n622), .A2(new_n623), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n629), .B1(new_n632), .B2(KEYINPUT99), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n630), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n594), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n567), .A2(new_n564), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n569), .A2(KEYINPUT95), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n575), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G57gat), .B(G64gat), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT9), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n580), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n608), .A2(new_n643), .A3(new_n614), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n604), .A2(new_n606), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n605), .B1(new_n611), .B2(new_n612), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT100), .B1(new_n647), .B2(new_n581), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n607), .A2(new_n639), .A3(new_n613), .A4(new_n642), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT100), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n644), .B1(new_n648), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G230gat), .A2(G233gat), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n656), .B(new_n657), .Z(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT10), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n662), .B(new_n644), .C1(new_n648), .C2(new_n651), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n617), .A2(KEYINPUT10), .A3(new_n581), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(KEYINPUT101), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n663), .A2(new_n667), .A3(new_n664), .ZN(new_n668));
  AND4_X1   g467(.A1(new_n661), .A2(new_n666), .A3(new_n653), .A4(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n654), .B1(new_n665), .B2(KEYINPUT101), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n661), .B1(new_n670), .B2(new_n668), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n660), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n665), .A2(new_n653), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n665), .A2(KEYINPUT103), .A3(new_n653), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n659), .B1(new_n677), .B2(new_n655), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n636), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n563), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(new_n437), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(new_n492), .ZN(G1324gat));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684));
  INV_X1    g483(.A(new_n486), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT16), .B(G8gat), .Z(new_n687));
  AOI21_X1  g486(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(G8gat), .B1(new_n681), .B2(new_n685), .ZN(new_n689));
  NOR2_X1   g488(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n690));
  MUX2_X1   g489(.A(KEYINPUT104), .B(new_n690), .S(new_n687), .Z(new_n691));
  AOI22_X1  g490(.A1(new_n688), .A2(new_n689), .B1(new_n686), .B2(new_n691), .ZN(G1325gat));
  NAND2_X1  g491(.A1(new_n459), .A2(G15gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT106), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n681), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n494), .B1(new_n681), .B2(new_n274), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n695), .B1(new_n698), .B2(new_n699), .ZN(G1326gat));
  NAND3_X1  g499(.A1(new_n563), .A2(new_n460), .A3(new_n680), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n701), .A2(KEYINPUT107), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(KEYINPUT107), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT43), .B(G22gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  NOR2_X1   g505(.A1(new_n491), .A2(new_n635), .ZN(new_n707));
  INV_X1    g506(.A(new_n437), .ZN(new_n708));
  INV_X1    g507(.A(new_n594), .ZN(new_n709));
  INV_X1    g508(.A(new_n679), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n562), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n707), .A2(new_n526), .A3(new_n708), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT45), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n715), .B1(new_n491), .B2(new_n635), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n461), .A2(new_n490), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n399), .A2(new_n402), .A3(KEYINPUT79), .ZN(new_n718));
  AOI21_X1  g517(.A(KEYINPUT79), .B1(new_n399), .B2(new_n402), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI22_X1  g519(.A1(new_n435), .A2(new_n436), .B1(new_n438), .B2(new_n400), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n489), .A2(new_n720), .A3(new_n275), .A4(new_n721), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n722), .A2(KEYINPUT35), .B1(new_n447), .B2(new_n455), .ZN(new_n723));
  OAI211_X1 g522(.A(KEYINPUT44), .B(new_n634), .C1(new_n717), .C2(new_n723), .ZN(new_n724));
  AND4_X1   g523(.A1(new_n708), .A2(new_n716), .A3(new_n712), .A4(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n714), .B1(new_n526), .B2(new_n725), .ZN(G1328gat));
  NAND4_X1  g525(.A1(new_n707), .A2(new_n524), .A3(new_n486), .A4(new_n712), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n727), .A2(KEYINPUT46), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n716), .A2(new_n724), .A3(new_n712), .ZN(new_n729));
  OAI21_X1  g528(.A(G36gat), .B1(new_n729), .B2(new_n685), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n727), .A2(KEYINPUT46), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n728), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT108), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n728), .A2(new_n730), .A3(new_n734), .A4(new_n731), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(G1329gat));
  NAND3_X1  g535(.A1(new_n707), .A2(new_n275), .A3(new_n712), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n260), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n459), .A2(G43gat), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n729), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g540(.A(new_n534), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n729), .B2(new_n489), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n711), .A2(new_n742), .A3(new_n635), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n563), .A2(new_n460), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT48), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n746), .B(new_n748), .ZN(G1331gat));
  NAND2_X1  g548(.A1(new_n442), .A2(new_n456), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n461), .A2(new_n490), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n636), .A2(new_n710), .A3(new_n561), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n437), .ZN(new_n755));
  XOR2_X1   g554(.A(KEYINPUT110), .B(G57gat), .Z(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(G1332gat));
  NOR2_X1   g556(.A1(new_n754), .A2(new_n685), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  AND2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n758), .B2(new_n759), .ZN(G1333gat));
  INV_X1    g561(.A(new_n459), .ZN(new_n763));
  OAI21_X1  g562(.A(G71gat), .B1(new_n754), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n275), .A2(new_n565), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n754), .B2(new_n765), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g566(.A1(new_n754), .A2(new_n489), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(new_n566), .ZN(G1335gat));
  NOR2_X1   g568(.A1(new_n594), .A2(new_n561), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n634), .B(new_n770), .C1(new_n717), .C2(new_n723), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT51), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n752), .A2(new_n634), .A3(new_n770), .A4(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n710), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n778), .A2(new_n600), .A3(new_n708), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n770), .A2(new_n679), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT111), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n716), .A2(new_n724), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n716), .A2(new_n724), .A3(KEYINPUT112), .A4(new_n781), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n784), .A2(new_n708), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n779), .B1(new_n786), .B2(new_n600), .ZN(G1336gat));
  NAND2_X1  g586(.A1(new_n774), .A2(new_n777), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n685), .A2(G92gat), .A3(new_n710), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(G92gat), .B1(new_n782), .B2(new_n685), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n789), .B(KEYINPUT114), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(new_n774), .B2(new_n777), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n784), .A2(new_n486), .A3(new_n785), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n796), .B2(G92gat), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n793), .B1(new_n797), .B2(new_n792), .ZN(G1337gat));
  INV_X1    g597(.A(G99gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n778), .A2(new_n799), .A3(new_n275), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n784), .A2(new_n459), .A3(new_n785), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n801), .B2(new_n799), .ZN(G1338gat));
  NOR2_X1   g601(.A1(new_n489), .A2(G106gat), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n778), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805));
  OAI21_X1  g604(.A(G106gat), .B1(new_n782), .B2(new_n489), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n803), .ZN(new_n808));
  AOI211_X1 g607(.A(new_n710), .B(new_n808), .C1(new_n774), .C2(new_n777), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n784), .A2(new_n460), .A3(new_n785), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n809), .B1(new_n810), .B2(G106gat), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n807), .B1(new_n811), .B2(new_n805), .ZN(G1339gat));
  NAND3_X1  g611(.A1(new_n666), .A2(new_n653), .A3(new_n668), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT102), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n670), .A2(new_n661), .A3(new_n668), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI22_X1  g615(.A1(new_n559), .A2(new_n560), .B1(new_n816), .B2(new_n660), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n663), .A2(new_n654), .A3(new_n664), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT54), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n820), .B1(new_n814), .B2(new_n815), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT103), .B1(new_n665), .B2(new_n653), .ZN(new_n823));
  AOI211_X1 g622(.A(new_n674), .B(new_n654), .C1(new_n663), .C2(new_n664), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n659), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n818), .B1(new_n821), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(KEYINPUT55), .A3(new_n659), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n821), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n825), .A2(KEYINPUT55), .A3(new_n659), .ZN(new_n831));
  INV_X1    g630(.A(new_n820), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n832), .B1(new_n669), .B2(new_n671), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT115), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n817), .B(new_n827), .C1(new_n830), .C2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n541), .B1(new_n550), .B2(new_n540), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n547), .A2(new_n548), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n556), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n560), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n679), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n634), .B1(new_n835), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n634), .A2(new_n827), .A3(new_n840), .A4(new_n672), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n830), .A2(new_n834), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n709), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n636), .A2(new_n561), .A3(new_n679), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n489), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n708), .A2(new_n275), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n850), .A2(new_n486), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(G113gat), .B1(new_n852), .B2(new_n561), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n852), .B(KEYINPUT116), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n561), .A2(G113gat), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(G1340gat));
  AOI21_X1  g655(.A(G120gat), .B1(new_n852), .B2(new_n679), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n679), .A2(G120gat), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n854), .B2(new_n858), .ZN(G1341gat));
  INV_X1    g658(.A(G127gat), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n852), .A2(new_n860), .A3(new_n594), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n854), .A2(new_n594), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n861), .B1(new_n862), .B2(new_n860), .ZN(G1342gat));
  NOR2_X1   g662(.A1(new_n635), .A2(new_n486), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT117), .ZN(new_n865));
  NOR4_X1   g664(.A1(new_n850), .A2(G134gat), .A3(new_n851), .A4(new_n865), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT56), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n854), .A2(new_n634), .ZN(new_n868));
  INV_X1    g667(.A(G134gat), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(G1343gat));
  NOR3_X1   g669(.A1(new_n459), .A2(new_n437), .A3(new_n486), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n460), .A2(KEYINPUT57), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n843), .A2(new_n844), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT118), .B1(new_n821), .B2(new_n826), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n658), .B1(new_n677), .B2(new_n822), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n833), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n874), .A2(new_n818), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n829), .B1(new_n821), .B2(new_n828), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n831), .A2(new_n833), .A3(KEYINPUT115), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n878), .A2(new_n881), .A3(new_n817), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n634), .B1(new_n882), .B2(new_n841), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n873), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n841), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n549), .A2(new_n557), .A3(new_n551), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n557), .B1(new_n549), .B2(new_n551), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n672), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n889), .B1(new_n879), .B2(new_n880), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n886), .B1(new_n890), .B2(new_n878), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n891), .A2(KEYINPUT119), .A3(new_n634), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n709), .B1(new_n885), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n872), .B1(new_n893), .B2(new_n848), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n489), .B1(new_n846), .B2(new_n848), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(KEYINPUT57), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n871), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(G141gat), .B1(new_n897), .B2(new_n562), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n895), .A2(new_n871), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n561), .A2(new_n297), .ZN(new_n900));
  XOR2_X1   g699(.A(new_n900), .B(KEYINPUT120), .Z(new_n901));
  AOI21_X1  g700(.A(KEYINPUT121), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT58), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT58), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n898), .A2(new_n905), .A3(new_n902), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(G1344gat));
  OAI211_X1 g706(.A(new_n679), .B(new_n871), .C1(new_n894), .C2(new_n896), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n293), .A2(KEYINPUT59), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT57), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n873), .B1(new_n891), .B2(new_n634), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n847), .B1(new_n912), .B2(new_n709), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n460), .A2(new_n911), .ZN(new_n914));
  OAI22_X1  g713(.A1(new_n895), .A2(new_n911), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n871), .A2(new_n679), .ZN(new_n916));
  OAI21_X1  g715(.A(G148gat), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g716(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n910), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n899), .A2(new_n293), .A3(new_n679), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AOI22_X1  g722(.A1(new_n908), .A2(new_n909), .B1(new_n917), .B2(new_n918), .ZN(new_n924));
  INV_X1    g723(.A(new_n922), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT123), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n923), .A2(new_n926), .ZN(G1345gat));
  OAI21_X1  g726(.A(new_n290), .B1(new_n897), .B2(new_n709), .ZN(new_n928));
  INV_X1    g727(.A(new_n290), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n899), .A2(new_n929), .A3(new_n594), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1346gat));
  OAI21_X1  g730(.A(G162gat), .B1(new_n897), .B2(new_n635), .ZN(new_n932));
  INV_X1    g731(.A(new_n895), .ZN(new_n933));
  OR4_X1    g732(.A1(G162gat), .A2(new_n865), .A3(new_n437), .A4(new_n459), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(G1347gat));
  NOR2_X1   g734(.A1(new_n708), .A2(new_n685), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n275), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n850), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(G169gat), .B1(new_n938), .B2(new_n561), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n460), .B1(new_n846), .B2(new_n848), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n937), .B(KEYINPUT124), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n941), .B1(new_n942), .B2(new_n940), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n562), .A2(new_n202), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n939), .B1(new_n945), .B2(new_n946), .ZN(G1348gat));
  NAND3_X1  g746(.A1(new_n938), .A2(new_n203), .A3(new_n679), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n943), .A2(new_n944), .A3(new_n710), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(new_n203), .ZN(G1349gat));
  AND2_X1   g749(.A1(new_n594), .A2(new_n223), .ZN(new_n951));
  AOI21_X1  g750(.A(KEYINPUT126), .B1(new_n938), .B2(new_n951), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n943), .A2(new_n944), .A3(new_n709), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n953), .B2(new_n211), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT60), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT60), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n956), .B(new_n952), .C1(new_n953), .C2(new_n211), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(G1350gat));
  NAND3_X1  g757(.A1(new_n938), .A2(new_n224), .A3(new_n634), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n634), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n960), .B1(new_n961), .B2(G190gat), .ZN(new_n962));
  AOI211_X1 g761(.A(KEYINPUT61), .B(new_n224), .C1(new_n945), .C2(new_n634), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(G1351gat));
  NAND2_X1  g763(.A1(new_n763), .A2(new_n936), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n933), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g765(.A(G197gat), .B1(new_n966), .B2(new_n561), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n915), .A2(new_n965), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n561), .A2(G197gat), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(G1352gat));
  NOR4_X1   g769(.A1(new_n933), .A2(G204gat), .A3(new_n710), .A4(new_n965), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT62), .ZN(new_n972));
  INV_X1    g771(.A(new_n968), .ZN(new_n973));
  OAI21_X1  g772(.A(G204gat), .B1(new_n973), .B2(new_n710), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n974), .ZN(G1353gat));
  INV_X1    g774(.A(G211gat), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n966), .A2(new_n976), .A3(new_n594), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n968), .A2(new_n594), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n978), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n979));
  AOI21_X1  g778(.A(KEYINPUT63), .B1(new_n978), .B2(G211gat), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(G1354gat));
  AOI21_X1  g780(.A(G218gat), .B1(new_n966), .B2(new_n634), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n968), .A2(KEYINPUT127), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n634), .A2(new_n279), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n984), .B1(new_n968), .B2(KEYINPUT127), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n982), .B1(new_n983), .B2(new_n985), .ZN(G1355gat));
endmodule


