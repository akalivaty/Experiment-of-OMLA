//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n563, new_n565, new_n566, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n621, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1240, new_n1241, new_n1242, new_n1243;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n454), .A2(new_n458), .B1(new_n459), .B2(new_n455), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT69), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT3), .ZN(new_n466));
  OR2_X1    g041(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(G137), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(new_n465), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT68), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n472), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n471), .A2(new_n477), .ZN(G160));
  AND3_X1   g053(.A1(new_n466), .A2(KEYINPUT70), .A3(new_n467), .ZN(new_n479));
  AOI21_X1  g054(.A(KEYINPUT70), .B1(new_n466), .B2(new_n467), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n472), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n472), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI22_X1  g059(.A1(new_n481), .A2(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(G2105), .B1(new_n479), .B2(new_n480), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(KEYINPUT71), .B(G2105), .C1(new_n479), .C2(new_n480), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n485), .B1(new_n490), .B2(G124), .ZN(G162));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n472), .A2(G138), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n473), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n466), .A2(new_n467), .A3(new_n493), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT72), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n496), .A2(new_n499), .A3(KEYINPUT4), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n495), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n466), .A2(G126), .A3(G2105), .A4(new_n467), .ZN(new_n502));
  OR2_X1    g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n503), .B(G2104), .C1(G114), .C2(new_n472), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n501), .A2(new_n505), .ZN(G164));
  XNOR2_X1  g081(.A(KEYINPUT5), .B(G543), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n507), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n511));
  XOR2_X1   g086(.A(KEYINPUT6), .B(G651), .Z(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n510), .A2(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  INV_X1    g090(.A(new_n507), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n507), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n517), .A2(G63), .A3(G651), .A4(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n512), .A2(KEYINPUT74), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT6), .B(G651), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT74), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n521), .A2(G543), .A3(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n520), .B(KEYINPUT75), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT76), .B(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n528), .B(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n516), .A2(new_n512), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n530), .B1(G89), .B2(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n520), .B1(new_n525), .B2(new_n526), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT75), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n533), .A2(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  NAND2_X1  g113(.A1(new_n517), .A2(new_n519), .ZN(new_n539));
  INV_X1    g114(.A(G64), .ZN(new_n540));
  INV_X1    g115(.A(G77), .ZN(new_n541));
  INV_X1    g116(.A(G543), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n539), .A2(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT77), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI221_X1 g120(.A(KEYINPUT77), .B1(new_n541), .B2(new_n542), .C1(new_n539), .C2(new_n540), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n545), .A2(G651), .A3(new_n546), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n521), .A2(G543), .A3(new_n524), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n548), .A2(G52), .B1(G90), .B2(new_n531), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n539), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G651), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n521), .A2(G43), .A3(G543), .A4(new_n524), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n531), .A2(G81), .ZN(new_n557));
  AND3_X1   g132(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT78), .ZN(new_n558));
  AOI21_X1  g133(.A(KEYINPUT78), .B1(new_n556), .B2(new_n557), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n555), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  AND3_X1   g137(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G36), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n563), .A2(new_n566), .ZN(G188));
  INV_X1    g142(.A(G53), .ZN(new_n568));
  OR3_X1    g143(.A1(new_n525), .A2(KEYINPUT9), .A3(new_n568), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT9), .B1(new_n525), .B2(new_n568), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n516), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n574), .A2(G651), .B1(new_n531), .B2(G91), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n571), .A2(new_n575), .ZN(G299));
  NAND2_X1  g151(.A1(new_n548), .A2(G49), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n507), .B(KEYINPUT73), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n578), .B2(G74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n531), .A2(G87), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(G288));
  AOI22_X1  g156(.A1(new_n507), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n512), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n507), .A2(G61), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT79), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n509), .B1(new_n584), .B2(new_n585), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT79), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n583), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G305));
  NAND2_X1  g168(.A1(new_n531), .A2(G85), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n525), .B2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G72), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G60), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n539), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n509), .B1(new_n600), .B2(KEYINPUT80), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT80), .ZN(new_n602));
  OAI211_X1 g177(.A(new_n602), .B(new_n598), .C1(new_n539), .C2(new_n599), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n601), .A2(KEYINPUT81), .A3(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(KEYINPUT81), .B1(new_n601), .B2(new_n603), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n597), .B1(new_n605), .B2(new_n606), .ZN(G290));
  AOI22_X1  g182(.A1(new_n507), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(new_n509), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(new_n548), .B2(G54), .ZN(new_n610));
  AND3_X1   g185(.A1(new_n507), .A2(new_n522), .A3(G92), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G171), .B2(new_n614), .ZN(G284));
  OAI21_X1  g191(.A(new_n615), .B1(G171), .B2(new_n614), .ZN(G321));
  NAND2_X1  g192(.A1(G299), .A2(new_n614), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G168), .B2(new_n614), .ZN(G280));
  XOR2_X1   g194(.A(G280), .B(KEYINPUT82), .Z(G297));
  AND2_X1   g195(.A1(new_n610), .A2(new_n612), .ZN(new_n621));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT83), .ZN(new_n625));
  MUX2_X1   g200(.A(new_n560), .B(new_n625), .S(G868), .Z(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g202(.A(G135), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n472), .A2(G111), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  OAI22_X1  g205(.A1(new_n481), .A2(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(new_n490), .B2(G123), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(KEYINPUT86), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(KEYINPUT86), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n635), .A2(G2096), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(G2096), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n469), .A2(new_n473), .A3(new_n472), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT12), .Z(new_n639));
  XOR2_X1   g214(.A(KEYINPUT84), .B(KEYINPUT13), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT85), .B(G2100), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n636), .A2(new_n637), .A3(new_n643), .ZN(G156));
  INV_X1    g219(.A(KEYINPUT14), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(new_n648), .B2(new_n647), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n650), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  AND3_X1   g233(.A1(new_n657), .A2(G14), .A3(new_n658), .ZN(G401));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  NAND3_X1  g238(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT18), .Z(new_n665));
  INV_X1    g240(.A(new_n662), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n663), .B1(new_n666), .B2(new_n660), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n667), .A2(KEYINPUT87), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(KEYINPUT87), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n660), .B(KEYINPUT17), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n668), .B(new_n669), .C1(new_n666), .C2(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(new_n666), .A3(new_n663), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n665), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2096), .B(G2100), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(G1971), .B(G1976), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n677), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n677), .A2(new_n680), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT20), .Z(new_n684));
  AOI211_X1 g259(.A(new_n682), .B(new_n684), .C1(new_n677), .C2(new_n681), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT88), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1991), .B(G1996), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n692), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(G229));
  XNOR2_X1  g270(.A(KEYINPUT27), .B(G1996), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT97), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT26), .Z(new_n700));
  NAND3_X1  g275(.A1(new_n469), .A2(G105), .A3(new_n472), .ZN(new_n701));
  INV_X1    g276(.A(G141), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n700), .B(new_n701), .C1(new_n481), .C2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n490), .B2(G129), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT96), .Z(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G29), .ZN(new_n706));
  OR2_X1    g281(.A1(G29), .A2(G32), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n698), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n696), .A2(new_n697), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n708), .B(new_n709), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n621), .A2(G16), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G4), .B2(G16), .ZN(new_n712));
  INV_X1    g287(.A(G1348), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT31), .B(G11), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT30), .B(G28), .Z(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(G29), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n712), .B2(new_n713), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NOR2_X1   g294(.A1(G171), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G5), .B2(new_n719), .ZN(new_n721));
  INV_X1    g296(.A(G1961), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n714), .B(new_n718), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G33), .ZN(new_n725));
  INV_X1    g300(.A(new_n481), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G139), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n473), .A2(G127), .ZN(new_n728));
  INV_X1    g303(.A(G115), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n462), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT25), .ZN(new_n731));
  NAND2_X1  g306(.A1(G103), .A2(G2104), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(G2105), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n472), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n730), .A2(G2105), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n727), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n725), .B1(new_n737), .B2(new_n724), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(G2072), .Z(new_n739));
  INV_X1    g314(.A(G160), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT24), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n741), .A2(G34), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n724), .B1(new_n741), .B2(G34), .ZN(new_n743));
  OAI22_X1  g318(.A1(new_n740), .A2(new_n724), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G2084), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n739), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n723), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n635), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G29), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n724), .A2(G35), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G162), .B2(new_n724), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT29), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n747), .B(new_n749), .C1(G2090), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n724), .A2(G27), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G164), .B2(new_n724), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G2078), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n719), .A2(G19), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n561), .B2(new_n719), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n758), .A2(G1341), .ZN(new_n759));
  AOI211_X1 g334(.A(new_n756), .B(new_n759), .C1(new_n721), .C2(new_n722), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n724), .A2(G26), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT28), .ZN(new_n762));
  INV_X1    g337(.A(G128), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n488), .B2(new_n489), .ZN(new_n764));
  OAI21_X1  g339(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n765));
  INV_X1    g340(.A(G116), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n765), .B1(new_n766), .B2(G2105), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G140), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n481), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n764), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n762), .B1(new_n771), .B2(new_n724), .ZN(new_n772));
  INV_X1    g347(.A(G2067), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n758), .A2(G1341), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n719), .A2(G21), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G168), .B2(new_n719), .ZN(new_n777));
  INV_X1    g352(.A(G1966), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n760), .A2(new_n774), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  NOR3_X1   g355(.A1(new_n710), .A2(new_n753), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n752), .A2(G2090), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT98), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n719), .A2(G20), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT23), .Z(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G299), .B2(G16), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT99), .ZN(new_n787));
  INV_X1    g362(.A(G1956), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n783), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(KEYINPUT100), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT100), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n783), .A2(new_n792), .A3(new_n789), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n781), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n719), .A2(G22), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G166), .B2(new_n719), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1971), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n719), .A2(G23), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G288), .B2(G16), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT93), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT33), .B(G1976), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n797), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n804), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n801), .B2(new_n802), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n719), .A2(G6), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n592), .B2(new_n719), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT92), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT32), .B(G1981), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(KEYINPUT94), .B1(new_n808), .B2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n812), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n811), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT94), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n816), .A2(new_n817), .A3(new_n807), .A4(new_n805), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n814), .A2(KEYINPUT34), .A3(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT95), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n814), .A2(new_n818), .A3(KEYINPUT95), .A4(KEYINPUT34), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(KEYINPUT34), .B1(new_n814), .B2(new_n818), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n719), .A2(G24), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n603), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT81), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n596), .B1(new_n828), .B2(new_n604), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n825), .B1(new_n829), .B2(new_n719), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(G1986), .Z(new_n831));
  OR2_X1    g406(.A1(G25), .A2(G29), .ZN(new_n832));
  OAI21_X1  g407(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n833));
  INV_X1    g408(.A(G107), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(G2105), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n726), .B2(G131), .ZN(new_n836));
  AOI21_X1  g411(.A(KEYINPUT89), .B1(new_n490), .B2(G119), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT89), .ZN(new_n838));
  INV_X1    g413(.A(G119), .ZN(new_n839));
  AOI211_X1 g414(.A(new_n838), .B(new_n839), .C1(new_n488), .C2(new_n489), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n836), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n832), .B1(new_n841), .B2(new_n724), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT35), .B(G1991), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT91), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT90), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n842), .A2(new_n845), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n831), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n824), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n823), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(KEYINPUT36), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT36), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n823), .A2(new_n852), .A3(new_n849), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n794), .B1(new_n851), .B2(new_n853), .ZN(G311));
  NAND2_X1  g429(.A1(new_n851), .A2(new_n853), .ZN(new_n855));
  INV_X1    g430(.A(new_n794), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(G150));
  NAND2_X1  g432(.A1(new_n621), .A2(G559), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT38), .ZN(new_n859));
  INV_X1    g434(.A(G55), .ZN(new_n860));
  INV_X1    g435(.A(new_n531), .ZN(new_n861));
  XNOR2_X1  g436(.A(KEYINPUT101), .B(G93), .ZN(new_n862));
  OAI22_X1  g437(.A1(new_n525), .A2(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n517), .A2(G67), .A3(new_n519), .ZN(new_n864));
  NAND2_X1  g439(.A1(G80), .A2(G543), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n509), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(new_n560), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n867), .B(new_n555), .C1(new_n559), .C2(new_n558), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n859), .B(new_n871), .Z(new_n872));
  AND2_X1   g447(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n873), .A2(new_n874), .A3(G860), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n868), .A2(G860), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT102), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(KEYINPUT37), .Z(new_n878));
  OR2_X1    g453(.A1(new_n875), .A2(new_n878), .ZN(G145));
  NAND2_X1  g454(.A1(new_n704), .A2(new_n736), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(new_n705), .B2(new_n736), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n841), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n466), .A2(new_n467), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT70), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n466), .A2(KEYINPUT70), .A3(new_n467), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT71), .B1(new_n889), .B2(G2105), .ZN(new_n890));
  INV_X1    g465(.A(new_n489), .ZN(new_n891));
  OAI21_X1  g466(.A(G119), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n838), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n490), .A2(KEYINPUT89), .A3(G119), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n895), .A2(KEYINPUT105), .A3(new_n836), .ZN(new_n896));
  INV_X1    g471(.A(new_n639), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n884), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n897), .B1(new_n884), .B2(new_n896), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n496), .A2(new_n499), .A3(KEYINPUT4), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n499), .B1(new_n496), .B2(KEYINPUT4), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n494), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n502), .A2(KEYINPUT103), .A3(new_n504), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT103), .B1(new_n502), .B2(new_n504), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n902), .B(new_n905), .C1(new_n764), .C2(new_n770), .ZN(new_n906));
  OAI21_X1  g481(.A(G128), .B1(new_n890), .B2(new_n891), .ZN(new_n907));
  INV_X1    g482(.A(new_n770), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n902), .A2(new_n905), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n490), .A2(G130), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n490), .A2(KEYINPUT104), .A3(G130), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n917));
  INV_X1    g492(.A(G118), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n917), .B1(new_n918), .B2(G2105), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n919), .B1(new_n726), .B2(G142), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n911), .A2(new_n916), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT104), .B1(new_n490), .B2(G130), .ZN(new_n922));
  INV_X1    g497(.A(G130), .ZN(new_n923));
  AOI211_X1 g498(.A(new_n913), .B(new_n923), .C1(new_n488), .C2(new_n489), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n920), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n925), .A2(new_n910), .A3(new_n906), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n921), .A2(new_n926), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n898), .A2(new_n899), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT105), .B1(new_n895), .B2(new_n836), .ZN(new_n929));
  INV_X1    g504(.A(new_n836), .ZN(new_n930));
  AOI211_X1 g505(.A(new_n883), .B(new_n930), .C1(new_n893), .C2(new_n894), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n639), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n884), .A2(new_n896), .A3(new_n897), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n932), .A2(new_n933), .B1(new_n926), .B2(new_n921), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n882), .B1(new_n928), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n635), .B(new_n740), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(G162), .ZN(new_n937));
  INV_X1    g512(.A(G162), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n748), .A2(new_n740), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n635), .A2(G160), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n927), .B1(new_n898), .B2(new_n899), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n932), .A2(new_n933), .A3(new_n926), .A4(new_n921), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(new_n944), .A3(new_n881), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n935), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n935), .A2(KEYINPUT106), .A3(new_n942), .A4(new_n945), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n942), .B1(new_n935), .B2(new_n945), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(G37), .ZN(new_n952));
  XNOR2_X1  g527(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n950), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n953), .B1(new_n950), .B2(new_n952), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(G395));
  NOR2_X1   g531(.A1(new_n868), .A2(G868), .ZN(new_n957));
  XNOR2_X1  g532(.A(G288), .B(G303), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n829), .A2(G305), .ZN(new_n960));
  AOI211_X1 g535(.A(new_n592), .B(new_n596), .C1(new_n828), .C2(new_n604), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(G290), .A2(new_n592), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n829), .A2(G305), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(new_n964), .A3(new_n958), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT42), .ZN(new_n967));
  OR3_X1    g542(.A1(new_n966), .A2(KEYINPUT111), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n967), .B1(new_n966), .B2(KEYINPUT111), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT112), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n968), .A2(KEYINPUT112), .A3(new_n969), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n974));
  XOR2_X1   g549(.A(new_n625), .B(new_n871), .Z(new_n975));
  NAND2_X1  g550(.A1(G299), .A2(new_n613), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n621), .A2(new_n571), .A3(new_n575), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(KEYINPUT109), .B(KEYINPUT41), .Z(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(new_n978), .B2(KEYINPUT41), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n974), .B1(new_n975), .B2(new_n982), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n976), .A2(KEYINPUT108), .A3(new_n977), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT108), .B1(new_n976), .B2(new_n977), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n983), .B1(new_n975), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n975), .A2(new_n974), .A3(new_n982), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n972), .A2(new_n973), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n987), .A2(new_n988), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n990), .A2(new_n971), .A3(new_n970), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n957), .B1(new_n992), .B2(G868), .ZN(G295));
  AOI21_X1  g568(.A(new_n957), .B1(new_n992), .B2(G868), .ZN(G331));
  NAND4_X1  g569(.A1(new_n547), .A2(new_n533), .A3(new_n536), .A4(new_n549), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n547), .A2(new_n549), .B1(new_n533), .B2(new_n536), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n871), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(G301), .A2(G286), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n999), .A2(new_n869), .A3(new_n870), .A4(new_n995), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n998), .A2(KEYINPUT114), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n871), .B(new_n1002), .C1(new_n996), .C2(new_n997), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(new_n982), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n978), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n998), .A2(new_n1005), .A3(new_n1000), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n966), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n966), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1011));
  INV_X1    g586(.A(G37), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT43), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n998), .A2(new_n1000), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1005), .A2(new_n980), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1015), .B(new_n1016), .C1(KEYINPUT41), .C2(new_n1005), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n986), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI211_X1 g595(.A(KEYINPUT115), .B(new_n986), .C1(new_n1001), .C2(new_n1003), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1008), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1014), .B1(new_n1024), .B2(KEYINPUT43), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT113), .B(KEYINPUT44), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1024), .A2(KEYINPUT43), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT43), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1009), .A2(new_n1030), .A3(new_n1012), .A4(new_n1011), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1031), .A2(KEYINPUT44), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1028), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1030), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1031), .A2(KEYINPUT44), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1034), .A2(new_n1035), .A3(KEYINPUT116), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1027), .B1(new_n1033), .B2(new_n1036), .ZN(G397));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n1038));
  INV_X1    g613(.A(G40), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n471), .A2(new_n1039), .A3(new_n477), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1384), .B1(new_n902), .B2(new_n905), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(KEYINPUT45), .ZN(new_n1042));
  INV_X1    g617(.A(G1384), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1043), .B1(new_n501), .B2(new_n505), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT45), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1038), .B(new_n778), .C1(new_n1042), .C2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1040), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT50), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1048), .B1(new_n1041), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1044), .A2(KEYINPUT50), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1047), .B1(G2084), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n909), .A2(new_n1043), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1048), .B1(new_n1054), .B2(new_n1045), .ZN(new_n1055));
  INV_X1    g630(.A(new_n505), .ZN(new_n1056));
  AOI21_X1  g631(.A(G1384), .B1(new_n902), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT45), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1038), .B1(new_n1059), .B2(new_n778), .ZN(new_n1060));
  OAI21_X1  g635(.A(G8), .B1(new_n1053), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G8), .ZN(new_n1062));
  NOR2_X1   g637(.A1(G168), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT51), .B1(new_n1064), .B2(KEYINPUT124), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1061), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1052), .A2(G2084), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n778), .B1(new_n1042), .B2(new_n1046), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT119), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(new_n1070), .A3(new_n1047), .ZN(new_n1071));
  OAI211_X1 g646(.A(G8), .B(new_n1065), .C1(new_n1071), .C2(G286), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1063), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1067), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT62), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT125), .B(KEYINPUT53), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT103), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n505), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n502), .A2(KEYINPUT103), .A3(new_n504), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g655(.A(KEYINPUT45), .B(new_n1043), .C1(new_n501), .C2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1081), .B(new_n1040), .C1(KEYINPUT45), .C2(new_n1057), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1076), .B1(new_n1082), .B2(G2078), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT126), .ZN(new_n1084));
  XNOR2_X1  g659(.A(new_n1083), .B(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1052), .A2(new_n722), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1087), .A2(G2078), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1055), .A2(new_n1058), .A3(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1085), .A2(new_n1086), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(G303), .A2(G8), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1091), .B(KEYINPUT55), .ZN(new_n1092));
  INV_X1    g667(.A(G1971), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1082), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1054), .A2(KEYINPUT50), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1048), .B1(new_n1057), .B2(new_n1049), .ZN(new_n1096));
  INV_X1    g671(.A(G2090), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1092), .B1(new_n1099), .B2(new_n1062), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1050), .A2(new_n1097), .A3(new_n1051), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1062), .B1(new_n1094), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1092), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1043), .B(new_n1040), .C1(new_n501), .C2(new_n1080), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1106), .A2(new_n1062), .ZN(new_n1107));
  OAI21_X1  g682(.A(G1981), .B1(new_n583), .B2(new_n589), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(G305), .B2(G1981), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT49), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(KEYINPUT49), .B(new_n1108), .C1(G305), .C2(G1981), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1107), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G288), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(G1976), .ZN(new_n1115));
  INV_X1    g690(.A(G1976), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT52), .B1(G288), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1107), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1115), .A2(G8), .A3(new_n1105), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT52), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1113), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1100), .A2(new_n1104), .A3(new_n1122), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1090), .A2(new_n1123), .A3(G301), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1067), .A2(new_n1072), .A3(new_n1125), .A4(new_n1073), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1075), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1113), .A2(new_n1116), .A3(new_n1114), .ZN(new_n1128));
  NOR2_X1   g703(.A1(G305), .A2(G1981), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1107), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n1104), .B2(new_n1121), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1071), .A2(G8), .A3(G168), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1122), .B(new_n1134), .C1(new_n1103), .C2(new_n1102), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT63), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1136), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT120), .B1(new_n1138), .B2(new_n1121), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1133), .A2(new_n1135), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1136), .B1(new_n1123), .B2(new_n1132), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1131), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  XOR2_X1   g717(.A(G299), .B(KEYINPUT57), .Z(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(KEYINPUT56), .B(G2072), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT121), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT122), .B1(new_n1082), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1048), .B1(new_n1041), .B2(KEYINPUT45), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1146), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1049), .B(new_n1043), .C1(new_n501), .C2(new_n505), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n1040), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1049), .B1(new_n909), .B2(new_n1043), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n788), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1153), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1144), .B1(new_n1148), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n1160));
  AOI21_X1  g735(.A(G1348), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1105), .A2(G2067), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1049), .B(new_n1043), .C1(new_n501), .C2(new_n1080), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1040), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1057), .A2(new_n1049), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n713), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1162), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1167), .A2(KEYINPUT123), .A3(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1163), .A2(new_n621), .A3(new_n1169), .ZN(new_n1170));
  AND4_X1   g745(.A1(new_n1143), .A2(new_n1147), .A3(new_n1153), .A4(new_n1157), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1159), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n1153), .A2(new_n1157), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1143), .B1(new_n1174), .B2(new_n1147), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1173), .B1(new_n1175), .B2(new_n1171), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n1161), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1177));
  AOI21_X1  g752(.A(KEYINPUT123), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT60), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT60), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1163), .A2(new_n1180), .A3(new_n1169), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1179), .A2(new_n621), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1174), .A2(new_n1143), .A3(new_n1147), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1183), .A2(new_n1159), .A3(KEYINPUT61), .ZN(new_n1184));
  AND3_X1   g759(.A1(new_n1176), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(KEYINPUT58), .B(G1341), .ZN(new_n1186));
  OAI22_X1  g761(.A1(new_n1082), .A2(G1996), .B1(new_n1106), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(new_n561), .ZN(new_n1188));
  XOR2_X1   g763(.A(new_n1188), .B(KEYINPUT59), .Z(new_n1189));
  AOI211_X1 g764(.A(new_n1180), .B(new_n621), .C1(new_n1163), .C2(new_n1169), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1172), .B1(new_n1185), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1055), .A2(new_n1081), .A3(new_n1088), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1085), .A2(new_n1086), .A3(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g769(.A(G301), .B(KEYINPUT54), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1085), .A2(new_n1086), .A3(new_n1089), .A4(new_n1195), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1123), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1199), .A2(new_n1074), .A3(new_n1200), .ZN(new_n1201));
  OAI211_X1 g776(.A(new_n1127), .B(new_n1142), .C1(new_n1192), .C2(new_n1201), .ZN(new_n1202));
  NOR3_X1   g777(.A1(new_n1041), .A2(KEYINPUT45), .A3(new_n1048), .ZN(new_n1203));
  AND2_X1   g778(.A1(new_n841), .A2(new_n844), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n841), .A2(new_n844), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1203), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n771), .B(new_n773), .ZN(new_n1207));
  INV_X1    g782(.A(G1996), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n704), .A2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1203), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT117), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1203), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1211), .B1(new_n1212), .B2(G1996), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1203), .A2(KEYINPUT117), .A3(new_n1208), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT118), .ZN(new_n1216));
  AND3_X1   g791(.A1(new_n1215), .A2(new_n1216), .A3(new_n705), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1216), .B1(new_n1215), .B2(new_n705), .ZN(new_n1218));
  OAI211_X1 g793(.A(new_n1206), .B(new_n1210), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1219));
  XNOR2_X1  g794(.A(G290), .B(G1986), .ZN(new_n1220));
  AOI21_X1  g795(.A(new_n1219), .B1(new_n1203), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1202), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT46), .ZN(new_n1223));
  XNOR2_X1  g798(.A(new_n1215), .B(new_n1223), .ZN(new_n1224));
  INV_X1    g799(.A(KEYINPUT47), .ZN(new_n1225));
  INV_X1    g800(.A(new_n704), .ZN(new_n1226));
  OAI21_X1  g801(.A(new_n1203), .B1(new_n1207), .B2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1224), .A2(new_n1225), .A3(new_n1227), .ZN(new_n1228));
  INV_X1    g803(.A(new_n1228), .ZN(new_n1229));
  AOI21_X1  g804(.A(new_n1225), .B1(new_n1224), .B2(new_n1227), .ZN(new_n1230));
  NOR3_X1   g805(.A1(G290), .A2(new_n1212), .A3(G1986), .ZN(new_n1231));
  XNOR2_X1  g806(.A(new_n1231), .B(KEYINPUT48), .ZN(new_n1232));
  OAI22_X1  g807(.A1(new_n1229), .A2(new_n1230), .B1(new_n1219), .B2(new_n1232), .ZN(new_n1233));
  OAI211_X1 g808(.A(new_n1205), .B(new_n1210), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n771), .A2(new_n773), .ZN(new_n1235));
  AOI21_X1  g810(.A(new_n1212), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NOR2_X1   g811(.A1(new_n1233), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1222), .A2(new_n1237), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g813(.A1(new_n950), .A2(new_n952), .ZN(new_n1240));
  INV_X1    g814(.A(G319), .ZN(new_n1241));
  NOR3_X1   g815(.A1(G401), .A2(new_n1241), .A3(G227), .ZN(new_n1242));
  AND3_X1   g816(.A1(new_n693), .A2(new_n694), .A3(new_n1242), .ZN(new_n1243));
  NAND3_X1  g817(.A1(new_n1240), .A2(new_n1243), .A3(new_n1025), .ZN(G225));
  INV_X1    g818(.A(G225), .ZN(G308));
endmodule


