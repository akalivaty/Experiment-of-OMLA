//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 1 0 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n547, new_n549, new_n550, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n593, new_n596, new_n597,
    new_n599, new_n600, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n465), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(G101), .A3(G2104), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT67), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n468), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT68), .ZN(G160));
  NAND2_X1  g050(.A1(new_n469), .A2(KEYINPUT69), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n477), .B1(new_n465), .B2(G2105), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n465), .A2(new_n471), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n461), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  AOI22_X1  g059(.A1(new_n481), .A2(G124), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND4_X1  g062(.A1(new_n462), .A2(new_n464), .A3(KEYINPUT4), .A4(G138), .ZN(new_n488));
  NAND2_X1  g063(.A1(G102), .A2(G2104), .ZN(new_n489));
  AOI21_X1  g064(.A(G2105), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  XNOR2_X1  g065(.A(KEYINPUT3), .B(G2104), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n491), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT4), .B1(new_n492), .B2(new_n471), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n491), .A2(G138), .A3(new_n471), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(G164));
  INV_X1    g070(.A(G50), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(G651), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(G651), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  OAI21_X1  g081(.A(G543), .B1(new_n506), .B2(KEYINPUT71), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT5), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n504), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n496), .A2(new_n505), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(G62), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n500), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n514), .A2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  INV_X1    g096(.A(G51), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n504), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n507), .A2(new_n510), .ZN(new_n524));
  OAI221_X1 g099(.A(new_n521), .B1(new_n505), .B2(new_n522), .C1(new_n523), .C2(new_n524), .ZN(G286));
  INV_X1    g100(.A(G286), .ZN(G168));
  AOI22_X1  g101(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n527), .A2(new_n500), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n502), .A2(new_n503), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n524), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G90), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n529), .A2(new_n509), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G52), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n528), .A2(new_n531), .A3(new_n533), .ZN(G171));
  NAND2_X1  g109(.A1(new_n530), .A2(G81), .ZN(new_n535));
  XOR2_X1   g110(.A(KEYINPUT72), .B(G43), .Z(new_n536));
  NAND2_X1  g111(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(G68), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G56), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n524), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n535), .A2(new_n537), .A3(new_n541), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(KEYINPUT73), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(KEYINPUT73), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(G188));
  NAND4_X1  g126(.A1(new_n502), .A2(G53), .A3(G543), .A4(new_n503), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT9), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n530), .A2(G91), .ZN(new_n554));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n524), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n553), .A2(new_n554), .A3(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  NAND2_X1  g135(.A1(new_n530), .A2(G87), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n532), .A2(G49), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(G288));
  NAND2_X1  g139(.A1(G73), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G61), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n524), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n532), .A2(G48), .B1(new_n567), .B2(G651), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n530), .A2(G86), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT74), .ZN(G305));
  INV_X1    g146(.A(G47), .ZN(new_n572));
  INV_X1    g147(.A(G85), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n572), .A2(new_n505), .B1(new_n512), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n574), .A2(new_n575), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  OAI22_X1  g153(.A1(new_n576), .A2(new_n577), .B1(new_n500), .B2(new_n578), .ZN(G290));
  XOR2_X1   g154(.A(KEYINPUT76), .B(KEYINPUT10), .Z(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(G92), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n512), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(new_n500), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n530), .A2(G92), .A3(new_n580), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n532), .A2(G54), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n583), .A2(new_n585), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n590), .B1(new_n589), .B2(G171), .ZN(G284));
  OAI21_X1  g166(.A(new_n590), .B1(new_n589), .B2(G171), .ZN(G321));
  NAND2_X1  g167(.A1(G299), .A2(new_n589), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(G168), .B2(new_n589), .ZN(G297));
  OAI21_X1  g169(.A(new_n593), .B1(G168), .B2(new_n589), .ZN(G280));
  INV_X1    g170(.A(new_n588), .ZN(new_n596));
  INV_X1    g171(.A(G559), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(G860), .ZN(G148));
  NOR2_X1   g173(.A1(new_n588), .A2(G559), .ZN(new_n599));
  MUX2_X1   g174(.A(new_n599), .B(new_n545), .S(new_n589), .Z(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT77), .ZN(G323));
  XNOR2_X1  g176(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g177(.A1(new_n479), .A2(G135), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n481), .A2(G123), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n471), .A2(G111), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT78), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n461), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI221_X1 g182(.A(new_n607), .B1(new_n606), .B2(new_n605), .C1(G99), .C2(G2105), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n603), .A2(new_n604), .A3(new_n608), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(G2096), .Z(new_n610));
  NAND3_X1  g185(.A1(new_n471), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2100), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n610), .A2(new_n614), .ZN(G156));
  XNOR2_X1  g190(.A(G2427), .B(G2438), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(G2430), .ZN(new_n617));
  XOR2_X1   g192(.A(KEYINPUT15), .B(G2435), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(KEYINPUT14), .ZN(new_n620));
  XNOR2_X1  g195(.A(G2451), .B(G2454), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT79), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT16), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n620), .B(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(G1341), .B(G1348), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2443), .B(G2446), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n626), .B(new_n627), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G14), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(G401));
  XOR2_X1   g205(.A(G2084), .B(G2090), .Z(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2067), .B(G2678), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT80), .Z(new_n634));
  XNOR2_X1  g209(.A(G2072), .B(G2078), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT81), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n632), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT82), .Z(new_n638));
  INV_X1    g213(.A(new_n634), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n636), .B(KEYINPUT17), .Z(new_n640));
  OAI21_X1  g215(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n634), .A2(new_n636), .A3(new_n631), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT18), .Z(new_n643));
  NAND3_X1  g218(.A1(new_n640), .A2(new_n639), .A3(new_n631), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n641), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2096), .B(G2100), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(G227));
  XNOR2_X1  g222(.A(G1971), .B(G1976), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT19), .ZN(new_n649));
  XOR2_X1   g224(.A(G1956), .B(G2474), .Z(new_n650));
  XOR2_X1   g225(.A(G1961), .B(G1966), .Z(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n649), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n650), .A2(new_n651), .ZN(new_n655));
  AOI22_X1  g230(.A1(new_n653), .A2(KEYINPUT20), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n657), .A2(new_n649), .A3(new_n652), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n656), .B(new_n658), .C1(KEYINPUT20), .C2(new_n653), .ZN(new_n659));
  XOR2_X1   g234(.A(G1991), .B(G1996), .Z(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT83), .B(G1986), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G1981), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n663), .B(new_n665), .ZN(G229));
  INV_X1    g241(.A(G19), .ZN(new_n667));
  OAI21_X1  g242(.A(KEYINPUT89), .B1(new_n667), .B2(G16), .ZN(new_n668));
  OR3_X1    g243(.A1(new_n667), .A2(KEYINPUT89), .A3(G16), .ZN(new_n669));
  INV_X1    g244(.A(G16), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n668), .B(new_n669), .C1(new_n545), .C2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT90), .B(G1341), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  AND2_X1   g248(.A1(KEYINPUT84), .A2(G29), .ZN(new_n674));
  NOR2_X1   g249(.A1(KEYINPUT84), .A2(G29), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(G26), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n479), .A2(G140), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT91), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(G104), .A2(G2105), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n684), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n481), .A2(G128), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT92), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n680), .B1(new_n689), .B2(G29), .ZN(new_n690));
  INV_X1    g265(.A(G2067), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n670), .A2(G4), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(new_n596), .B2(new_n670), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n694), .A2(G1348), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(G1348), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n677), .A2(G35), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G162), .B2(new_n677), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT29), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n696), .B1(new_n699), .B2(G2090), .ZN(new_n700));
  NOR3_X1   g275(.A1(new_n692), .A2(new_n695), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n670), .A2(G20), .ZN(new_n702));
  AND3_X1   g277(.A1(new_n553), .A2(new_n554), .A3(new_n558), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n670), .ZN(new_n704));
  MUX2_X1   g279(.A(new_n702), .B(new_n704), .S(KEYINPUT23), .Z(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT100), .B(G1956), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n699), .A2(G2090), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n709), .A2(KEYINPUT101), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(KEYINPUT101), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n701), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(G29), .A2(G32), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n479), .A2(G141), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT95), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n471), .A2(G105), .A3(G2104), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n481), .A2(G129), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT26), .ZN(new_n718));
  NAND3_X1  g293(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT96), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n717), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n718), .B2(new_n720), .ZN(new_n722));
  AND3_X1   g297(.A1(new_n715), .A2(new_n716), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n713), .B1(new_n723), .B2(G29), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT27), .B(G1996), .Z(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n670), .A2(G21), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G168), .B2(new_n670), .ZN(new_n728));
  INV_X1    g303(.A(G1966), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT98), .B(G28), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT30), .ZN(new_n732));
  OAI22_X1  g307(.A1(new_n609), .A2(new_n677), .B1(G29), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(G171), .A2(G16), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G5), .B2(G16), .ZN(new_n735));
  INV_X1    g310(.A(G1961), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n733), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n726), .A2(new_n730), .A3(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT31), .B(G11), .Z(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT24), .B(G34), .ZN(new_n740));
  AOI22_X1  g315(.A1(G160), .A2(G29), .B1(new_n677), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G2084), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n736), .B2(new_n735), .ZN(new_n743));
  NOR2_X1   g318(.A1(G164), .A2(new_n677), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G27), .B2(new_n677), .ZN(new_n745));
  INV_X1    g320(.A(G2078), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n747), .B(new_n748), .C1(G2084), .C2(new_n741), .ZN(new_n749));
  NOR4_X1   g324(.A1(new_n738), .A2(new_n739), .A3(new_n743), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n479), .A2(G139), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT25), .Z(new_n753));
  AOI22_X1  g328(.A1(new_n491), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT94), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n751), .B(new_n753), .C1(new_n471), .C2(new_n755), .ZN(new_n756));
  MUX2_X1   g331(.A(G33), .B(new_n756), .S(G29), .Z(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(G2072), .Z(new_n758));
  NOR2_X1   g333(.A1(new_n724), .A2(new_n725), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT97), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n750), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(KEYINPUT99), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(KEYINPUT99), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n712), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT86), .ZN(new_n765));
  NAND2_X1  g340(.A1(G288), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n562), .A2(new_n561), .A3(KEYINPUT86), .A4(new_n563), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(G16), .ZN(new_n769));
  INV_X1    g344(.A(G23), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(G16), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT33), .B(G1976), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n670), .A2(G22), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G166), .B2(new_n670), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n776), .A2(G1971), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n769), .B(new_n772), .C1(G16), .C2(new_n770), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(G1971), .ZN(new_n779));
  AND4_X1   g354(.A1(new_n774), .A2(new_n777), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n670), .A2(G6), .ZN(new_n781));
  INV_X1    g356(.A(G305), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(new_n670), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT32), .B(G1981), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n780), .A2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT34), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT87), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n676), .A2(G25), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n479), .A2(G131), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n481), .A2(G119), .ZN(new_n793));
  NOR2_X1   g368(.A1(G95), .A2(G2105), .ZN(new_n794));
  OAI21_X1  g369(.A(G2104), .B1(new_n471), .B2(G107), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n792), .B(new_n793), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT85), .Z(new_n797));
  AOI21_X1  g372(.A(new_n791), .B1(new_n797), .B2(new_n676), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT35), .B(G1991), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n798), .B(new_n800), .ZN(new_n801));
  MUX2_X1   g376(.A(G24), .B(G290), .S(G16), .Z(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(G1986), .Z(new_n803));
  NAND4_X1  g378(.A1(new_n789), .A2(new_n790), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n780), .A2(new_n785), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n801), .B(new_n803), .C1(new_n805), .C2(KEYINPUT34), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(KEYINPUT87), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n788), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n809), .ZN(new_n811));
  AOI211_X1 g386(.A(new_n788), .B(new_n811), .C1(new_n804), .C2(new_n807), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n673), .B(new_n764), .C1(new_n810), .C2(new_n812), .ZN(G150));
  INV_X1    g388(.A(G150), .ZN(G311));
  INV_X1    g389(.A(KEYINPUT104), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n504), .A2(G55), .A3(G543), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT102), .B(G93), .Z(new_n817));
  NAND3_X1  g392(.A1(new_n504), .A2(new_n511), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(KEYINPUT103), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n816), .A2(new_n818), .A3(KEYINPUT103), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(new_n500), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n815), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  AND3_X1   g400(.A1(new_n816), .A2(new_n818), .A3(KEYINPUT103), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n815), .B(new_n824), .C1(new_n826), .C2(new_n819), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n542), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n544), .A2(new_n543), .B1(new_n822), .B2(new_n824), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n588), .A2(new_n597), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n836), .A2(G860), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT105), .Z(new_n838));
  NOR2_X1   g413(.A1(new_n825), .A2(new_n828), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G860), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT106), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT37), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n838), .A2(new_n842), .ZN(G145));
  XNOR2_X1  g418(.A(G160), .B(new_n609), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n486), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT108), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n612), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n723), .ZN(new_n849));
  INV_X1    g424(.A(new_n689), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n479), .A2(G142), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n481), .A2(G130), .ZN(new_n852));
  NOR2_X1   g427(.A1(G106), .A2(G2105), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(new_n471), .B2(G118), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n851), .B(new_n852), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n850), .A2(new_n855), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n849), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n689), .B(new_n855), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(new_n723), .ZN(new_n860));
  XNOR2_X1  g435(.A(G164), .B(KEYINPUT107), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n858), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n862), .B1(new_n858), .B2(new_n860), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n756), .B(new_n796), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n858), .A2(new_n860), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n861), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n866), .B1(new_n870), .B2(new_n863), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n848), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(G37), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n867), .B1(new_n864), .B2(new_n865), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n870), .A2(new_n866), .A3(new_n863), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(new_n847), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n872), .A2(new_n873), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(KEYINPUT40), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n872), .A2(new_n879), .A3(new_n873), .A4(new_n876), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(G395));
  NAND2_X1  g456(.A1(new_n839), .A2(new_n589), .ZN(new_n882));
  INV_X1    g457(.A(new_n768), .ZN(new_n883));
  XNOR2_X1  g458(.A(G290), .B(G303), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n884), .A2(new_n782), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n782), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n884), .A2(new_n782), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n884), .A2(new_n782), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n768), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT42), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n832), .B(new_n599), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n703), .A2(new_n588), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n586), .A2(new_n587), .ZN(new_n895));
  NAND4_X1  g470(.A1(G299), .A2(new_n895), .A3(new_n585), .A4(new_n583), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT41), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT110), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n894), .A2(new_n896), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n703), .A2(KEYINPUT109), .A3(new_n588), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n900), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT110), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n897), .A2(new_n906), .A3(KEYINPUT41), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n901), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n899), .B1(new_n893), .B2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n892), .B(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n882), .B1(new_n910), .B2(new_n589), .ZN(G295));
  OAI21_X1  g486(.A(new_n882), .B1(new_n910), .B2(new_n589), .ZN(G331));
  NAND3_X1  g487(.A1(new_n829), .A2(new_n831), .A3(G301), .ZN(new_n913));
  INV_X1    g488(.A(new_n542), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n824), .B1(new_n826), .B2(new_n819), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT104), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n914), .B1(new_n916), .B2(new_n827), .ZN(new_n917));
  OAI21_X1  g492(.A(G171), .B1(new_n917), .B2(new_n830), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n913), .A2(new_n918), .A3(G168), .ZN(new_n919));
  AOI21_X1  g494(.A(G168), .B1(new_n913), .B2(new_n918), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n908), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(G301), .B1(new_n829), .B2(new_n831), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n917), .A2(new_n830), .A3(G171), .ZN(new_n923));
  OAI21_X1  g498(.A(G286), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n913), .A2(new_n918), .A3(G168), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n897), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n921), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(G37), .B1(new_n927), .B2(new_n891), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n887), .A2(new_n890), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n924), .A2(new_n925), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n897), .B1(new_n930), .B2(KEYINPUT41), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT111), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n933), .B1(new_n925), .B2(new_n924), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n929), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n928), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT112), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n929), .A2(new_n921), .A3(new_n926), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n928), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT112), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n928), .A2(new_n935), .A3(new_n942), .A4(new_n936), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n938), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n928), .A2(new_n935), .A3(KEYINPUT43), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT43), .B1(new_n928), .B2(new_n939), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT44), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n946), .A2(new_n949), .ZN(G397));
  NAND3_X1  g525(.A1(new_n462), .A2(new_n464), .A3(G126), .ZN(new_n951));
  NAND2_X1  g526(.A1(G114), .A2(G2104), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n471), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT4), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n494), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n490), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G1384), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  AND4_X1   g537(.A1(G40), .A2(new_n468), .A3(new_n470), .A4(new_n473), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n689), .B(new_n691), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n723), .B(G1996), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n797), .A2(new_n800), .ZN(new_n968));
  OAI22_X1  g543(.A1(new_n967), .A2(new_n968), .B1(G2067), .B2(new_n689), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT126), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n964), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n969), .A2(new_n970), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n964), .A2(G1996), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT46), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n965), .A2(new_n723), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n976), .B1(new_n977), .B2(new_n972), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n978), .B(KEYINPUT47), .Z(new_n979));
  XNOR2_X1  g554(.A(new_n796), .B(new_n799), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n967), .B1(new_n972), .B2(new_n980), .ZN(new_n981));
  OR2_X1    g556(.A1(G290), .A2(G1986), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(new_n964), .ZN(new_n983));
  XOR2_X1   g558(.A(new_n983), .B(KEYINPUT48), .Z(new_n984));
  NAND2_X1  g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n974), .A2(new_n979), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT125), .ZN(new_n987));
  INV_X1    g562(.A(G8), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n989));
  AOI21_X1  g564(.A(G1384), .B1(new_n955), .B2(new_n956), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n989), .A2(new_n963), .A3(new_n992), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n993), .A2(G2090), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n959), .A2(KEYINPUT113), .A3(new_n960), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(new_n990), .B2(KEYINPUT45), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n990), .A2(KEYINPUT45), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n995), .A2(new_n997), .A3(new_n963), .A4(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1971), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n988), .B1(new_n994), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT114), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n1005));
  NAND4_X1  g580(.A1(G303), .A2(new_n1005), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1006));
  NOR2_X1   g581(.A1(G166), .A2(new_n988), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1004), .B(new_n1006), .C1(new_n1007), .C2(KEYINPUT55), .ZN(new_n1008));
  OR2_X1    g583(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n990), .A2(new_n963), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(G8), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1976), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT52), .B1(G288), .B2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1013), .B(new_n1015), .C1(new_n768), .C2(new_n1014), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT49), .ZN(new_n1017));
  INV_X1    g592(.A(G1981), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n568), .A2(new_n1018), .A3(new_n569), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  XOR2_X1   g595(.A(KEYINPUT115), .B(G86), .Z(new_n1021));
  NAND2_X1  g596(.A1(new_n530), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1018), .B1(new_n568), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1017), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n568), .A2(new_n1022), .ZN(new_n1025));
  OAI211_X1 g600(.A(KEYINPUT49), .B(new_n1019), .C1(new_n1025), .C2(new_n1018), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1024), .A2(new_n1013), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1014), .B1(new_n766), .B2(new_n767), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT52), .B1(new_n1028), .B2(new_n1012), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1016), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1009), .A2(new_n1010), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1033), .B1(new_n999), .B2(G2078), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n993), .A2(new_n736), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1033), .A2(G2078), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n961), .A2(new_n963), .A3(new_n998), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(G171), .B(KEYINPUT54), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n963), .B1(new_n990), .B2(KEYINPUT45), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n1043), .A2(KEYINPUT124), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(KEYINPUT124), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1044), .A2(new_n998), .A3(new_n1045), .A4(new_n1037), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1036), .A2(new_n1040), .A3(new_n1046), .ZN(new_n1047));
  AOI211_X1 g622(.A(new_n960), .B(G1384), .C1(new_n955), .C2(new_n956), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n729), .B1(new_n1043), .B2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT119), .B(G2084), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n989), .A2(new_n992), .A3(new_n963), .A4(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1049), .A2(G168), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(G8), .ZN(new_n1053));
  AOI21_X1  g628(.A(G168), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n988), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT51), .B1(new_n1056), .B2(KEYINPUT123), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G8), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT123), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1053), .B1(new_n1062), .B2(KEYINPUT51), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1042), .B(new_n1047), .C1(new_n1058), .C2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G1956), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n993), .A2(new_n1065), .ZN(new_n1066));
  XOR2_X1   g641(.A(KEYINPUT56), .B(G2072), .Z(new_n1067));
  OAI21_X1  g642(.A(new_n1066), .B1(new_n999), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n1069));
  AND3_X1   g644(.A1(G299), .A2(new_n1069), .A3(KEYINPUT57), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT57), .B1(G299), .B2(new_n1069), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1068), .A2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1072), .B(new_n1066), .C1(new_n999), .C2(new_n1067), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1074), .A2(KEYINPUT61), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT61), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n990), .A2(new_n963), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT58), .B(G1341), .ZN(new_n1080));
  OAI22_X1  g655(.A1(new_n999), .A2(G1996), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n545), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1082), .B(KEYINPUT59), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1011), .A2(G2067), .ZN(new_n1084));
  INV_X1    g659(.A(G1348), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n993), .B2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1086), .A2(KEYINPUT122), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n1088));
  AOI211_X1 g663(.A(new_n1088), .B(new_n1084), .C1(new_n1085), .C2(new_n993), .ZN(new_n1089));
  OAI211_X1 g664(.A(KEYINPUT60), .B(new_n588), .C1(new_n1087), .C2(new_n1089), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1086), .A2(KEYINPUT122), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT60), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1086), .A2(KEYINPUT122), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT60), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1094), .A2(new_n1095), .A3(new_n596), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1078), .A2(new_n1083), .A3(new_n1090), .A4(new_n1096), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1075), .A2(new_n596), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1098), .A2(new_n1099), .B1(new_n1073), .B2(new_n1068), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1064), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT62), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1053), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n1057), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT62), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1104), .B(new_n1105), .C1(new_n1057), .C2(new_n1055), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1102), .A2(G171), .A3(new_n1039), .A4(new_n1106), .ZN(new_n1107));
  OR3_X1    g682(.A1(new_n1060), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1032), .B1(new_n1101), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1030), .A2(KEYINPUT116), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT116), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1016), .A2(new_n1027), .A3(new_n1029), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1114), .A2(new_n1010), .ZN(new_n1115));
  NOR2_X1   g690(.A1(G288), .A2(G1976), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1116), .B(KEYINPUT118), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1027), .A2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1019), .B(KEYINPUT117), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1012), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1121), .B1(new_n1114), .B2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1009), .A2(KEYINPUT120), .A3(new_n1111), .A4(new_n1113), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1060), .A2(G286), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .A4(new_n1010), .ZN(new_n1126));
  AOI211_X1 g701(.A(new_n1115), .B(new_n1120), .C1(new_n1126), .C2(KEYINPUT63), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1110), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(G290), .A2(G1986), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n982), .A2(new_n1129), .ZN(new_n1130));
  OR2_X1    g705(.A1(new_n1130), .A2(new_n964), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n981), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n987), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1134));
  AOI211_X1 g709(.A(KEYINPUT125), .B(new_n1132), .C1(new_n1110), .C2(new_n1127), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n986), .B1(new_n1134), .B2(new_n1135), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g711(.A(G229), .ZN(new_n1138));
  INV_X1    g712(.A(G319), .ZN(new_n1139));
  NOR2_X1   g713(.A1(G227), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g714(.A1(new_n629), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g715(.A(new_n1138), .B1(new_n1141), .B2(KEYINPUT127), .ZN(new_n1142));
  AOI21_X1  g716(.A(new_n1142), .B1(KEYINPUT127), .B2(new_n1141), .ZN(new_n1143));
  AND3_X1   g717(.A1(new_n944), .A2(new_n877), .A3(new_n1143), .ZN(G308));
  NAND3_X1  g718(.A1(new_n944), .A2(new_n877), .A3(new_n1143), .ZN(G225));
endmodule


