//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1285,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  INV_X1    g0003(.A(G107), .ZN(new_n204));
  INV_X1    g0004(.A(G264), .ZN(new_n205));
  INV_X1    g0005(.A(G116), .ZN(new_n206));
  INV_X1    g0006(.A(G270), .ZN(new_n207));
  OAI22_X1  g0007(.A1(new_n204), .A2(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(KEYINPUT65), .B(G244), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n208), .B(new_n213), .C1(G77), .C2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AND2_X1   g0020(.A1(G50), .A2(G226), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n203), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n203), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  AOI211_X1 g0025(.A(new_n212), .B(new_n225), .C1(new_n219), .C2(new_n205), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n226), .A2(KEYINPUT0), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n216), .A2(new_n209), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n230), .A2(G20), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n226), .A2(KEYINPUT0), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n227), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT64), .Z(new_n236));
  NOR2_X1   g0036(.A1(new_n223), .A2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G226), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G264), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n207), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  AND2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR3_X1   g0055(.A1(new_n254), .A2(new_n255), .A3(KEYINPUT67), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT67), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(G232), .B(G1698), .C1(new_n256), .C2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT70), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n259), .A2(new_n218), .ZN(new_n265));
  OAI21_X1  g0065(.A(KEYINPUT67), .B1(new_n254), .B2(new_n255), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n260), .A2(new_n257), .A3(new_n261), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1698), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n265), .B1(new_n268), .B2(G226), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(new_n267), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT70), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n270), .A2(new_n271), .A3(G232), .A4(G1698), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n264), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G1), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n276), .B1(G41), .B2(G45), .ZN(new_n277));
  INV_X1    g0077(.A(G274), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n274), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n277), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n280), .B1(new_n282), .B2(new_n210), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n275), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT13), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT13), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n275), .A2(new_n287), .A3(new_n284), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(G190), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n287), .B1(new_n275), .B2(new_n284), .ZN(new_n290));
  AOI211_X1 g0090(.A(KEYINPUT13), .B(new_n283), .C1(new_n273), .C2(new_n274), .ZN(new_n291));
  OAI21_X1  g0091(.A(G200), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n231), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT68), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n209), .A2(G20), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G20), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G50), .ZN(new_n300));
  INV_X1    g0100(.A(G20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G33), .ZN(new_n302));
  INV_X1    g0102(.A(G77), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n299), .A2(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n295), .B1(new_n297), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT11), .ZN(new_n306));
  INV_X1    g0106(.A(G13), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(G1), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT71), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT12), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(KEYINPUT71), .A2(KEYINPUT12), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n297), .A2(new_n308), .A3(new_n311), .A4(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n294), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n301), .A2(G1), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(G68), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n297), .A2(new_n308), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n318), .A2(new_n309), .A3(new_n310), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n306), .A2(new_n313), .A3(new_n317), .A4(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n289), .A2(new_n292), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n286), .A2(G179), .A3(new_n288), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT72), .ZN(new_n325));
  OAI21_X1  g0125(.A(G169), .B1(new_n290), .B2(new_n291), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT14), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT14), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n328), .B(G169), .C1(new_n290), .C2(new_n291), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT72), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n286), .A2(new_n330), .A3(G179), .A4(new_n288), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n325), .A2(new_n327), .A3(new_n329), .A4(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n323), .B1(new_n332), .B2(new_n320), .ZN(new_n333));
  INV_X1    g0133(.A(new_n282), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n279), .B1(new_n334), .B2(new_n214), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n270), .B1(new_n217), .B2(G1698), .ZN(new_n336));
  INV_X1    g0136(.A(G1698), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n210), .A2(new_n337), .ZN(new_n338));
  OAI22_X1  g0138(.A1(new_n336), .A2(new_n338), .B1(G107), .B2(new_n270), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n335), .B1(new_n339), .B2(new_n281), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n340), .A2(G179), .ZN(new_n341));
  INV_X1    g0141(.A(G169), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n341), .B1(new_n342), .B2(new_n340), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n294), .A2(new_n315), .A3(new_n303), .ZN(new_n344));
  XNOR2_X1  g0144(.A(KEYINPUT8), .B(G58), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n346), .A2(new_n298), .B1(G20), .B2(G77), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT15), .B(G87), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n347), .B1(new_n302), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n344), .B1(new_n349), .B2(new_n294), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n307), .A2(new_n301), .A3(G1), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n303), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n343), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n333), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(G20), .B1(new_n228), .B2(G50), .ZN(new_n356));
  INV_X1    g0156(.A(G150), .ZN(new_n357));
  OAI221_X1 g0157(.A(new_n356), .B1(new_n357), .B2(new_n299), .C1(new_n302), .C2(new_n345), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n295), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n359), .B(KEYINPUT69), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n295), .A2(new_n351), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(G50), .A3(new_n316), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n308), .A2(G20), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n362), .B1(G50), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n337), .A2(G222), .ZN(new_n366));
  NAND2_X1  g0166(.A1(G223), .A2(G1698), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n270), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n368), .B(new_n274), .C1(G77), .C2(new_n270), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n334), .A2(G226), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n369), .A2(new_n280), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n365), .A2(KEYINPUT9), .B1(new_n372), .B2(G190), .ZN(new_n373));
  OR2_X1    g0173(.A1(new_n360), .A2(new_n364), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT9), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n371), .A2(G200), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n373), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT10), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT10), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n373), .A2(new_n376), .A3(new_n380), .A4(new_n377), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n371), .A2(new_n342), .ZN(new_n383));
  INV_X1    g0183(.A(G179), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n372), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n374), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n346), .A2(new_n316), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n361), .A2(new_n389), .B1(new_n351), .B2(new_n345), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n216), .A2(new_n209), .ZN(new_n392));
  NOR2_X1   g0192(.A1(G58), .A2(G68), .ZN(new_n393));
  OAI21_X1  g0193(.A(G20), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n298), .A2(G159), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n260), .A2(new_n261), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  NOR3_X1   g0199(.A1(new_n398), .A2(new_n399), .A3(G20), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n266), .A2(new_n267), .A3(new_n301), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n400), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n397), .B1(new_n402), .B2(new_n209), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT16), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n399), .B1(new_n398), .B2(G20), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n254), .A2(new_n255), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(KEYINPUT7), .A3(new_n301), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n209), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n409), .A2(new_n396), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n314), .B1(new_n410), .B2(KEYINPUT16), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n391), .B1(new_n405), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n398), .B1(G226), .B2(new_n337), .ZN(new_n413));
  NOR2_X1   g0213(.A1(G223), .A2(G1698), .ZN(new_n414));
  OAI22_X1  g0214(.A1(new_n413), .A2(new_n414), .B1(new_n259), .B2(new_n211), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n279), .B1(new_n415), .B2(new_n274), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n334), .A2(G232), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G200), .ZN(new_n419));
  INV_X1    g0219(.A(new_n418), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G190), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n412), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT17), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n412), .A2(KEYINPUT17), .A3(new_n421), .A4(new_n419), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT18), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n418), .A2(G169), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n416), .A2(G179), .A3(new_n417), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n428), .B1(new_n431), .B2(new_n412), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n405), .A2(new_n411), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n390), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n430), .B1(new_n420), .B2(new_n342), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(KEYINPUT18), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n427), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n340), .A2(G200), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n350), .A2(new_n352), .ZN(new_n440));
  INV_X1    g0240(.A(G190), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n439), .B(new_n440), .C1(new_n441), .C2(new_n340), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  OR4_X1    g0243(.A1(new_n355), .A2(new_n387), .A3(new_n438), .A4(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n301), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT75), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n211), .A2(new_n218), .A3(new_n204), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n445), .A2(KEYINPUT75), .A3(new_n301), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n398), .A2(new_n301), .A3(G68), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n302), .A2(new_n218), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n451), .B(new_n452), .C1(KEYINPUT19), .C2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n294), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n348), .A2(new_n351), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT68), .ZN(new_n457));
  XNOR2_X1  g0257(.A(new_n294), .B(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n276), .A2(G33), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(new_n363), .A3(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n455), .B(new_n456), .C1(new_n211), .C2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT76), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n210), .A2(new_n337), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n398), .B(new_n463), .C1(G244), .C2(new_n337), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G116), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n281), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(G45), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n212), .B1(new_n467), .B2(G1), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n276), .A2(new_n278), .A3(G45), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n281), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n462), .B1(new_n471), .B2(G190), .ZN(new_n472));
  NOR4_X1   g0272(.A1(new_n466), .A2(new_n470), .A3(KEYINPUT76), .A4(new_n441), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n461), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n466), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n281), .A2(new_n468), .A3(new_n469), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G200), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n466), .A2(G179), .A3(new_n470), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n455), .A2(new_n456), .ZN(new_n480));
  INV_X1    g0280(.A(new_n460), .ZN(new_n481));
  INV_X1    g0281(.A(new_n348), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n479), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n477), .A2(new_n342), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n474), .A2(new_n478), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n398), .A2(G244), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT4), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n487), .A2(new_n488), .B1(G33), .B2(G283), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n270), .A2(KEYINPUT4), .A3(G244), .A4(new_n337), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n488), .B1(new_n270), .B2(G250), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n489), .B(new_n490), .C1(new_n491), .C2(new_n337), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n274), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT5), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT74), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT74), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT5), .ZN(new_n497));
  AOI21_X1  g0297(.A(G41), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(G41), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n276), .B(G45), .C1(new_n499), .C2(KEYINPUT5), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n281), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G257), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n498), .A2(new_n278), .A3(new_n274), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n500), .B(KEYINPUT73), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n493), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n342), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n460), .A2(new_n218), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n298), .A2(G77), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n204), .A2(KEYINPUT6), .A3(G97), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n218), .A2(new_n204), .ZN(new_n512));
  NOR2_X1   g0312(.A1(G97), .A2(G107), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n511), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G20), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n510), .B(new_n516), .C1(new_n402), .C2(new_n204), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n509), .B1(new_n517), .B2(new_n294), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n363), .A2(G97), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n493), .A2(new_n384), .A3(new_n503), .A4(new_n506), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n508), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n507), .A2(G200), .ZN(new_n524));
  AOI211_X1 g0324(.A(new_n519), .B(new_n509), .C1(new_n517), .C2(new_n294), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n493), .A2(G190), .A3(new_n503), .A4(new_n506), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n486), .A2(new_n523), .A3(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT77), .ZN(new_n529));
  XNOR2_X1  g0329(.A(new_n528), .B(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G283), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n531), .B(new_n301), .C1(G33), .C2(new_n218), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n532), .B(new_n294), .C1(new_n301), .C2(G116), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT20), .ZN(new_n534));
  OR2_X1    g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n351), .A2(new_n294), .A3(new_n206), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n537), .A2(KEYINPUT78), .A3(new_n459), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n314), .A2(new_n363), .A3(G116), .A4(new_n459), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT78), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n535), .A2(new_n536), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n351), .A2(new_n206), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n342), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n219), .A2(new_n337), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n398), .B(new_n545), .C1(G264), .C2(new_n337), .ZN(new_n546));
  INV_X1    g0346(.A(G303), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(new_n270), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n274), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n502), .A2(G270), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(new_n506), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n544), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT21), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n542), .A2(new_n543), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n551), .A2(G200), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n556), .B(new_n557), .C1(new_n441), .C2(new_n551), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n549), .A2(new_n506), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n555), .A2(G179), .A3(new_n550), .A4(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n544), .A2(KEYINPUT21), .A3(new_n551), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n554), .A2(new_n558), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT79), .ZN(new_n563));
  AND4_X1   g0363(.A1(KEYINPUT21), .A2(new_n555), .A3(G169), .A4(new_n551), .ZN(new_n564));
  AOI21_X1  g0364(.A(KEYINPUT21), .B1(new_n544), .B2(new_n551), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT79), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n566), .A2(new_n567), .A3(new_n560), .A4(new_n558), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n481), .A2(G107), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n308), .A2(G20), .A3(new_n204), .ZN(new_n571));
  XOR2_X1   g0371(.A(new_n571), .B(KEYINPUT25), .Z(new_n572));
  AND2_X1   g0372(.A1(KEYINPUT82), .A2(KEYINPUT24), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT23), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n301), .B2(G107), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n204), .A2(KEYINPUT23), .A3(G20), .ZN(new_n576));
  INV_X1    g0376(.A(new_n465), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n575), .A2(new_n576), .B1(new_n577), .B2(new_n301), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n211), .A2(G20), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n254), .B2(new_n255), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT80), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n579), .B(KEYINPUT80), .C1(new_n255), .C2(new_n254), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(KEYINPUT22), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT81), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT22), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n586), .B(new_n579), .C1(new_n256), .C2(new_n262), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n585), .B1(new_n584), .B2(new_n587), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n578), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(KEYINPUT82), .A2(KEYINPUT24), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI221_X1 g0392(.A(new_n578), .B1(KEYINPUT82), .B2(KEYINPUT24), .C1(new_n588), .C2(new_n589), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n573), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n570), .B(new_n572), .C1(new_n594), .C2(new_n314), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n398), .B1(G257), .B2(new_n337), .ZN(new_n597));
  NOR2_X1   g0397(.A1(G250), .A2(G1698), .ZN(new_n598));
  XNOR2_X1  g0398(.A(KEYINPUT83), .B(G294), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n597), .A2(new_n598), .B1(new_n259), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n274), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n502), .A2(G264), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n603), .A3(new_n506), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT84), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n602), .A2(new_n603), .A3(KEYINPUT84), .A4(new_n506), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(KEYINPUT86), .B1(new_n608), .B2(G190), .ZN(new_n609));
  INV_X1    g0409(.A(G200), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT86), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n606), .A2(new_n612), .A3(new_n441), .A4(new_n607), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n609), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n596), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT85), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n608), .A2(G169), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n384), .B2(new_n604), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n595), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n616), .B1(new_n595), .B2(new_n618), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n569), .B(new_n615), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n444), .A2(new_n530), .A3(new_n621), .ZN(G372));
  INV_X1    g0422(.A(new_n386), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT89), .ZN(new_n624));
  INV_X1    g0424(.A(new_n354), .ZN(new_n625));
  AOI211_X1 g0425(.A(new_n625), .B(new_n323), .C1(new_n332), .C2(new_n320), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n624), .B1(new_n626), .B2(new_n323), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n332), .A2(new_n320), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n323), .B1(new_n628), .B2(new_n354), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT89), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n627), .A2(new_n427), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n437), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n623), .B1(new_n632), .B2(new_n382), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n476), .A2(KEYINPUT87), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n476), .A2(KEYINPUT87), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n475), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n342), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n484), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT88), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n523), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n508), .A2(new_n521), .A3(KEYINPUT88), .A4(new_n522), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n523), .A2(new_n527), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n609), .A2(new_n611), .A3(new_n613), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n645), .B1(new_n646), .B2(new_n595), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n554), .A2(new_n560), .A3(new_n561), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n648), .B1(new_n595), .B2(new_n618), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n644), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n636), .A2(G200), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n474), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n639), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n486), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT26), .B1(new_n654), .B2(new_n523), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n633), .B1(new_n444), .B2(new_n656), .ZN(G369));
  NOR2_X1   g0457(.A1(new_n646), .A2(new_n595), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n595), .A2(new_n618), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(KEYINPUT85), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n595), .A2(new_n616), .A3(new_n618), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n308), .A2(new_n301), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT90), .ZN(new_n664));
  OR3_X1    g0464(.A1(new_n663), .A2(new_n664), .A3(KEYINPUT27), .ZN(new_n665));
  INV_X1    g0465(.A(G213), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n666), .B1(new_n663), .B2(KEYINPUT27), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n664), .B1(new_n663), .B2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n662), .B1(new_n596), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n659), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n671), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n556), .A2(new_n672), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n563), .B2(new_n568), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n648), .B2(new_n677), .ZN(new_n679));
  INV_X1    g0479(.A(G330), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n648), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(new_n671), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n662), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n674), .A2(new_n672), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n682), .A2(new_n688), .ZN(G399));
  NOR2_X1   g0489(.A1(new_n225), .A2(G41), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n449), .A2(G116), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G1), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n229), .B2(new_n691), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT28), .Z(new_n695));
  AOI211_X1 g0495(.A(KEYINPUT29), .B(new_n671), .C1(new_n653), .C2(new_n655), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n641), .A2(new_n652), .A3(new_n643), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT26), .ZN(new_n698));
  INV_X1    g0498(.A(new_n523), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(new_n642), .A3(new_n486), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n698), .A2(new_n638), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n647), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n648), .B1(new_n660), .B2(new_n661), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT93), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n652), .A2(new_n638), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n683), .B1(new_n619), .B2(new_n620), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n708), .B1(new_n709), .B2(KEYINPUT93), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n702), .B1(new_n706), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n672), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n696), .B1(new_n712), .B2(KEYINPUT29), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n528), .B(KEYINPUT77), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n662), .A2(new_n714), .A3(new_n569), .A4(new_n672), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  INV_X1    g0516(.A(new_n506), .ZN(new_n717));
  AOI221_X4 g0517(.A(new_n717), .B1(G257), .B2(new_n502), .C1(new_n492), .C2(new_n274), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n551), .A2(new_n477), .A3(new_n384), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n602), .A2(new_n603), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n718), .A2(new_n719), .A3(KEYINPUT30), .A4(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n493), .A2(new_n720), .A3(new_n503), .A4(new_n506), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n559), .A2(G179), .A3(new_n471), .A4(new_n550), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n551), .A2(new_n636), .A3(new_n384), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(new_n507), .A3(new_n604), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT91), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n722), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n726), .A2(new_n728), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(KEYINPUT91), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n716), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n726), .A2(new_n721), .A3(new_n728), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT92), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT92), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n726), .A2(new_n721), .A3(new_n728), .A4(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n736), .A2(new_n671), .A3(new_n738), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n734), .A2(new_n671), .B1(new_n716), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n715), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G330), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n713), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n695), .B1(new_n744), .B2(new_n276), .ZN(new_n745));
  XOR2_X1   g0545(.A(new_n745), .B(KEYINPUT94), .Z(G364));
  NOR2_X1   g0546(.A1(new_n307), .A2(G20), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G45), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n691), .A2(G1), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n749), .B1(new_n679), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n301), .A2(G190), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G179), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G159), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n755), .A2(G190), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n758), .A2(KEYINPUT32), .B1(new_n218), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n270), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(KEYINPUT32), .B2(new_n758), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n301), .A2(new_n441), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n384), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n754), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n767), .A2(new_n216), .B1(new_n768), .B2(new_n303), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT97), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n610), .A2(G179), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n765), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G87), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n769), .A2(new_n770), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n764), .A2(new_n771), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n384), .A2(new_n610), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n778), .A2(new_n754), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n762), .B(new_n777), .C1(G68), .C2(new_n779), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n765), .A2(new_n778), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n754), .A2(new_n772), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n780), .B1(new_n300), .B2(new_n782), .C1(new_n204), .C2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n768), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n785), .A2(G311), .B1(new_n760), .B2(new_n599), .ZN(new_n786));
  INV_X1    g0586(.A(G326), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(new_n787), .B2(new_n782), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT98), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n270), .B(new_n789), .C1(G303), .C2(new_n774), .ZN(new_n790));
  INV_X1    g0590(.A(new_n779), .ZN(new_n791));
  INV_X1    g0591(.A(G317), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n791), .B1(KEYINPUT33), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(KEYINPUT33), .B2(new_n792), .ZN(new_n794));
  INV_X1    g0594(.A(new_n783), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G283), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n757), .A2(KEYINPUT99), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n757), .A2(KEYINPUT99), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G329), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n790), .A2(new_n794), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n767), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n802), .A2(G322), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n784), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n231), .B1(G20), .B2(new_n342), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n225), .A2(new_n398), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(new_n467), .B2(new_n230), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n249), .B2(new_n467), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n270), .A2(G355), .A3(new_n224), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n810), .B(new_n811), .C1(G116), .C2(new_n224), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n752), .A2(new_n805), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n753), .A2(new_n806), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n679), .A2(KEYINPUT95), .A3(new_n680), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n749), .ZN(new_n817));
  AOI21_X1  g0617(.A(KEYINPUT95), .B1(new_n679), .B2(new_n680), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n681), .A2(KEYINPUT96), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT96), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n679), .B2(new_n680), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n815), .B1(new_n819), .B2(new_n824), .ZN(G396));
  NAND2_X1  g0625(.A1(new_n650), .A2(new_n652), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n826), .A2(new_n655), .A3(new_n638), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n625), .A2(new_n672), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n442), .B1(new_n440), .B2(new_n672), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n354), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n827), .A2(new_n672), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n671), .B1(new_n653), .B2(new_n655), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n831), .A2(KEYINPUT103), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT103), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n828), .A2(new_n836), .A3(new_n830), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n833), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT104), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(G330), .A3(new_n741), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n742), .B1(new_n840), .B2(new_n841), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n843), .B(new_n749), .C1(new_n844), .C2(new_n842), .ZN(new_n845));
  AOI22_X1  g0645(.A1(G143), .A2(new_n802), .B1(new_n785), .B2(G159), .ZN(new_n846));
  INV_X1    g0646(.A(G137), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n846), .B1(new_n847), .B2(new_n782), .C1(new_n357), .C2(new_n791), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT34), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n783), .A2(new_n209), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n407), .B(new_n850), .C1(G50), .C2(new_n774), .ZN(new_n851));
  INV_X1    g0651(.A(G132), .ZN(new_n852));
  INV_X1    g0652(.A(new_n799), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n849), .B(new_n851), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n761), .A2(new_n216), .ZN(new_n855));
  INV_X1    g0655(.A(G294), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n761), .A2(new_n218), .B1(new_n767), .B2(new_n856), .ZN(new_n857));
  XNOR2_X1  g0657(.A(KEYINPUT101), .B(G283), .ZN(new_n858));
  AOI22_X1  g0658(.A1(G303), .A2(new_n781), .B1(new_n779), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n211), .B2(new_n783), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n857), .B(new_n860), .C1(G311), .C2(new_n799), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n206), .B2(new_n768), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n763), .B1(new_n204), .B2(new_n773), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT102), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n854), .A2(new_n855), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n805), .ZN(new_n866));
  INV_X1    g0666(.A(new_n749), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n805), .A2(new_n750), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n867), .B1(G77), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT100), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n866), .B(new_n871), .C1(new_n832), .C2(new_n751), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n845), .A2(new_n872), .ZN(G384));
  NOR2_X1   g0673(.A1(new_n321), .A2(new_n672), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n333), .A2(KEYINPUT105), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n875), .B1(new_n333), .B2(KEYINPUT105), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n833), .B2(new_n828), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT106), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n828), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n834), .B2(new_n832), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT106), .B1(new_n883), .B2(new_n878), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n410), .A2(KEYINPUT16), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n404), .B1(new_n409), .B2(new_n396), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(new_n295), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n390), .ZN(new_n888));
  INV_X1    g0688(.A(new_n669), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n432), .A2(new_n436), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n891), .B1(new_n892), .B2(new_n426), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n435), .A2(new_n888), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n422), .A2(new_n894), .A3(new_n890), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT37), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n434), .B1(new_n435), .B2(new_n889), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT37), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n897), .A2(new_n898), .A3(new_n422), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n896), .A2(new_n899), .A3(KEYINPUT107), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT107), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n895), .A2(new_n901), .A3(KEYINPUT37), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n893), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT38), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n893), .A2(new_n900), .A3(KEYINPUT38), .A4(new_n902), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n881), .A2(new_n884), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n892), .A2(new_n669), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n628), .A2(new_n671), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n434), .A2(new_n889), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n427), .B2(new_n437), .ZN(new_n912));
  INV_X1    g0712(.A(new_n899), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n898), .B1(new_n897), .B2(new_n422), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n904), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT39), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n916), .A2(new_n917), .A3(new_n906), .ZN(new_n918));
  AOI22_X1  g0718(.A1(KEYINPUT39), .A2(new_n907), .B1(new_n918), .B2(KEYINPUT108), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n907), .A2(KEYINPUT108), .A3(KEYINPUT39), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n910), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n908), .A2(new_n909), .A3(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT111), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n707), .B1(new_n704), .B2(new_n705), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n647), .B1(new_n709), .B2(KEYINPUT93), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n701), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT29), .B1(new_n926), .B2(new_n671), .ZN(new_n927));
  INV_X1    g0727(.A(new_n696), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n444), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n629), .A2(KEYINPUT89), .ZN(new_n930));
  AOI211_X1 g0730(.A(new_n624), .B(new_n323), .C1(new_n628), .C2(new_n354), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n930), .A2(new_n931), .A3(new_n426), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n382), .B1(new_n932), .B2(new_n892), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n386), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n923), .B(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n907), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n628), .A2(KEYINPUT105), .A3(new_n322), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n874), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n333), .A2(KEYINPUT105), .A3(new_n875), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n831), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n716), .A2(KEYINPUT109), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n739), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n715), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT110), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n937), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n941), .B(new_n944), .C1(KEYINPUT110), .C2(KEYINPUT40), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n916), .A2(new_n906), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n941), .A2(new_n944), .A3(new_n949), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n947), .A2(new_n948), .B1(KEYINPUT40), .B2(new_n950), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n621), .A2(new_n530), .A3(new_n671), .ZN(new_n952));
  INV_X1    g0752(.A(new_n942), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n739), .B(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n955), .A2(new_n444), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n951), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(G330), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n936), .B(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n276), .B2(new_n747), .ZN(new_n960));
  OAI211_X1 g0760(.A(G20), .B(new_n232), .C1(new_n515), .C2(KEYINPUT35), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n206), .B(new_n961), .C1(KEYINPUT35), .C2(new_n515), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT36), .Z(new_n963));
  OAI21_X1  g0763(.A(G77), .B1(new_n216), .B2(new_n209), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n229), .A2(new_n964), .B1(G50), .B2(new_n209), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n965), .A2(G1), .A3(new_n307), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n960), .A2(new_n963), .A3(new_n966), .ZN(G367));
  INV_X1    g0767(.A(new_n682), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n645), .B1(new_n525), .B2(new_n672), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n699), .A2(new_n671), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT114), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n645), .ZN(new_n975));
  OAI21_X1  g0775(.A(KEYINPUT42), .B1(new_n685), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n660), .A2(new_n661), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n523), .B1(new_n977), .B2(new_n969), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n672), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(KEYINPUT112), .ZN(new_n981));
  OR3_X1    g0781(.A1(new_n685), .A2(KEYINPUT42), .A3(new_n975), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT112), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n976), .A2(new_n983), .A3(new_n979), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n981), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n461), .A2(new_n671), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n708), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n638), .B2(new_n986), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT43), .ZN(new_n990));
  AND3_X1   g0790(.A1(new_n985), .A2(KEYINPUT113), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n990), .B1(new_n985), .B2(KEYINPUT113), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n985), .A2(KEYINPUT113), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n985), .A2(KEYINPUT113), .A3(new_n990), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n995), .A2(new_n996), .A3(new_n988), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n993), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n972), .A2(new_n973), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n974), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT115), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n1001), .B(KEYINPUT44), .C1(new_n688), .C2(new_n971), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n685), .A2(new_n686), .A3(new_n971), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(KEYINPUT45), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1003), .A2(KEYINPUT45), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(KEYINPUT115), .B(KEYINPUT44), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n687), .A2(new_n969), .A3(new_n970), .A4(new_n1006), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .A4(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n968), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1003), .B(KEYINPUT45), .Z(new_n1010));
  NAND4_X1  g0810(.A1(new_n1010), .A2(new_n682), .A3(new_n1002), .A4(new_n1007), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n676), .A2(new_n684), .ZN(new_n1013));
  AND3_X1   g0813(.A1(new_n1013), .A2(new_n681), .A3(new_n685), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n1013), .A2(new_n685), .B1(new_n822), .B2(new_n820), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n743), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n690), .B(KEYINPUT41), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n748), .A2(G1), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n993), .A2(new_n997), .A3(new_n973), .A4(new_n972), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1000), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n783), .A2(new_n218), .B1(new_n756), .B2(new_n792), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n407), .B1(new_n767), .B2(new_n547), .C1(new_n761), .C2(new_n204), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(new_n785), .C2(new_n858), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n774), .A2(G116), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT46), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1027), .B(new_n1029), .C1(new_n600), .C2(new_n791), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G311), .B2(new_n781), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n785), .A2(G50), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n774), .A2(G58), .B1(new_n781), .B2(G143), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n847), .B2(new_n756), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G68), .B2(new_n760), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n795), .A2(G77), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n763), .B1(G159), .B2(new_n779), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(G150), .B2(new_n802), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1031), .B1(new_n1032), .B2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT47), .Z(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n805), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n987), .B(new_n752), .C1(new_n638), .C2(new_n986), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n813), .B1(new_n224), .B2(new_n348), .C1(new_n245), .C2(new_n808), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1042), .A2(new_n867), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1024), .A2(new_n1045), .ZN(G387));
  NOR2_X1   g0846(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n743), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n690), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT117), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n744), .A2(new_n1016), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1048), .A2(KEYINPUT117), .A3(new_n690), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n802), .A2(G50), .B1(new_n482), .B2(new_n760), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n303), .B2(new_n773), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n209), .A2(new_n768), .B1(new_n783), .B2(new_n218), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n346), .B2(new_n779), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n757), .A2(G150), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n407), .B1(new_n781), .B2(G159), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1057), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G322), .A2(new_n781), .B1(new_n779), .B2(G311), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1063), .B1(new_n547), .B2(new_n768), .C1(new_n792), .C2(new_n767), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT48), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n858), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1065), .B1(new_n600), .B2(new_n773), .C1(new_n761), .C2(new_n1066), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT49), .Z(new_n1068));
  OAI221_X1 g0868(.A(new_n407), .B1(new_n756), .B2(new_n787), .C1(new_n206), .C2(new_n783), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1062), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT116), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n805), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n673), .A2(new_n675), .A3(new_n752), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n807), .B1(new_n242), .B2(new_n467), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n692), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n270), .A2(new_n1075), .A3(new_n224), .ZN(new_n1076));
  AOI211_X1 g0876(.A(G45), .B(new_n1075), .C1(G68), .C2(G77), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n345), .A2(G50), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT50), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1074), .A2(new_n1076), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n224), .A2(G107), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n813), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AND4_X1   g0882(.A1(new_n867), .A2(new_n1072), .A3(new_n1073), .A4(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n1047), .B2(new_n1020), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1054), .A2(new_n1084), .ZN(G393));
  NAND3_X1  g0885(.A1(new_n1009), .A2(new_n1011), .A3(new_n1020), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n969), .A2(new_n752), .A3(new_n970), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n802), .A2(G311), .B1(new_n781), .B2(G317), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT52), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n757), .A2(G322), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n763), .B1(new_n856), .B2(new_n768), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n791), .A2(new_n547), .B1(new_n783), .B2(new_n204), .ZN(new_n1092));
  NOR4_X1   g0892(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1093), .B1(new_n206), .B2(new_n761), .C1(new_n773), .C2(new_n1066), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n407), .B1(new_n757), .B2(G143), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1095), .B1(new_n209), .B2(new_n773), .C1(new_n211), .C2(new_n783), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT118), .Z(new_n1097));
  INV_X1    g0897(.A(G159), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n782), .A2(new_n357), .B1(new_n767), .B2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT51), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n779), .A2(G50), .B1(new_n760), .B2(G77), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n345), .B2(new_n768), .ZN(new_n1103));
  XOR2_X1   g0903(.A(new_n1103), .B(KEYINPUT119), .Z(new_n1104));
  OAI21_X1  g0904(.A(new_n1094), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n805), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n813), .B1(new_n218), .B2(new_n224), .C1(new_n252), .C2(new_n808), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1087), .A2(new_n867), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1086), .A2(new_n1108), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1048), .A2(new_n1012), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n691), .B1(new_n1048), .B2(new_n1012), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(G390));
  NAND2_X1  g0913(.A1(new_n939), .A2(new_n940), .ZN(new_n1114));
  AND4_X1   g0914(.A1(G330), .A2(new_n741), .A3(new_n832), .A4(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n680), .B1(new_n715), .B2(new_n943), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1114), .B1(new_n1116), .B2(new_n839), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n926), .A2(new_n671), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n882), .B1(new_n1119), .B2(new_n830), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n833), .A2(new_n828), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1116), .A2(new_n941), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n680), .B(new_n831), .C1(new_n715), .C2(new_n740), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1122), .B1(new_n1123), .B2(new_n1114), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1118), .A2(new_n1120), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n956), .A2(G330), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n633), .B(new_n1126), .C1(new_n713), .C2(new_n444), .ZN(new_n1127));
  OAI21_X1  g0927(.A(KEYINPUT120), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n741), .A2(G330), .A3(new_n832), .A4(new_n1114), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n680), .B(new_n838), .C1(new_n715), .C2(new_n943), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1129), .B1(new_n1130), .B2(new_n1114), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n711), .A2(new_n672), .A3(new_n830), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n828), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n734), .A2(new_n671), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n739), .A2(new_n716), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g0936(.A(G330), .B(new_n832), .C1(new_n952), .C2(new_n1136), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1137), .A2(new_n878), .B1(new_n1116), .B2(new_n941), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n1131), .A2(new_n1133), .B1(new_n1138), .B2(new_n883), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT120), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n935), .A2(new_n1139), .A3(new_n1140), .A4(new_n1126), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1128), .A2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n919), .A2(new_n920), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n879), .B2(new_n910), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n878), .B1(new_n1132), .B2(new_n828), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n910), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n949), .A2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1144), .B(new_n1115), .C1(new_n1145), .C2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1133), .A2(new_n1114), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1147), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1146), .B1(new_n883), .B2(new_n878), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1149), .A2(new_n1150), .B1(new_n1151), .B2(new_n1143), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1122), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1148), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n691), .B1(new_n1142), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1144), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n1122), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1128), .A2(new_n1157), .A3(new_n1141), .A4(new_n1148), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1021), .B1(new_n1157), .B2(new_n1148), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1143), .A2(new_n750), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n775), .B1(new_n206), .B2(new_n767), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n850), .B(new_n1162), .C1(G77), .C2(new_n760), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n785), .A2(G97), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n799), .A2(G294), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n270), .B1(G283), .B2(new_n781), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n791), .A2(new_n204), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT54), .B(G143), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n768), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n799), .A2(G125), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n791), .A2(new_n847), .B1(new_n852), .B2(new_n767), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT53), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n773), .B2(new_n357), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n774), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1172), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n760), .A2(G159), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n270), .B1(new_n300), .B2(new_n783), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G128), .B2(new_n781), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1171), .A2(new_n1176), .A3(new_n1177), .A4(new_n1179), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n1167), .A2(new_n1168), .B1(new_n1170), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n805), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1161), .A2(new_n867), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n345), .B2(new_n868), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1160), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1159), .A2(new_n1185), .ZN(G378));
  XOR2_X1   g0986(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n387), .B(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n374), .A2(new_n889), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1189), .B(new_n1190), .Z(new_n1191));
  AOI21_X1  g0991(.A(new_n749), .B1(new_n1191), .B2(new_n750), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n767), .A2(new_n204), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT122), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n209), .B2(new_n761), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n799), .A2(G283), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G77), .A2(new_n774), .B1(new_n795), .B2(G58), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1196), .A2(new_n499), .A3(new_n407), .A4(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT121), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1195), .B(new_n1199), .C1(new_n482), .C2(new_n785), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n218), .B2(new_n791), .C1(new_n206), .C2(new_n782), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT58), .Z(new_n1202));
  OAI21_X1  g1002(.A(new_n300), .B1(new_n254), .B2(G41), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n768), .A2(new_n847), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n761), .A2(new_n357), .B1(new_n773), .B2(new_n1169), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(G128), .C2(new_n802), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n781), .A2(G125), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n852), .C2(new_n791), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT59), .ZN(new_n1209));
  AOI211_X1 g1009(.A(G33), .B(G41), .C1(new_n757), .C2(G124), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n1098), .B2(new_n783), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1203), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n805), .B1(new_n1202), .B2(new_n1212), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1192), .B(new_n1213), .C1(G50), .C2(new_n869), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT123), .Z(new_n1215));
  XNOR2_X1  g1015(.A(new_n1189), .B(new_n1190), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n951), .B2(new_n680), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n832), .B1(new_n876), .B2(new_n877), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n946), .B1(new_n955), .B2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1219), .A2(new_n948), .A3(new_n907), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n950), .A2(KEYINPUT40), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1222), .A2(G330), .A3(new_n1191), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1217), .A2(KEYINPUT124), .A3(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n922), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n922), .A2(KEYINPUT124), .A3(new_n1217), .A4(new_n1223), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1215), .B1(new_n1228), .B2(new_n1020), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1125), .A2(new_n1127), .A3(KEYINPUT120), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n955), .A2(new_n444), .A3(new_n680), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n929), .A2(new_n934), .A3(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1140), .B1(new_n1232), .B2(new_n1139), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1154), .B1(new_n1230), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1232), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT57), .B1(new_n1235), .B2(new_n1228), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1127), .B1(new_n1142), .B2(new_n1154), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n921), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n880), .B1(new_n1121), .B2(new_n1114), .ZN(new_n1239));
  AOI211_X1 g1039(.A(KEYINPUT106), .B(new_n878), .C1(new_n833), .C2(new_n828), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1238), .B1(new_n1241), .B2(new_n907), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1242), .A2(new_n909), .A3(new_n1217), .A4(new_n1223), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1191), .B1(new_n1222), .B2(G330), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n680), .B(new_n1216), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n922), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1243), .A2(KEYINPUT57), .A3(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n690), .B1(new_n1237), .B2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1229), .B1(new_n1236), .B2(new_n1248), .ZN(G375));
  NAND2_X1  g1049(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1128), .A2(new_n1141), .A3(new_n1018), .A4(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n878), .A2(new_n750), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n868), .A2(new_n209), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n781), .A2(G132), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n1254), .B1(new_n847), .B2(new_n767), .C1(new_n791), .C2(new_n1169), .ZN(new_n1255));
  XOR2_X1   g1055(.A(new_n1255), .B(KEYINPUT126), .Z(new_n1256));
  NOR2_X1   g1056(.A1(new_n1256), .A2(new_n407), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n774), .A2(G159), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(G58), .A2(new_n795), .B1(new_n785), .B2(G150), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n799), .A2(G128), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .A4(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n761), .A2(new_n300), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n802), .A2(G283), .B1(new_n482), .B2(new_n760), .ZN(new_n1263));
  XOR2_X1   g1063(.A(new_n1263), .B(KEYINPUT125), .Z(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(G294), .B2(new_n781), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(G97), .A2(new_n774), .B1(new_n785), .B2(G107), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n779), .A2(G116), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1265), .A2(new_n1036), .A3(new_n1266), .A4(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n763), .B1(new_n853), .B2(new_n547), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n1261), .A2(new_n1262), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n805), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1252), .A2(new_n867), .A3(new_n1253), .A4(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1125), .B2(new_n1021), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1251), .A2(new_n1274), .ZN(G381));
  INV_X1    g1075(.A(G375), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n1160), .B(new_n1184), .C1(new_n1155), .C2(new_n1158), .ZN(new_n1277));
  INV_X1    g1077(.A(G396), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1054), .A2(new_n1278), .A3(new_n1084), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1024), .A2(new_n1045), .A3(new_n1112), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1276), .A2(new_n1277), .A3(new_n1279), .A4(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(G381), .A2(G384), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  OR2_X1    g1083(.A1(new_n1281), .A2(new_n1283), .ZN(G407));
  NAND3_X1  g1084(.A1(new_n1276), .A2(new_n670), .A3(new_n1277), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(G407), .A2(G213), .A3(new_n1285), .ZN(G409));
  OAI211_X1 g1086(.A(G378), .B(new_n1229), .C1(new_n1236), .C2(new_n1248), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1128), .A2(new_n1141), .B1(new_n1157), .B2(new_n1148), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1228), .B(new_n1018), .C1(new_n1127), .C2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1243), .A2(new_n1020), .A3(new_n1246), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1214), .B(KEYINPUT123), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1289), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1277), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1287), .A2(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n666), .A2(G343), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT60), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1128), .A2(new_n1141), .A3(new_n1250), .ZN(new_n1299));
  AOI211_X1 g1099(.A(new_n691), .B(new_n1298), .C1(new_n1299), .C2(KEYINPUT60), .ZN(new_n1300));
  INV_X1    g1100(.A(G384), .ZN(new_n1301));
  NOR3_X1   g1101(.A1(new_n1300), .A2(new_n1301), .A3(new_n1273), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1299), .A2(KEYINPUT60), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1298), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n690), .A3(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(G384), .B1(new_n1305), .B2(new_n1274), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1302), .A2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1295), .A2(new_n1297), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(KEYINPUT62), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1301), .B1(new_n1300), .B2(new_n1273), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1305), .A2(G384), .A3(new_n1274), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1296), .A2(G2897), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1311), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1313), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1310), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT61), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1296), .B1(new_n1287), .B2(new_n1294), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT62), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1319), .A2(new_n1320), .A3(new_n1307), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1309), .A2(new_n1317), .A3(new_n1318), .A4(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1278), .B1(new_n1054), .B2(new_n1084), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1279), .A2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1112), .B1(new_n1024), .B2(new_n1045), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1324), .B1(new_n1280), .B2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(G387), .A2(G390), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1024), .A2(new_n1045), .A3(new_n1112), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(G393), .A2(G396), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1054), .A2(new_n1278), .A3(new_n1084), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1327), .A2(new_n1328), .A3(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1326), .A2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1322), .A2(new_n1333), .ZN(new_n1334));
  OAI211_X1 g1134(.A(G2897), .B(new_n1296), .C1(new_n1302), .C2(new_n1306), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1311), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  OAI21_X1  g1137(.A(KEYINPUT63), .B1(new_n1337), .B2(new_n1319), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1338), .A2(new_n1308), .ZN(new_n1339));
  AND2_X1   g1139(.A1(new_n1326), .A2(new_n1332), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1295), .A2(KEYINPUT63), .A3(new_n1297), .A4(new_n1307), .ZN(new_n1341));
  AND2_X1   g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1339), .A2(new_n1342), .A3(new_n1318), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1334), .A2(new_n1343), .ZN(G405));
  INV_X1    g1144(.A(KEYINPUT127), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1307), .A2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1333), .A2(new_n1346), .ZN(new_n1347));
  OAI211_X1 g1147(.A(new_n1326), .B(new_n1332), .C1(new_n1345), .C2(new_n1307), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1307), .A2(new_n1345), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(G375), .A2(new_n1277), .ZN(new_n1351));
  AND3_X1   g1151(.A1(new_n1350), .A2(new_n1287), .A3(new_n1351), .ZN(new_n1352));
  XNOR2_X1  g1152(.A(new_n1349), .B(new_n1352), .ZN(G402));
endmodule


