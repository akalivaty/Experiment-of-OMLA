//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT89), .ZN(new_n190));
  NOR2_X1   g004(.A1(G237), .A2(G953), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n188), .A2(new_n190), .A3(G214), .A4(new_n191), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n191), .A2(G214), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(new_n188), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT68), .B(G131), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT17), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n194), .B(new_n195), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(KEYINPUT17), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT76), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n200), .B1(new_n202), .B2(KEYINPUT16), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n204), .A2(new_n201), .A3(KEYINPUT76), .A4(G125), .ZN(new_n205));
  INV_X1    g019(.A(G125), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G140), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n202), .A2(new_n207), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n203), .B(new_n205), .C1(new_n204), .C2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n209), .B(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n199), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(new_n208), .B(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT18), .A2(G131), .ZN(new_n214));
  XOR2_X1   g028(.A(new_n194), .B(new_n214), .Z(new_n215));
  AOI21_X1  g029(.A(new_n212), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  XOR2_X1   g030(.A(G113), .B(G122), .Z(new_n217));
  XNOR2_X1  g031(.A(new_n217), .B(KEYINPUT90), .ZN(new_n218));
  INV_X1    g032(.A(G104), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n218), .B(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n208), .B(KEYINPUT19), .ZN(new_n222));
  MUX2_X1   g036(.A(new_n209), .B(new_n222), .S(new_n210), .Z(new_n223));
  AOI22_X1  g037(.A1(new_n213), .A2(new_n215), .B1(new_n223), .B2(new_n198), .ZN(new_n224));
  OR2_X1    g038(.A1(new_n224), .A2(new_n220), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G475), .ZN(new_n227));
  INV_X1    g041(.A(G902), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT20), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT20), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n226), .A2(new_n231), .A3(new_n227), .A4(new_n228), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n216), .B(new_n220), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n228), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n230), .A2(new_n232), .B1(G475), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G953), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G952), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n237), .B1(G234), .B2(G237), .ZN(new_n238));
  XOR2_X1   g052(.A(KEYINPUT21), .B(G898), .Z(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(G234), .A2(G237), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(G902), .A3(G953), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n238), .B1(new_n240), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  XOR2_X1   g059(.A(KEYINPUT9), .B(G234), .Z(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G217), .ZN(new_n248));
  NOR3_X1   g062(.A1(new_n247), .A2(new_n248), .A3(G953), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G122), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT91), .B1(new_n251), .B2(G116), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT91), .ZN(new_n253));
  INV_X1    g067(.A(G116), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(G122), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G107), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n254), .A2(G122), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n256), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(G128), .B(G143), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n262), .B(G134), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT93), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n252), .A2(new_n255), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT14), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n264), .B(new_n259), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n266), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n266), .B1(new_n252), .B2(new_n255), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT93), .B1(new_n269), .B2(new_n258), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  AOI211_X1 g085(.A(new_n261), .B(new_n263), .C1(new_n271), .C2(G107), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n257), .B1(new_n256), .B2(new_n259), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT92), .B1(new_n261), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n273), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT92), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n276), .A3(new_n260), .ZN(new_n277));
  INV_X1    g091(.A(G134), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n262), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G128), .ZN(new_n280));
  NOR3_X1   g094(.A1(new_n280), .A2(KEYINPUT13), .A3(G143), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n281), .B1(new_n262), .B2(KEYINPUT13), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n279), .B1(G134), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n274), .A2(new_n277), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n250), .B1(new_n272), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n263), .B1(new_n271), .B2(G107), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n260), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(new_n284), .A3(new_n249), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n286), .A2(new_n289), .A3(KEYINPUT94), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT94), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n291), .B(new_n250), .C1(new_n272), .C2(new_n285), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n290), .A2(new_n228), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G478), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT95), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(KEYINPUT15), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(KEYINPUT15), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n294), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  OR2_X1    g113(.A1(new_n293), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n293), .A2(new_n299), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n235), .A2(new_n245), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G214), .B1(G237), .B2(G902), .ZN(new_n305));
  XOR2_X1   g119(.A(new_n305), .B(KEYINPUT84), .Z(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(G210), .B1(G237), .B2(G902), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  OR2_X1    g123(.A1(new_n280), .A2(KEYINPUT1), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(new_n189), .A3(G146), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n210), .A2(G143), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n189), .A2(G146), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI221_X1 g128(.A(new_n311), .B1(G128), .B2(new_n312), .C1(new_n314), .C2(new_n310), .ZN(new_n315));
  NAND2_X1  g129(.A1(KEYINPUT0), .A2(G128), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(KEYINPUT65), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT65), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(KEYINPUT0), .A3(G128), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  OR2_X1    g135(.A1(KEYINPUT0), .A2(G128), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(new_n314), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT66), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n321), .A2(new_n314), .A3(KEYINPUT66), .A4(new_n322), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n317), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  MUX2_X1   g141(.A(new_n315), .B(new_n327), .S(G125), .Z(new_n328));
  NAND2_X1  g142(.A1(new_n236), .A2(G224), .ZN(new_n329));
  XOR2_X1   g143(.A(new_n328), .B(new_n329), .Z(new_n330));
  XOR2_X1   g144(.A(G110), .B(G122), .Z(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT3), .B1(new_n219), .B2(G107), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT3), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n257), .A3(G104), .ZN(new_n335));
  INV_X1    g149(.A(G101), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n219), .A2(G107), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n333), .A2(new_n335), .A3(new_n336), .A4(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT79), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n338), .B(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n337), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n219), .A2(G107), .ZN(new_n342));
  OAI21_X1  g156(.A(G101), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT85), .B(KEYINPUT5), .ZN(new_n345));
  INV_X1    g159(.A(G119), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G116), .ZN(new_n347));
  OAI21_X1  g161(.A(G113), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(G116), .B(G119), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n345), .ZN(new_n351));
  XOR2_X1   g165(.A(KEYINPUT2), .B(G113), .Z(new_n352));
  AOI22_X1  g166(.A1(new_n349), .A2(new_n351), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n344), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(new_n350), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT2), .B(G113), .ZN(new_n357));
  INV_X1    g171(.A(new_n347), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n346), .A2(G116), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n338), .A2(new_n339), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n338), .A2(new_n339), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT4), .ZN(new_n364));
  NOR3_X1   g178(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n333), .A2(new_n335), .A3(new_n337), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G101), .ZN(new_n367));
  NAND2_X1  g181(.A1(KEYINPUT78), .A2(KEYINPUT4), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n366), .A2(KEYINPUT78), .A3(KEYINPUT4), .A4(G101), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n361), .B1(new_n365), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT86), .B1(new_n355), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT86), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n354), .A2(new_n375), .A3(new_n372), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n332), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  OR2_X1    g191(.A1(new_n377), .A2(KEYINPUT6), .ZN(new_n378));
  NOR3_X1   g192(.A1(new_n355), .A2(new_n373), .A3(new_n331), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT6), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n330), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT7), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n328), .B1(KEYINPUT88), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n329), .A2(KEYINPUT7), .ZN(new_n384));
  XOR2_X1   g198(.A(new_n383), .B(new_n384), .Z(new_n385));
  AND2_X1   g199(.A1(new_n350), .A2(KEYINPUT5), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n344), .B(new_n356), .C1(new_n348), .C2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n387), .B1(new_n344), .B2(new_n353), .ZN(new_n388));
  XOR2_X1   g202(.A(KEYINPUT87), .B(KEYINPUT8), .Z(new_n389));
  XNOR2_X1  g203(.A(new_n331), .B(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n379), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n385), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n228), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n309), .B1(new_n381), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n381), .A2(new_n393), .A3(new_n309), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n307), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(G221), .B1(new_n247), .B2(G902), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n340), .A2(new_n315), .A3(new_n343), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT10), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n327), .B1(new_n365), .B2(new_n371), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n340), .A2(KEYINPUT10), .A3(new_n315), .A4(new_n343), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G137), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(KEYINPUT11), .A3(G134), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n278), .A2(G137), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n278), .A2(G137), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT67), .B1(new_n410), .B2(KEYINPUT11), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n405), .A2(G134), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT67), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT11), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n409), .A2(new_n411), .A3(new_n415), .A4(new_n195), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n413), .B1(new_n412), .B2(new_n414), .ZN(new_n417));
  AOI211_X1 g231(.A(KEYINPUT67), .B(KEYINPUT11), .C1(new_n405), .C2(G134), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n417), .A2(new_n418), .A3(new_n408), .ZN(new_n419));
  INV_X1    g233(.A(G131), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n416), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n404), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT80), .ZN(new_n423));
  INV_X1    g237(.A(new_n421), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n401), .A2(new_n402), .A3(new_n424), .A4(new_n403), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n422), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G110), .B(G140), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n236), .A2(G227), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n427), .B(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n404), .A2(KEYINPUT80), .A3(new_n421), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n426), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n344), .A2(new_n315), .ZN(new_n432));
  INV_X1    g246(.A(new_n399), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n421), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT12), .ZN(new_n435));
  INV_X1    g249(.A(new_n429), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT12), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n437), .B(new_n421), .C1(new_n432), .C2(new_n433), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n435), .A2(new_n436), .A3(new_n425), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n431), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT81), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n431), .A2(KEYINPUT81), .A3(new_n439), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(G469), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n435), .A2(new_n429), .A3(new_n425), .A4(new_n438), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n446), .A2(KEYINPUT82), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n426), .A2(new_n436), .A3(new_n430), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(KEYINPUT82), .A3(new_n446), .ZN(new_n449));
  INV_X1    g263(.A(G469), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n447), .A2(new_n449), .A3(new_n450), .A4(new_n228), .ZN(new_n451));
  NAND2_X1  g265(.A1(G469), .A2(G902), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n398), .B1(new_n445), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT83), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT83), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n456), .B(new_n398), .C1(new_n445), .C2(new_n453), .ZN(new_n457));
  AOI211_X1 g271(.A(new_n304), .B(new_n397), .C1(new_n455), .C2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G472), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n327), .A2(new_n421), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n412), .A2(new_n407), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n315), .B(new_n416), .C1(new_n420), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(KEYINPUT30), .B1(new_n463), .B2(KEYINPUT64), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT64), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT30), .ZN(new_n466));
  AOI211_X1 g280(.A(new_n465), .B(new_n466), .C1(new_n460), .C2(new_n462), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n361), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT69), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT70), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n361), .B(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n460), .A2(new_n472), .A3(new_n462), .ZN(new_n473));
  XOR2_X1   g287(.A(KEYINPUT26), .B(G101), .Z(new_n474));
  NAND2_X1  g288(.A1(new_n191), .A2(G210), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n476), .B(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(KEYINPUT69), .B(new_n361), .C1(new_n464), .C2(new_n467), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n470), .A2(new_n473), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT31), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT28), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n473), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n460), .A2(new_n472), .A3(KEYINPUT28), .A4(new_n462), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n463), .A2(new_n361), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n478), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n489), .B1(new_n481), .B2(KEYINPUT31), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n459), .B(new_n228), .C1(new_n483), .C2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT72), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT75), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT32), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(KEYINPUT75), .A2(KEYINPUT32), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT29), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(new_n488), .B2(new_n478), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n470), .A2(new_n480), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n473), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n500), .B1(new_n502), .B2(new_n478), .ZN(new_n503));
  INV_X1    g317(.A(new_n472), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT73), .B1(new_n463), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n505), .A2(new_n485), .A3(new_n486), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n460), .A2(new_n472), .A3(KEYINPUT73), .A4(new_n462), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(KEYINPUT29), .A3(new_n479), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n228), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT74), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT74), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n512), .A3(new_n228), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(G472), .B1(new_n503), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n493), .A2(KEYINPUT75), .A3(KEYINPUT32), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n498), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n346), .A2(G128), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n518), .A2(KEYINPUT23), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(KEYINPUT23), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n519), .B(new_n520), .C1(G119), .C2(new_n280), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(G110), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT24), .B(G110), .Z(new_n523));
  XNOR2_X1  g337(.A(G119), .B(G128), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n211), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  OAI22_X1  g340(.A1(new_n521), .A2(G110), .B1(new_n524), .B2(new_n523), .ZN(new_n527));
  OR2_X1    g341(.A1(new_n209), .A2(new_n210), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n527), .B(new_n528), .C1(G146), .C2(new_n208), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT22), .B(G137), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(KEYINPUT77), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n236), .A2(G221), .A3(G234), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n530), .B(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(G902), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(KEYINPUT25), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n248), .B1(G234), .B2(new_n228), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n536), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n539), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n458), .A2(new_n517), .A3(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(G101), .ZN(G3));
  NOR2_X1   g358(.A1(new_n294), .A2(G902), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n249), .B1(new_n288), .B2(new_n284), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n289), .B1(new_n547), .B2(KEYINPUT98), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT98), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT33), .B1(new_n286), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT96), .B(KEYINPUT33), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n290), .A2(new_n292), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT97), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT97), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n290), .A2(new_n555), .A3(new_n292), .A4(new_n552), .ZN(new_n556));
  AOI211_X1 g370(.A(new_n546), .B(new_n551), .C1(new_n554), .C2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT99), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n293), .A2(new_n558), .A3(new_n294), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n558), .B1(new_n293), .B2(new_n294), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT100), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n554), .A2(new_n556), .ZN(new_n563));
  INV_X1    g377(.A(new_n551), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n545), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n560), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n293), .A2(new_n558), .A3(new_n294), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT100), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n565), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n235), .B1(new_n562), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n572), .A2(new_n397), .A3(new_n244), .ZN(new_n573));
  OR2_X1    g387(.A1(new_n481), .A2(KEYINPUT31), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n574), .A2(new_n482), .A3(new_n489), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n228), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(G472), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n491), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n541), .B1(new_n455), .B2(new_n457), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n573), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  XOR2_X1   g395(.A(KEYINPUT34), .B(G104), .Z(new_n582));
  XNOR2_X1  g396(.A(new_n581), .B(new_n582), .ZN(G6));
  INV_X1    g397(.A(new_n381), .ZN(new_n584));
  INV_X1    g398(.A(new_n393), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n585), .A3(new_n308), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n306), .B1(new_n586), .B2(new_n394), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n234), .A2(G475), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT101), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT101), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n234), .A2(new_n590), .A3(G475), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n589), .A2(new_n591), .B1(new_n230), .B2(new_n232), .ZN(new_n592));
  XOR2_X1   g406(.A(new_n244), .B(KEYINPUT102), .Z(new_n593));
  AND4_X1   g407(.A1(new_n587), .A2(new_n592), .A3(new_n302), .A4(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n580), .A2(new_n594), .A3(new_n579), .ZN(new_n595));
  XOR2_X1   g409(.A(KEYINPUT35), .B(G107), .Z(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(G9));
  NOR2_X1   g411(.A1(new_n534), .A2(KEYINPUT36), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n530), .B(new_n598), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n599), .B(new_n228), .C1(new_n248), .C2(G234), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n539), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n458), .A2(new_n579), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT37), .ZN(new_n603));
  XOR2_X1   g417(.A(new_n603), .B(G110), .Z(G12));
  NAND2_X1  g418(.A1(new_n455), .A2(new_n457), .ZN(new_n605));
  INV_X1    g419(.A(new_n238), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n606), .B1(G900), .B2(new_n242), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n592), .A2(new_n607), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n608), .A2(new_n302), .ZN(new_n609));
  INV_X1    g423(.A(new_n601), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n397), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n517), .A2(new_n605), .A3(new_n609), .A4(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(G128), .ZN(G30));
  XNOR2_X1  g427(.A(new_n607), .B(KEYINPUT39), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n605), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT40), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n502), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n478), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n505), .A2(new_n473), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n620), .A2(new_n507), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n228), .B1(new_n621), .B2(new_n479), .ZN(new_n622));
  OAI21_X1  g436(.A(G472), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n498), .A2(new_n516), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT38), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n586), .A2(new_n394), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n627), .B1(new_n586), .B2(new_n394), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT103), .B1(new_n395), .B2(new_n396), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n586), .A2(new_n394), .A3(new_n627), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n631), .A2(KEYINPUT38), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n625), .A2(new_n634), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n601), .A2(new_n235), .A3(new_n303), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n617), .A2(new_n635), .A3(new_n307), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G143), .ZN(G45));
  AND3_X1   g452(.A1(new_n571), .A2(KEYINPUT104), .A3(new_n607), .ZN(new_n639));
  AOI21_X1  g453(.A(KEYINPUT104), .B1(new_n571), .B2(new_n607), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n641), .A2(new_n517), .A3(new_n605), .A4(new_n611), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT105), .B(G146), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G48));
  AND2_X1   g458(.A1(new_n447), .A2(new_n449), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n228), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(G469), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n647), .A2(new_n398), .A3(new_n451), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n517), .A2(new_n542), .A3(new_n573), .A4(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT41), .B(G113), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G15));
  NAND4_X1  g465(.A1(new_n517), .A2(new_n542), .A3(new_n594), .A4(new_n648), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G116), .ZN(G18));
  NOR2_X1   g467(.A1(new_n304), .A2(new_n610), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n647), .A2(new_n451), .ZN(new_n655));
  INV_X1    g469(.A(new_n398), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n397), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n517), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G119), .ZN(G21));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n508), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n478), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n482), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT107), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n662), .A2(new_n665), .A3(new_n482), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n664), .A2(new_n574), .A3(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(G472), .A2(G902), .ZN(new_n668));
  AOI221_X4 g482(.A(new_n541), .B1(G472), .B2(new_n576), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n587), .A2(new_n593), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n235), .A2(new_n303), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n669), .A2(new_n670), .A3(new_n671), .A4(new_n648), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G122), .ZN(G24));
  NAND2_X1  g487(.A1(new_n667), .A2(new_n668), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n674), .A2(new_n577), .A3(new_n601), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n641), .A2(new_n675), .A3(new_n657), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G125), .ZN(G27));
  INV_X1    g491(.A(KEYINPUT42), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n440), .A2(G469), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n451), .A2(new_n452), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n398), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n395), .A2(new_n396), .A3(new_n306), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n517), .A2(new_n542), .A3(new_n682), .A4(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n641), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n678), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n491), .A2(new_n495), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n515), .A2(KEYINPUT32), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n687), .B1(new_n688), .B2(new_n491), .ZN(new_n689));
  OAI21_X1  g503(.A(KEYINPUT108), .B1(new_n689), .B2(new_n541), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n691));
  INV_X1    g505(.A(new_n576), .ZN(new_n692));
  AOI22_X1  g506(.A1(new_n692), .A2(new_n459), .B1(new_n515), .B2(KEYINPUT32), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n691), .B(new_n542), .C1(new_n693), .C2(new_n687), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n639), .A2(new_n640), .A3(new_n681), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n695), .A2(KEYINPUT42), .A3(new_n696), .A4(new_n683), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n686), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G131), .ZN(G33));
  INV_X1    g513(.A(new_n609), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n684), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n278), .ZN(G36));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n431), .A2(KEYINPUT81), .A3(new_n439), .ZN(new_n704));
  AOI21_X1  g518(.A(KEYINPUT81), .B1(new_n431), .B2(new_n439), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n703), .B(G469), .C1(new_n706), .C2(KEYINPUT45), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n440), .A2(KEYINPUT45), .ZN(new_n708));
  NAND2_X1  g522(.A1(KEYINPUT45), .A2(G469), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n444), .A2(KEYINPUT109), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT46), .B1(new_n711), .B2(new_n452), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n712), .A2(KEYINPUT111), .ZN(new_n713));
  INV_X1    g527(.A(new_n451), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n711), .A2(KEYINPUT46), .A3(new_n452), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT110), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n711), .A2(KEYINPUT110), .A3(KEYINPUT46), .A4(new_n452), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n712), .A2(KEYINPUT111), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n713), .A2(new_n717), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n398), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n683), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n562), .A2(new_n570), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n235), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n724), .A2(KEYINPUT43), .A3(new_n235), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n578), .A3(new_n601), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n723), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OR2_X1    g546(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n722), .A2(new_n614), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G137), .ZN(G39));
  NOR3_X1   g549(.A1(new_n517), .A2(new_n542), .A3(new_n723), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n720), .A2(KEYINPUT47), .A3(new_n398), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT47), .B1(new_n720), .B2(new_n398), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n641), .B(new_n736), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G140), .ZN(G42));
  AND3_X1   g554(.A1(new_n648), .A2(new_n238), .A3(new_n683), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n625), .A2(new_n542), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n571), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n695), .A2(new_n729), .A3(new_n741), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n744), .A2(KEYINPUT48), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(KEYINPUT48), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n237), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT47), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n721), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n720), .A2(KEYINPUT47), .A3(new_n398), .ZN(new_n750));
  INV_X1    g564(.A(new_n655), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n656), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n606), .B1(new_n727), .B2(new_n728), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n669), .A3(new_n683), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n307), .B1(new_n630), .B2(new_n633), .ZN(new_n759));
  AND4_X1   g573(.A1(new_n542), .A2(new_n674), .A3(new_n577), .A4(new_n648), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n759), .A2(new_n760), .A3(new_n754), .A4(KEYINPUT50), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n761), .A2(KEYINPUT117), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(KEYINPUT117), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n759), .A2(new_n760), .A3(new_n754), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n764), .A2(KEYINPUT116), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT116), .B1(new_n764), .B2(new_n765), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n762), .B(new_n763), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n675), .A2(new_n741), .A3(new_n729), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n742), .A2(new_n235), .A3(new_n562), .A4(new_n570), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(KEYINPUT115), .B(KEYINPUT51), .C1(new_n758), .C2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n757), .A2(new_n769), .A3(new_n768), .A4(new_n770), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT51), .B1(new_n774), .B2(KEYINPUT115), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n743), .B(new_n747), .C1(new_n773), .C2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n701), .B1(new_n686), .B2(new_n697), .ZN(new_n779));
  INV_X1    g593(.A(new_n607), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n681), .A2(new_n601), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n587), .A2(new_n671), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n784), .B1(new_n781), .B2(new_n782), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n624), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n642), .A2(new_n612), .A3(new_n676), .A4(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(KEYINPUT114), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n649), .A2(new_n652), .A3(new_n658), .A4(new_n672), .ZN(new_n790));
  INV_X1    g604(.A(new_n235), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n572), .B1(new_n303), .B2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n792), .A2(new_n580), .A3(new_n579), .A4(new_n670), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n543), .A2(new_n602), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n641), .A2(new_n577), .A3(new_n674), .A4(new_n682), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n517), .A2(new_n605), .A3(new_n303), .A4(new_n608), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(new_n601), .A3(new_n683), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n779), .A2(new_n789), .A3(new_n795), .A4(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n612), .A2(new_n676), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n801), .A2(KEYINPUT52), .A3(new_n642), .A4(new_n786), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n787), .A2(new_n788), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n778), .B1(new_n800), .B2(new_n805), .ZN(new_n806));
  AOI211_X1 g620(.A(new_n610), .B(new_n723), .C1(new_n796), .C2(new_n797), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n807), .A2(new_n790), .A3(new_n794), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n802), .A2(new_n804), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n808), .A2(new_n809), .A3(new_n778), .A4(new_n779), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n777), .B1(new_n806), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT53), .B1(new_n800), .B2(new_n805), .ZN(new_n813));
  AND4_X1   g627(.A1(KEYINPUT53), .A2(new_n808), .A3(new_n809), .A4(new_n779), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT54), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n754), .A2(new_n657), .A3(new_n669), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n812), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  OAI22_X1  g631(.A1(new_n776), .A2(new_n817), .B1(G952), .B2(G953), .ZN(new_n818));
  XNOR2_X1  g632(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n819));
  AOI211_X1 g633(.A(new_n656), .B(new_n725), .C1(new_n751), .C2(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n820), .A2(new_n307), .A3(new_n634), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n655), .B1(KEYINPUT112), .B2(KEYINPUT49), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n821), .A2(new_n542), .A3(new_n625), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n818), .A2(new_n823), .ZN(G75));
  AND3_X1   g638(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n779), .A2(new_n789), .A3(new_n795), .A4(new_n799), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT53), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(G210), .A3(G902), .A4(new_n810), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT56), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT118), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n236), .A2(G952), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n828), .A2(KEYINPUT118), .A3(new_n829), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n378), .A2(new_n380), .A3(new_n330), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n584), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT55), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n835), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n828), .A2(KEYINPUT118), .A3(new_n829), .A4(new_n837), .ZN(new_n838));
  AOI211_X1 g652(.A(new_n830), .B(new_n831), .C1(new_n836), .C2(new_n838), .ZN(G51));
  OR2_X1    g653(.A1(new_n452), .A2(KEYINPUT57), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n452), .A2(KEYINPUT57), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n827), .A2(KEYINPUT54), .A3(new_n810), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT54), .B1(new_n827), .B2(new_n810), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n840), .B(new_n841), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n645), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n711), .B(KEYINPUT119), .Z(new_n846));
  NAND4_X1  g660(.A1(new_n827), .A2(G902), .A3(new_n810), .A4(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n831), .B1(new_n845), .B2(new_n847), .ZN(G54));
  NAND4_X1  g662(.A1(new_n827), .A2(KEYINPUT58), .A3(G902), .A4(new_n810), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n227), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT120), .B1(new_n850), .B2(new_n226), .ZN(new_n851));
  INV_X1    g665(.A(new_n226), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n852), .B1(new_n849), .B2(new_n227), .ZN(new_n853));
  INV_X1    g667(.A(new_n831), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n849), .A2(new_n856), .A3(new_n227), .A4(new_n852), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n851), .A2(new_n855), .A3(new_n857), .ZN(G60));
  NAND2_X1  g672(.A1(new_n563), .A2(new_n564), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(G478), .A2(G902), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n861), .B(KEYINPUT59), .Z(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n860), .B(new_n863), .C1(new_n842), .C2(new_n843), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n862), .B1(new_n812), .B2(new_n815), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n864), .B(new_n854), .C1(new_n865), .C2(new_n860), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(G63));
  NAND2_X1  g681(.A1(G217), .A2(G902), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT60), .Z(new_n869));
  NAND3_X1  g683(.A1(new_n827), .A2(new_n810), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n535), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n827), .A2(new_n599), .A3(new_n810), .A4(new_n869), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n854), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT61), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n871), .A2(KEYINPUT61), .A3(new_n854), .A4(new_n872), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(G66));
  INV_X1    g691(.A(G224), .ZN(new_n878));
  OAI21_X1  g692(.A(G953), .B1(new_n240), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n879), .B1(new_n795), .B2(G953), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n378), .B(new_n380), .C1(G898), .C2(new_n236), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT121), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n880), .B(new_n882), .ZN(G69));
  NAND3_X1  g697(.A1(new_n642), .A2(new_n612), .A3(new_n676), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT122), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n642), .A2(new_n612), .A3(new_n676), .A4(KEYINPUT122), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n739), .A2(new_n734), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n784), .B1(new_n690), .B2(new_n694), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n722), .A2(new_n614), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n779), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT125), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n886), .A2(new_n887), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n685), .B1(new_n749), .B2(new_n750), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n894), .B2(new_n736), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT125), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n890), .A2(new_n779), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n895), .A2(new_n896), .A3(new_n734), .A4(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n892), .A2(new_n898), .A3(new_n236), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n464), .A2(new_n467), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(new_n222), .Z(new_n901));
  NAND2_X1  g715(.A1(G900), .A2(G953), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n904));
  INV_X1    g718(.A(new_n637), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n904), .B1(new_n893), .B2(new_n905), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n886), .A2(new_n637), .A3(KEYINPUT62), .A4(new_n887), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n739), .A2(new_n734), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n517), .A2(new_n542), .A3(new_n683), .ZN(new_n910));
  INV_X1    g724(.A(new_n615), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n910), .A2(new_n911), .A3(new_n792), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n908), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n236), .ZN(new_n914));
  INV_X1    g728(.A(new_n901), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n903), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n236), .B1(G227), .B2(G900), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n914), .A2(new_n920), .A3(new_n915), .ZN(new_n921));
  INV_X1    g735(.A(new_n912), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n906), .B2(new_n907), .ZN(new_n923));
  AOI21_X1  g737(.A(G953), .B1(new_n923), .B2(new_n909), .ZN(new_n924));
  OAI21_X1  g738(.A(KEYINPUT123), .B1(new_n924), .B2(new_n901), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n918), .B(KEYINPUT124), .Z(new_n926));
  NAND4_X1  g740(.A1(new_n903), .A2(new_n921), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n919), .A2(new_n927), .ZN(G72));
  NAND4_X1  g742(.A1(new_n908), .A2(new_n795), .A3(new_n909), .A4(new_n912), .ZN(new_n929));
  XNOR2_X1  g743(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n459), .A2(new_n228), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n930), .B(new_n931), .Z(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(KEYINPUT127), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n929), .A2(new_n936), .A3(new_n933), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n935), .A2(new_n619), .A3(new_n937), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n892), .A2(new_n898), .A3(new_n795), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n478), .B(new_n618), .C1(new_n939), .C2(new_n932), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n813), .A2(new_n814), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n502), .A2(new_n478), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n932), .B1(new_n942), .B2(new_n481), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n831), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n938), .A2(new_n940), .A3(new_n944), .ZN(G57));
endmodule


