//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n800, new_n802, new_n803, new_n804, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913;
  XOR2_X1   g000(.A(G15gat), .B(G22gat), .Z(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT90), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(new_n207), .B2(new_n202), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT91), .ZN(new_n209));
  AOI21_X1  g008(.A(G8gat), .B1(new_n204), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n208), .B(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G71gat), .A2(G78gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT94), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OR2_X1    g013(.A1(G71gat), .A2(G78gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(KEYINPUT94), .A2(G71gat), .A3(G78gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT95), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT9), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n212), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G57gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(G64gat), .ZN(new_n222));
  INV_X1    g021(.A(G64gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n223), .A2(G57gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n220), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT95), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n214), .A2(new_n215), .A3(new_n226), .A4(new_n216), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n218), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n212), .B1(new_n215), .B2(new_n219), .ZN(new_n229));
  OR3_X1    g028(.A1(new_n223), .A2(KEYINPUT96), .A3(G57gat), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT96), .B1(new_n223), .B2(G57gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n229), .B1(new_n232), .B2(new_n222), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n228), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT21), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n211), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G183gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G127gat), .B(G155gat), .ZN(new_n241));
  INV_X1    g040(.A(G211gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n234), .A2(KEYINPUT21), .ZN(new_n245));
  NAND2_X1  g044(.A1(G231gat), .A2(G233gat), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n246), .B(KEYINPUT97), .Z(new_n247));
  XNOR2_X1  g046(.A(new_n245), .B(new_n247), .ZN(new_n248));
  OR2_X1    g047(.A1(new_n238), .A2(new_n239), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n238), .A2(new_n239), .ZN(new_n250));
  INV_X1    g049(.A(new_n243), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n244), .A2(new_n248), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n248), .B1(new_n244), .B2(new_n252), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G134gat), .B(G162gat), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT100), .ZN(new_n260));
  INV_X1    g059(.A(G85gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT98), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n262), .A2(G92gat), .ZN(new_n263));
  INV_X1    g062(.A(G92gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(KEYINPUT98), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n261), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G99gat), .B(G106gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(G99gat), .A2(G106gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT8), .ZN(new_n269));
  AND3_X1   g068(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n266), .A2(new_n267), .A3(new_n269), .A4(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT99), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n264), .A2(KEYINPUT98), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n262), .A2(G92gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n278), .A2(new_n261), .B1(KEYINPUT8), .B2(new_n268), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n267), .B1(new_n279), .B2(new_n272), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n266), .A2(new_n269), .A3(new_n272), .ZN(new_n282));
  INV_X1    g081(.A(new_n267), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(KEYINPUT99), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n260), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT98), .B(G92gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n269), .B1(new_n287), .B2(G85gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n272), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n283), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(new_n274), .A3(new_n273), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(KEYINPUT100), .A3(new_n284), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n286), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G50gat), .ZN(new_n294));
  OR2_X1    g093(.A1(new_n294), .A2(G43gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(G43gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(KEYINPUT15), .A3(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT89), .B(G43gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n294), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT15), .B1(new_n299), .B2(new_n295), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT14), .ZN(new_n301));
  OR3_X1    g100(.A1(new_n301), .A2(G29gat), .A3(G36gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n301), .B1(G29gat), .B2(G36gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT88), .B(G29gat), .ZN(new_n304));
  INV_X1    g103(.A(G36gat), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n302), .B(new_n303), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n297), .B1(new_n300), .B2(new_n306), .ZN(new_n307));
  OR2_X1    g106(.A1(new_n306), .A2(new_n297), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n308), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT17), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT17), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n307), .A2(new_n313), .A3(new_n308), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n286), .A2(new_n312), .A3(new_n314), .A4(new_n292), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n309), .A2(new_n310), .A3(new_n315), .ZN(new_n316));
  XOR2_X1   g115(.A(G190gat), .B(G218gat), .Z(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n259), .B1(new_n319), .B2(KEYINPUT101), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n316), .A2(new_n318), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n309), .A2(new_n317), .A3(new_n310), .A4(new_n315), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n321), .A2(KEYINPUT101), .A3(new_n322), .A4(new_n259), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n290), .A2(KEYINPUT102), .A3(new_n273), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT102), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n282), .A2(new_n328), .A3(new_n283), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n234), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n291), .A2(new_n284), .B1(new_n233), .B2(new_n228), .ZN(new_n331));
  INV_X1    g130(.A(G230gat), .ZN(new_n332));
  INV_X1    g131(.A(G233gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NOR3_X1   g134(.A1(new_n330), .A2(new_n331), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT103), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n228), .A2(new_n233), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(new_n281), .B2(new_n285), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n234), .A2(new_n327), .A3(new_n329), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT10), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT10), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n345), .B1(new_n286), .B2(new_n292), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n335), .B1(new_n342), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G120gat), .B(G148gat), .ZN(new_n348));
  INV_X1    g147(.A(G176gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G204gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n337), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n338), .A2(new_n347), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n343), .B1(new_n330), .B2(new_n331), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n291), .A2(KEYINPUT100), .A3(new_n284), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT100), .B1(new_n291), .B2(new_n284), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n344), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n334), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n352), .B1(new_n360), .B2(new_n336), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n256), .A2(new_n326), .A3(new_n362), .ZN(new_n363));
  OR2_X1    g162(.A1(new_n211), .A2(new_n311), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n312), .A2(new_n211), .A3(new_n314), .ZN(new_n365));
  NAND2_X1  g164(.A1(G229gat), .A2(G233gat), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT18), .A4(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(new_n366), .B(KEYINPUT13), .Z(new_n368));
  AND2_X1   g167(.A1(new_n211), .A2(new_n311), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n211), .A2(new_n311), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(new_n371), .A3(KEYINPUT92), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT11), .B(G169gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(G197gat), .ZN(new_n374));
  XOR2_X1   g173(.A(G113gat), .B(G141gat), .Z(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(KEYINPUT12), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT18), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n371), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n372), .B(new_n378), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n367), .A2(new_n371), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n385), .B(new_n381), .C1(KEYINPUT92), .C2(new_n377), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT93), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT93), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n363), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT0), .B(G57gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n395), .B(G85gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(G1gat), .B(G29gat), .ZN(new_n397));
  XOR2_X1   g196(.A(new_n396), .B(new_n397), .Z(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G127gat), .B(G134gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(KEYINPUT67), .ZN(new_n401));
  XNOR2_X1  g200(.A(G113gat), .B(G120gat), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n401), .B1(KEYINPUT1), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT68), .B(G120gat), .ZN(new_n405));
  INV_X1    g204(.A(G113gat), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n406), .A2(G120gat), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n404), .B(new_n400), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT78), .B(G141gat), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n411), .A2(KEYINPUT79), .A3(G148gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(G155gat), .A2(G162gat), .ZN(new_n413));
  INV_X1    g212(.A(G155gat), .ZN(new_n414));
  INV_X1    g213(.A(G162gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n413), .B1(new_n416), .B2(KEYINPUT2), .ZN(new_n417));
  INV_X1    g216(.A(new_n411), .ZN(new_n418));
  INV_X1    g217(.A(G148gat), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT79), .ZN(new_n421));
  INV_X1    g220(.A(G141gat), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(G148gat), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n412), .B(new_n417), .C1(new_n420), .C2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT76), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n416), .B(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G141gat), .B(G148gat), .ZN(new_n427));
  XOR2_X1   g226(.A(KEYINPUT77), .B(KEYINPUT2), .Z(new_n428));
  OAI211_X1 g227(.A(new_n426), .B(new_n413), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n410), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n403), .A2(new_n424), .A3(new_n429), .A4(new_n409), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(G225gat), .A2(G233gat), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT5), .ZN(new_n437));
  INV_X1    g236(.A(new_n432), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT4), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(KEYINPUT80), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n430), .A2(KEYINPUT3), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT3), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n424), .A2(new_n429), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n441), .A2(new_n410), .A3(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n438), .A2(new_n439), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT80), .B1(new_n432), .B2(KEYINPUT4), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n435), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT81), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n445), .A2(KEYINPUT81), .A3(new_n448), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n437), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n432), .B(KEYINPUT4), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n444), .ZN(new_n455));
  OR3_X1    g254(.A1(new_n455), .A2(KEYINPUT5), .A3(new_n435), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n399), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n437), .ZN(new_n459));
  INV_X1    g258(.A(new_n452), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT81), .B1(new_n445), .B2(new_n448), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(new_n398), .A3(new_n456), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n458), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(KEYINPUT6), .B(new_n399), .C1(new_n453), .C2(new_n457), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n410), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n469));
  INV_X1    g268(.A(G190gat), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n469), .B1(new_n237), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(G169gat), .A2(G176gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT23), .ZN(new_n475));
  INV_X1    g274(.A(G169gat), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT23), .B1(new_n476), .B2(new_n349), .ZN(new_n477));
  INV_X1    g276(.A(new_n474), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n473), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT25), .ZN(new_n481));
  XNOR2_X1  g280(.A(KEYINPUT27), .B(G183gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n470), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT28), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(G183gat), .A2(G190gat), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n478), .A2(KEYINPUT26), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT66), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n478), .A2(KEYINPUT26), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT66), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n490), .B1(G169gat), .B2(G176gat), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n488), .B(new_n489), .C1(new_n487), .C2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n485), .A2(new_n486), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n469), .B1(KEYINPUT64), .B2(new_n472), .ZN(new_n494));
  OAI221_X1 g293(.A(new_n494), .B1(KEYINPUT64), .B2(new_n472), .C1(G183gat), .C2(G190gat), .ZN(new_n495));
  XOR2_X1   g294(.A(new_n475), .B(KEYINPUT65), .Z(new_n496));
  INV_X1    g295(.A(KEYINPUT25), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n495), .A2(new_n496), .A3(new_n497), .A4(new_n479), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n468), .A2(new_n481), .A3(new_n493), .A4(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n493), .A2(new_n481), .A3(new_n498), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n410), .ZN(new_n501));
  AND2_X1   g300(.A1(G227gat), .A2(G233gat), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n499), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT71), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT34), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G15gat), .B(G43gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(G71gat), .B(G99gat), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n509), .B(new_n510), .Z(new_n511));
  AOI21_X1  g310(.A(new_n503), .B1(new_n499), .B2(new_n501), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(KEYINPUT33), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT32), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n513), .A2(new_n515), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n508), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n506), .B(KEYINPUT34), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n513), .A2(new_n515), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n521), .A3(new_n516), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(G228gat), .A2(G233gat), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT22), .ZN(new_n526));
  INV_X1    g325(.A(G218gat), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n526), .B1(new_n242), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G197gat), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n529), .A2(new_n351), .ZN(new_n530));
  NOR2_X1   g329(.A1(G197gat), .A2(G204gat), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n532), .A2(KEYINPUT82), .ZN(new_n533));
  XNOR2_X1  g332(.A(G211gat), .B(G218gat), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n532), .A2(KEYINPUT82), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n532), .A2(KEYINPUT82), .A3(new_n534), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT29), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT83), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n537), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n442), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n541), .B1(new_n537), .B2(new_n540), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n430), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n443), .A2(new_n539), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT73), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT72), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n547), .B1(new_n532), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n535), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT72), .B1(new_n535), .B2(KEYINPUT73), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(new_n532), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n546), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n525), .B1(new_n545), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n442), .B1(new_n553), .B2(KEYINPUT29), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(new_n430), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(new_n554), .A3(new_n525), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(G22gat), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G78gat), .B(G106gat), .Z(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT31), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(new_n294), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G22gat), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n545), .A2(new_n554), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n558), .B(new_n566), .C1(new_n567), .C2(new_n525), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT84), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n568), .A2(new_n560), .A3(new_n569), .A4(new_n564), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n555), .A2(new_n559), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n571), .B(new_n566), .C1(KEYINPUT84), .C2(new_n563), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n565), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  NOR3_X1   g372(.A1(new_n523), .A2(KEYINPUT35), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G8gat), .B(G36gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(new_n223), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(new_n264), .ZN(new_n577));
  INV_X1    g376(.A(new_n553), .ZN(new_n578));
  NAND2_X1  g377(.A1(G226gat), .A2(G233gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n500), .B1(KEYINPUT29), .B2(new_n580), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n493), .A2(new_n579), .A3(new_n481), .A4(new_n498), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n578), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n581), .A2(new_n578), .A3(new_n582), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(KEYINPUT74), .A3(new_n585), .ZN(new_n586));
  AOI211_X1 g385(.A(KEYINPUT74), .B(new_n578), .C1(new_n581), .C2(new_n582), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n577), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT30), .B1(new_n589), .B2(KEYINPUT75), .ZN(new_n590));
  INV_X1    g389(.A(new_n577), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n585), .A2(KEYINPUT74), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n592), .A2(new_n583), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n591), .B1(new_n593), .B2(new_n587), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT75), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT30), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n586), .A2(new_n588), .A3(new_n577), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n590), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n467), .A2(new_n574), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT87), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n508), .A2(new_n521), .A3(KEYINPUT70), .A4(new_n516), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT70), .ZN(new_n604));
  OAI22_X1  g403(.A1(new_n520), .A2(new_n604), .B1(new_n517), .B2(new_n518), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n573), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n467), .A2(new_n606), .A3(new_n600), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT35), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT87), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n467), .A2(new_n574), .A3(new_n609), .A4(new_n600), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n602), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n455), .A2(new_n435), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(KEYINPUT39), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n613), .A2(new_n399), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n612), .B(KEYINPUT39), .C1(new_n435), .C2(new_n433), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(KEYINPUT40), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT40), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n599), .A2(new_n616), .A3(new_n458), .A4(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n573), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT37), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n622), .B1(new_n593), .B2(new_n587), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n586), .A2(KEYINPUT37), .A3(new_n588), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(new_n577), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n589), .B1(new_n625), .B2(KEYINPUT38), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n465), .A2(new_n626), .A3(new_n466), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT85), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n584), .A2(new_n628), .A3(new_n585), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n629), .B(KEYINPUT37), .C1(new_n628), .C2(new_n584), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT38), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n630), .A2(new_n623), .A3(new_n631), .A4(new_n577), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(KEYINPUT86), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n586), .A2(new_n588), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n591), .B1(new_n634), .B2(new_n622), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT86), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n635), .A2(new_n636), .A3(new_n631), .A4(new_n630), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n620), .B(new_n621), .C1(new_n627), .C2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n467), .A2(new_n600), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n573), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n605), .A2(new_n603), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT36), .ZN(new_n643));
  INV_X1    g442(.A(new_n523), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n643), .B1(KEYINPUT36), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n639), .A2(new_n641), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n394), .B1(new_n611), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n467), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g449(.A(KEYINPUT16), .B(G8gat), .Z(new_n651));
  NAND3_X1  g450(.A1(new_n647), .A2(new_n599), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n653));
  AND2_X1   g452(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n647), .A2(new_n599), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n656), .A2(KEYINPUT105), .A3(G8gat), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT105), .B1(new_n656), .B2(G8gat), .ZN(new_n658));
  OAI221_X1 g457(.A(new_n655), .B1(new_n653), .B2(new_n652), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n659), .B(KEYINPUT106), .Z(G1325gat));
  AOI21_X1  g459(.A(G15gat), .B1(new_n647), .B2(new_n644), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT107), .ZN(new_n662));
  INV_X1    g461(.A(new_n645), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n647), .A2(G15gat), .A3(new_n663), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n662), .A2(new_n664), .ZN(G1326gat));
  NAND2_X1  g464(.A1(new_n647), .A2(new_n573), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT43), .B(G22gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1327gat));
  AND2_X1   g467(.A1(new_n324), .A2(new_n325), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n669), .B1(new_n611), .B2(new_n646), .ZN(new_n670));
  INV_X1    g469(.A(new_n362), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n256), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n672), .A2(new_n392), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n670), .A2(new_n648), .A3(new_n304), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT45), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n670), .B(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n672), .A2(new_n388), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n648), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n675), .B1(new_n681), .B2(new_n304), .ZN(G1328gat));
  NAND2_X1  g481(.A1(new_n670), .A2(new_n673), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n683), .A2(G36gat), .A3(new_n600), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT46), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n679), .A2(new_n599), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n687), .B2(new_n305), .ZN(G1329gat));
  NAND4_X1  g487(.A1(new_n677), .A2(new_n663), .A3(new_n298), .A4(new_n678), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n683), .A2(new_n523), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n689), .B1(new_n298), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g491(.A1(new_n683), .A2(KEYINPUT108), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n670), .A2(new_n694), .A3(new_n673), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n695), .A2(new_n294), .A3(new_n573), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n611), .A2(new_n646), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n676), .B1(new_n697), .B2(new_n326), .ZN(new_n698));
  AOI211_X1 g497(.A(KEYINPUT44), .B(new_n669), .C1(new_n611), .C2(new_n646), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n573), .B(new_n678), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  AOI22_X1  g499(.A1(new_n693), .A2(new_n696), .B1(new_n700), .B2(G50gat), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n701), .A2(KEYINPUT48), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n677), .A2(new_n703), .A3(new_n573), .A4(new_n678), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n700), .A2(KEYINPUT109), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(new_n705), .A3(G50gat), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT110), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT48), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(new_n696), .B2(new_n693), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n706), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n707), .B1(new_n706), .B2(new_n709), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n702), .B1(new_n710), .B2(new_n711), .ZN(G1331gat));
  NOR2_X1   g511(.A1(new_n387), .A2(new_n671), .ZN(new_n713));
  AND4_X1   g512(.A1(new_n697), .A2(new_n669), .A3(new_n255), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n648), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(G57gat), .ZN(G1332gat));
  INV_X1    g515(.A(KEYINPUT49), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n714), .B(new_n599), .C1(new_n717), .C2(new_n223), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n223), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1333gat));
  INV_X1    g519(.A(G71gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n714), .A2(new_n721), .A3(new_n644), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n714), .A2(new_n663), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n723), .B2(new_n721), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n724), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g524(.A1(new_n714), .A2(new_n573), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g526(.A1(new_n670), .A2(new_n388), .A3(new_n256), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n728), .A2(KEYINPUT51), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(KEYINPUT51), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n467), .A2(G85gat), .A3(new_n671), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT111), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n713), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n255), .A2(new_n735), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n677), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n648), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n734), .B1(new_n739), .B2(new_n261), .ZN(G1336gat));
  OAI211_X1 g539(.A(new_n599), .B(new_n736), .C1(new_n698), .C2(new_n699), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n287), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT113), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT52), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n599), .A2(new_n264), .A3(new_n362), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT112), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n730), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n742), .ZN(new_n748));
  XOR2_X1   g547(.A(new_n744), .B(new_n748), .Z(G1337gat));
  INV_X1    g548(.A(G99gat), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n731), .A2(new_n750), .A3(new_n644), .A4(new_n362), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n737), .A2(new_n663), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n753), .B2(new_n750), .ZN(G1338gat));
  NAND3_X1  g553(.A1(new_n677), .A2(new_n573), .A3(new_n736), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G106gat), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n729), .A2(new_n573), .A3(new_n362), .A4(new_n730), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n757), .B2(G106gat), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(new_n757), .B2(G106gat), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n758), .A2(new_n760), .A3(KEYINPUT53), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762));
  OAI221_X1 g561(.A(new_n756), .B1(new_n759), .B2(new_n762), .C1(new_n757), .C2(G106gat), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(G1339gat));
  NOR2_X1   g563(.A1(new_n467), .A2(new_n599), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT54), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n353), .B1(new_n360), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n356), .A2(new_n359), .A3(new_n334), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n347), .A2(KEYINPUT54), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n768), .A2(new_n770), .A3(KEYINPUT55), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n771), .A2(new_n355), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n768), .A2(new_n770), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT115), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n776));
  AOI211_X1 g575(.A(new_n776), .B(KEYINPUT55), .C1(new_n768), .C2(new_n770), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n772), .B(new_n387), .C1(new_n775), .C2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n385), .A2(new_n377), .A3(new_n381), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n369), .A2(new_n370), .A3(new_n368), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n366), .B1(new_n364), .B2(new_n365), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n376), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n362), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n326), .B1(new_n778), .B2(new_n784), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n772), .B(new_n783), .C1(new_n775), .C2(new_n777), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(new_n669), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n256), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n255), .A2(new_n388), .A3(new_n669), .A4(new_n671), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n766), .B1(new_n790), .B2(new_n621), .ZN(new_n791));
  AOI211_X1 g590(.A(KEYINPUT116), .B(new_n573), .C1(new_n788), .C2(new_n789), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n644), .B(new_n765), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(G113gat), .B1(new_n793), .B2(new_n392), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n790), .A2(new_n606), .A3(new_n765), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(new_n406), .A3(new_n387), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(G1340gat));
  OAI21_X1  g596(.A(G120gat), .B1(new_n793), .B2(new_n671), .ZN(new_n798));
  INV_X1    g597(.A(new_n405), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n795), .A2(new_n799), .A3(new_n362), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(G1341gat));
  AOI21_X1  g600(.A(G127gat), .B1(new_n795), .B2(new_n255), .ZN(new_n802));
  INV_X1    g601(.A(G127gat), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n793), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n802), .B1(new_n804), .B2(new_n255), .ZN(G1342gat));
  INV_X1    g604(.A(G134gat), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n795), .A2(new_n806), .A3(new_n326), .ZN(new_n807));
  XOR2_X1   g606(.A(new_n807), .B(KEYINPUT56), .Z(new_n808));
  OAI21_X1  g607(.A(G134gat), .B1(new_n793), .B2(new_n669), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(G1343gat));
  AOI21_X1  g609(.A(new_n621), .B1(new_n788), .B2(new_n789), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n765), .A2(new_n645), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n814), .A2(G141gat), .A3(new_n392), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n784), .B(KEYINPUT117), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n773), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n768), .A2(new_n770), .A3(KEYINPUT118), .ZN(new_n821));
  XOR2_X1   g620(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n389), .A2(new_n391), .A3(new_n772), .A4(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n326), .B1(new_n818), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n256), .B1(new_n825), .B2(new_n787), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n789), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n573), .ZN(new_n828));
  AOI211_X1 g627(.A(new_n812), .B(new_n817), .C1(new_n828), .C2(KEYINPUT57), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n387), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n815), .B1(new_n830), .B2(new_n418), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n411), .B1(new_n829), .B2(new_n393), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n815), .A2(KEYINPUT58), .ZN(new_n834));
  OAI22_X1  g633(.A1(new_n831), .A2(new_n832), .B1(new_n833), .B2(new_n834), .ZN(G1344gat));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n363), .A2(new_n392), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n826), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n816), .B1(new_n838), .B2(new_n621), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n811), .A2(KEYINPUT57), .ZN(new_n842));
  OAI211_X1 g641(.A(KEYINPUT121), .B(new_n816), .C1(new_n838), .C2(new_n621), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n812), .A2(KEYINPUT120), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n812), .A2(KEYINPUT120), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n844), .A2(new_n362), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n836), .B1(new_n847), .B2(G148gat), .ZN(new_n848));
  AOI211_X1 g647(.A(KEYINPUT59), .B(new_n419), .C1(new_n829), .C2(new_n362), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n362), .A2(new_n419), .ZN(new_n850));
  OAI22_X1  g649(.A1(new_n848), .A2(new_n849), .B1(new_n814), .B2(new_n850), .ZN(G1345gat));
  NAND3_X1  g650(.A1(new_n829), .A2(G155gat), .A3(new_n255), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n414), .B1(new_n814), .B2(new_n256), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(G1346gat));
  NAND3_X1  g653(.A1(new_n829), .A2(G162gat), .A3(new_n326), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n415), .B1(new_n814), .B2(new_n669), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(G1347gat));
  NAND2_X1  g656(.A1(new_n790), .A2(new_n467), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT122), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n859), .A2(new_n606), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n599), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n861), .A2(G169gat), .A3(new_n388), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n648), .A2(new_n600), .A3(new_n523), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(new_n791), .B2(new_n792), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT123), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT123), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n866), .B(new_n863), .C1(new_n791), .C2(new_n792), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n476), .B1(new_n868), .B2(new_n393), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n862), .A2(new_n869), .ZN(G1348gat));
  OAI21_X1  g669(.A(new_n349), .B1(new_n861), .B2(new_n671), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n868), .A2(G176gat), .A3(new_n362), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(G1349gat));
  NAND3_X1  g672(.A1(new_n865), .A2(new_n255), .A3(new_n867), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(G183gat), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n482), .A3(new_n599), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n876), .B2(new_n256), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g677(.A1(new_n865), .A2(new_n326), .A3(new_n867), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(G190gat), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT61), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n880), .A2(KEYINPUT124), .A3(KEYINPUT61), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT125), .B1(new_n880), .B2(KEYINPUT61), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT125), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT61), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n879), .A2(new_n886), .A3(new_n887), .A4(G190gat), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n883), .A2(new_n884), .A3(new_n885), .A4(new_n888), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n860), .A2(new_n470), .A3(new_n599), .A4(new_n326), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(G1351gat));
  NOR2_X1   g690(.A1(new_n663), .A2(new_n600), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n859), .A2(new_n573), .A3(new_n892), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT126), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n529), .A3(new_n387), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n663), .A2(new_n648), .A3(new_n600), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n844), .A2(new_n393), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n895), .B1(new_n529), .B2(new_n897), .ZN(G1352gat));
  OR3_X1    g697(.A1(new_n893), .A2(G204gat), .A3(new_n671), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT127), .ZN(new_n900));
  OR3_X1    g699(.A1(new_n899), .A2(new_n900), .A3(KEYINPUT62), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(KEYINPUT62), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n844), .A2(new_n362), .A3(new_n896), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(G204gat), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n900), .B1(new_n899), .B2(KEYINPUT62), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n901), .A2(new_n902), .A3(new_n904), .A4(new_n905), .ZN(G1353gat));
  NAND3_X1  g705(.A1(new_n894), .A2(new_n242), .A3(new_n255), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n844), .A2(new_n255), .A3(new_n896), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n908), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT63), .B1(new_n908), .B2(G211gat), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(G1354gat));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n527), .A3(new_n326), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n844), .A2(new_n326), .A3(new_n896), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n527), .B2(new_n913), .ZN(G1355gat));
endmodule


