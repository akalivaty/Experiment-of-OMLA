

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U323 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U324 ( .A(n340), .B(n339), .ZN(n344) );
  XNOR2_X1 U325 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n428) );
  XNOR2_X1 U326 ( .A(n429), .B(n428), .ZN(n462) );
  NOR2_X1 U327 ( .A1(n538), .A2(n453), .ZN(n574) );
  XNOR2_X1 U328 ( .A(n455), .B(G176GAT), .ZN(n456) );
  XNOR2_X1 U329 ( .A(n457), .B(n456), .ZN(G1349GAT) );
  XOR2_X1 U330 ( .A(KEYINPUT84), .B(KEYINPUT86), .Z(n292) );
  NAND2_X1 U331 ( .A1(G227GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U332 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U333 ( .A(n293), .B(KEYINPUT20), .Z(n295) );
  XOR2_X1 U334 ( .A(G190GAT), .B(G134GAT), .Z(n393) );
  XOR2_X1 U335 ( .A(KEYINPUT0), .B(G127GAT), .Z(n441) );
  XNOR2_X1 U336 ( .A(n393), .B(n441), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n295), .B(n294), .ZN(n297) );
  XNOR2_X1 U338 ( .A(G99GAT), .B(G71GAT), .ZN(n296) );
  XNOR2_X1 U339 ( .A(n296), .B(G120GAT), .ZN(n342) );
  XOR2_X1 U340 ( .A(n297), .B(n342), .Z(n305) );
  XOR2_X1 U341 ( .A(G15GAT), .B(G113GAT), .Z(n299) );
  XNOR2_X1 U342 ( .A(G169GAT), .B(G43GAT), .ZN(n298) );
  XNOR2_X1 U343 ( .A(n299), .B(n298), .ZN(n349) );
  XNOR2_X1 U344 ( .A(G183GAT), .B(KEYINPUT19), .ZN(n300) );
  XNOR2_X1 U345 ( .A(n300), .B(G176GAT), .ZN(n301) );
  XOR2_X1 U346 ( .A(n301), .B(KEYINPUT85), .Z(n303) );
  XNOR2_X1 U347 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n303), .B(n302), .ZN(n416) );
  XNOR2_X1 U349 ( .A(n349), .B(n416), .ZN(n304) );
  XNOR2_X1 U350 ( .A(n305), .B(n304), .ZN(n538) );
  XNOR2_X1 U351 ( .A(G211GAT), .B(G218GAT), .ZN(n306) );
  XNOR2_X1 U352 ( .A(n306), .B(KEYINPUT89), .ZN(n307) );
  XOR2_X1 U353 ( .A(n307), .B(KEYINPUT21), .Z(n309) );
  XNOR2_X1 U354 ( .A(G197GAT), .B(G204GAT), .ZN(n308) );
  XNOR2_X1 U355 ( .A(n309), .B(n308), .ZN(n415) );
  XOR2_X1 U356 ( .A(G141GAT), .B(G22GAT), .Z(n346) );
  XOR2_X1 U357 ( .A(KEYINPUT24), .B(KEYINPUT91), .Z(n311) );
  XNOR2_X1 U358 ( .A(G50GAT), .B(KEYINPUT22), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U360 ( .A(n346), .B(n312), .Z(n314) );
  NAND2_X1 U361 ( .A1(G228GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U363 ( .A(n315), .B(KEYINPUT23), .Z(n318) );
  XNOR2_X1 U364 ( .A(G106GAT), .B(G78GAT), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n316), .B(G148GAT), .ZN(n327) );
  XNOR2_X1 U366 ( .A(n327), .B(KEYINPUT88), .ZN(n317) );
  XNOR2_X1 U367 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n415), .B(n319), .ZN(n323) );
  XOR2_X1 U369 ( .A(KEYINPUT3), .B(G162GAT), .Z(n321) );
  XNOR2_X1 U370 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U372 ( .A(KEYINPUT90), .B(n322), .ZN(n449) );
  XNOR2_X1 U373 ( .A(n323), .B(n449), .ZN(n475) );
  XOR2_X1 U374 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n364) );
  XOR2_X1 U375 ( .A(KEYINPUT74), .B(KEYINPUT76), .Z(n325) );
  XOR2_X1 U376 ( .A(G92GAT), .B(G64GAT), .Z(n417) );
  XOR2_X1 U377 ( .A(KEYINPUT73), .B(G85GAT), .Z(n392) );
  XNOR2_X1 U378 ( .A(n417), .B(n392), .ZN(n324) );
  XOR2_X1 U379 ( .A(n325), .B(n324), .Z(n334) );
  INV_X1 U380 ( .A(n327), .ZN(n326) );
  NAND2_X1 U381 ( .A1(n326), .A2(KEYINPUT31), .ZN(n330) );
  INV_X1 U382 ( .A(KEYINPUT31), .ZN(n328) );
  NAND2_X1 U383 ( .A1(n328), .A2(n327), .ZN(n329) );
  NAND2_X1 U384 ( .A1(n330), .A2(n329), .ZN(n332) );
  NAND2_X1 U385 ( .A1(G230GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U386 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U387 ( .A(n334), .B(n333), .ZN(n340) );
  XOR2_X1 U388 ( .A(KEYINPUT32), .B(KEYINPUT72), .Z(n336) );
  XNOR2_X1 U389 ( .A(KEYINPUT33), .B(KEYINPUT75), .ZN(n335) );
  XOR2_X1 U390 ( .A(n336), .B(n335), .Z(n338) );
  XNOR2_X1 U391 ( .A(G176GAT), .B(G204GAT), .ZN(n337) );
  XNOR2_X1 U392 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n341) );
  XNOR2_X1 U393 ( .A(n341), .B(KEYINPUT13), .ZN(n376) );
  XNOR2_X1 U394 ( .A(n342), .B(n376), .ZN(n343) );
  XNOR2_X1 U395 ( .A(n344), .B(n343), .ZN(n468) );
  XNOR2_X1 U396 ( .A(KEYINPUT41), .B(n468), .ZN(n454) );
  XNOR2_X1 U397 ( .A(G8GAT), .B(G1GAT), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n345), .B(KEYINPUT68), .ZN(n365) );
  XOR2_X1 U399 ( .A(KEYINPUT69), .B(n365), .Z(n348) );
  XNOR2_X1 U400 ( .A(n346), .B(G197GAT), .ZN(n347) );
  XNOR2_X1 U401 ( .A(n348), .B(n347), .ZN(n353) );
  XOR2_X1 U402 ( .A(n349), .B(KEYINPUT30), .Z(n351) );
  NAND2_X1 U403 ( .A1(G229GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U404 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U405 ( .A(n353), .B(n352), .Z(n362) );
  XNOR2_X1 U406 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n354) );
  XNOR2_X1 U407 ( .A(n354), .B(G29GAT), .ZN(n355) );
  XOR2_X1 U408 ( .A(n355), .B(KEYINPUT8), .Z(n357) );
  XNOR2_X1 U409 ( .A(G50GAT), .B(KEYINPUT67), .ZN(n356) );
  XNOR2_X1 U410 ( .A(n357), .B(n356), .ZN(n402) );
  XOR2_X1 U411 ( .A(KEYINPUT29), .B(KEYINPUT64), .Z(n359) );
  XNOR2_X1 U412 ( .A(KEYINPUT66), .B(KEYINPUT65), .ZN(n358) );
  XNOR2_X1 U413 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U414 ( .A(n402), .B(n360), .ZN(n361) );
  XNOR2_X1 U415 ( .A(n362), .B(n361), .ZN(n554) );
  NOR2_X1 U416 ( .A1(n454), .A2(n554), .ZN(n363) );
  XNOR2_X1 U417 ( .A(n364), .B(n363), .ZN(n386) );
  XOR2_X1 U418 ( .A(KEYINPUT80), .B(n365), .Z(n367) );
  NAND2_X1 U419 ( .A1(G231GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U420 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U421 ( .A(KEYINPUT82), .B(KEYINPUT12), .Z(n369) );
  XNOR2_X1 U422 ( .A(G64GAT), .B(KEYINPUT81), .ZN(n368) );
  XNOR2_X1 U423 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U424 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U425 ( .A(G71GAT), .B(G127GAT), .Z(n373) );
  XNOR2_X1 U426 ( .A(G15GAT), .B(G183GAT), .ZN(n372) );
  XNOR2_X1 U427 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U428 ( .A(n375), .B(n374), .ZN(n380) );
  XOR2_X1 U429 ( .A(n376), .B(G78GAT), .Z(n378) );
  XNOR2_X1 U430 ( .A(G22GAT), .B(G155GAT), .ZN(n377) );
  XNOR2_X1 U431 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U432 ( .A(n380), .B(n379), .Z(n385) );
  XOR2_X1 U433 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n382) );
  XNOR2_X1 U434 ( .A(KEYINPUT14), .B(KEYINPUT15), .ZN(n381) );
  XNOR2_X1 U435 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U436 ( .A(G211GAT), .B(n383), .ZN(n384) );
  XNOR2_X1 U437 ( .A(n385), .B(n384), .ZN(n581) );
  NOR2_X1 U438 ( .A1(n386), .A2(n581), .ZN(n387) );
  XNOR2_X1 U439 ( .A(n387), .B(KEYINPUT112), .ZN(n405) );
  XOR2_X1 U440 ( .A(KEYINPUT77), .B(KEYINPUT11), .Z(n389) );
  XNOR2_X1 U441 ( .A(G43GAT), .B(G162GAT), .ZN(n388) );
  XNOR2_X1 U442 ( .A(n389), .B(n388), .ZN(n401) );
  XOR2_X1 U443 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n391) );
  XNOR2_X1 U444 ( .A(G99GAT), .B(G106GAT), .ZN(n390) );
  XNOR2_X1 U445 ( .A(n391), .B(n390), .ZN(n397) );
  XOR2_X1 U446 ( .A(n392), .B(G92GAT), .Z(n395) );
  XNOR2_X1 U447 ( .A(n393), .B(G218GAT), .ZN(n394) );
  XNOR2_X1 U448 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U449 ( .A(n397), .B(n396), .Z(n399) );
  NAND2_X1 U450 ( .A1(G232GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U451 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U452 ( .A(n401), .B(n400), .ZN(n404) );
  INV_X1 U453 ( .A(n402), .ZN(n403) );
  XOR2_X1 U454 ( .A(n404), .B(n403), .Z(n575) );
  INV_X1 U455 ( .A(n575), .ZN(n567) );
  NAND2_X1 U456 ( .A1(n405), .A2(n567), .ZN(n406) );
  XNOR2_X1 U457 ( .A(n406), .B(KEYINPUT113), .ZN(n407) );
  XNOR2_X1 U458 ( .A(n407), .B(KEYINPUT47), .ZN(n413) );
  INV_X1 U459 ( .A(n581), .ZN(n563) );
  XNOR2_X1 U460 ( .A(KEYINPUT36), .B(KEYINPUT104), .ZN(n408) );
  XNOR2_X1 U461 ( .A(n408), .B(n567), .ZN(n585) );
  NOR2_X1 U462 ( .A1(n563), .A2(n585), .ZN(n409) );
  XOR2_X1 U463 ( .A(KEYINPUT45), .B(n409), .Z(n410) );
  NOR2_X1 U464 ( .A1(n468), .A2(n410), .ZN(n411) );
  XOR2_X1 U465 ( .A(n554), .B(KEYINPUT70), .Z(n569) );
  INV_X1 U466 ( .A(n569), .ZN(n469) );
  NAND2_X1 U467 ( .A1(n411), .A2(n469), .ZN(n412) );
  NAND2_X1 U468 ( .A1(n413), .A2(n412), .ZN(n414) );
  XNOR2_X1 U469 ( .A(n414), .B(KEYINPUT48), .ZN(n537) );
  XNOR2_X1 U470 ( .A(n416), .B(n415), .ZN(n427) );
  XOR2_X1 U471 ( .A(G8GAT), .B(n417), .Z(n419) );
  NAND2_X1 U472 ( .A1(G226GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U473 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U474 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n421) );
  XNOR2_X1 U475 ( .A(G169GAT), .B(KEYINPUT95), .ZN(n420) );
  XNOR2_X1 U476 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U477 ( .A(n423), .B(n422), .Z(n425) );
  XNOR2_X1 U478 ( .A(G36GAT), .B(G190GAT), .ZN(n424) );
  XNOR2_X1 U479 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U480 ( .A(n427), .B(n426), .ZN(n505) );
  NAND2_X1 U481 ( .A1(n537), .A2(n505), .ZN(n429) );
  XOR2_X1 U482 ( .A(G120GAT), .B(G1GAT), .Z(n431) );
  XNOR2_X1 U483 ( .A(G113GAT), .B(G141GAT), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U485 ( .A(KEYINPUT94), .B(KEYINPUT4), .Z(n433) );
  XNOR2_X1 U486 ( .A(G57GAT), .B(KEYINPUT5), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U488 ( .A(n435), .B(n434), .Z(n447) );
  XOR2_X1 U489 ( .A(KEYINPUT1), .B(KEYINPUT93), .Z(n437) );
  XNOR2_X1 U490 ( .A(KEYINPUT6), .B(KEYINPUT92), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n445) );
  XOR2_X1 U492 ( .A(G85GAT), .B(G148GAT), .Z(n439) );
  XNOR2_X1 U493 ( .A(G29GAT), .B(G134GAT), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U495 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U496 ( .A1(G225GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n449), .B(n448), .ZN(n525) );
  NAND2_X1 U501 ( .A1(n462), .A2(n525), .ZN(n450) );
  NOR2_X1 U502 ( .A1(n475), .A2(n450), .ZN(n452) );
  XNOR2_X1 U503 ( .A(KEYINPUT55), .B(KEYINPUT122), .ZN(n451) );
  XNOR2_X1 U504 ( .A(n452), .B(n451), .ZN(n453) );
  INV_X1 U505 ( .A(n454), .ZN(n543) );
  NAND2_X1 U506 ( .A1(n574), .A2(n543), .ZN(n457) );
  XOR2_X1 U507 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n455) );
  NAND2_X1 U508 ( .A1(n475), .A2(n538), .ZN(n458) );
  XNOR2_X1 U509 ( .A(n458), .B(KEYINPUT26), .ZN(n459) );
  XNOR2_X1 U510 ( .A(KEYINPUT98), .B(n459), .ZN(n552) );
  INV_X1 U511 ( .A(n552), .ZN(n460) );
  AND2_X1 U512 ( .A1(n525), .A2(n460), .ZN(n461) );
  AND2_X1 U513 ( .A1(n462), .A2(n461), .ZN(n582) );
  INV_X1 U514 ( .A(n582), .ZN(n584) );
  NOR2_X1 U515 ( .A1(n554), .A2(n584), .ZN(n464) );
  XNOR2_X1 U516 ( .A(KEYINPUT60), .B(KEYINPUT126), .ZN(n463) );
  XNOR2_X1 U517 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U518 ( .A(n465), .B(KEYINPUT59), .ZN(n467) );
  XOR2_X1 U519 ( .A(G197GAT), .B(KEYINPUT125), .Z(n466) );
  XNOR2_X1 U520 ( .A(n467), .B(n466), .ZN(G1352GAT) );
  NOR2_X1 U521 ( .A1(n468), .A2(n469), .ZN(n500) );
  INV_X1 U522 ( .A(n525), .ZN(n502) );
  INV_X1 U523 ( .A(n505), .ZN(n528) );
  NOR2_X1 U524 ( .A1(n538), .A2(n528), .ZN(n470) );
  NOR2_X1 U525 ( .A1(n475), .A2(n470), .ZN(n471) );
  XOR2_X1 U526 ( .A(KEYINPUT25), .B(n471), .Z(n473) );
  XOR2_X1 U527 ( .A(n505), .B(KEYINPUT27), .Z(n476) );
  NOR2_X1 U528 ( .A1(n476), .A2(n552), .ZN(n472) );
  NOR2_X1 U529 ( .A1(n473), .A2(n472), .ZN(n474) );
  NOR2_X1 U530 ( .A1(n502), .A2(n474), .ZN(n480) );
  XNOR2_X1 U531 ( .A(KEYINPUT28), .B(n475), .ZN(n541) );
  NOR2_X1 U532 ( .A1(n525), .A2(n476), .ZN(n536) );
  XOR2_X1 U533 ( .A(n538), .B(KEYINPUT87), .Z(n477) );
  NAND2_X1 U534 ( .A1(n536), .A2(n477), .ZN(n478) );
  NOR2_X1 U535 ( .A1(n541), .A2(n478), .ZN(n479) );
  NOR2_X1 U536 ( .A1(n480), .A2(n479), .ZN(n496) );
  XOR2_X1 U537 ( .A(KEYINPUT83), .B(KEYINPUT16), .Z(n482) );
  NAND2_X1 U538 ( .A1(n581), .A2(n567), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(n483) );
  NOR2_X1 U540 ( .A1(n496), .A2(n483), .ZN(n484) );
  XOR2_X1 U541 ( .A(KEYINPUT99), .B(n484), .Z(n512) );
  NAND2_X1 U542 ( .A1(n500), .A2(n512), .ZN(n485) );
  XNOR2_X1 U543 ( .A(n485), .B(KEYINPUT100), .ZN(n492) );
  NOR2_X1 U544 ( .A1(n525), .A2(n492), .ZN(n486) );
  XOR2_X1 U545 ( .A(KEYINPUT34), .B(n486), .Z(n487) );
  XNOR2_X1 U546 ( .A(G1GAT), .B(n487), .ZN(G1324GAT) );
  NOR2_X1 U547 ( .A1(n492), .A2(n528), .ZN(n489) );
  XNOR2_X1 U548 ( .A(G8GAT), .B(KEYINPUT101), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(G1325GAT) );
  XNOR2_X1 U550 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n491) );
  NOR2_X1 U551 ( .A1(n538), .A2(n492), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n491), .B(n490), .ZN(G1326GAT) );
  INV_X1 U553 ( .A(n541), .ZN(n533) );
  NOR2_X1 U554 ( .A1(n492), .A2(n533), .ZN(n494) );
  XNOR2_X1 U555 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U557 ( .A(G22GAT), .B(n495), .ZN(G1327GAT) );
  XOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT39), .Z(n504) );
  XOR2_X1 U559 ( .A(KEYINPUT37), .B(KEYINPUT105), .Z(n499) );
  NOR2_X1 U560 ( .A1(n496), .A2(n585), .ZN(n497) );
  NAND2_X1 U561 ( .A1(n497), .A2(n563), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n499), .B(n498), .ZN(n524) );
  NAND2_X1 U563 ( .A1(n524), .A2(n500), .ZN(n501) );
  XOR2_X1 U564 ( .A(KEYINPUT38), .B(n501), .Z(n510) );
  NAND2_X1 U565 ( .A1(n510), .A2(n502), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n504), .B(n503), .ZN(G1328GAT) );
  NAND2_X1 U567 ( .A1(n510), .A2(n505), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n506), .B(G36GAT), .ZN(G1329GAT) );
  INV_X1 U569 ( .A(n538), .ZN(n507) );
  NAND2_X1 U570 ( .A1(n507), .A2(n510), .ZN(n508) );
  XNOR2_X1 U571 ( .A(KEYINPUT40), .B(n508), .ZN(n509) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(n509), .ZN(G1330GAT) );
  NAND2_X1 U573 ( .A1(n510), .A2(n541), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n511), .B(G50GAT), .ZN(G1331GAT) );
  AND2_X1 U575 ( .A1(n554), .A2(n543), .ZN(n523) );
  NAND2_X1 U576 ( .A1(n512), .A2(n523), .ZN(n519) );
  NOR2_X1 U577 ( .A1(n525), .A2(n519), .ZN(n513) );
  XOR2_X1 U578 ( .A(G57GAT), .B(n513), .Z(n514) );
  XNOR2_X1 U579 ( .A(KEYINPUT42), .B(n514), .ZN(G1332GAT) );
  NOR2_X1 U580 ( .A1(n528), .A2(n519), .ZN(n515) );
  XOR2_X1 U581 ( .A(G64GAT), .B(n515), .Z(G1333GAT) );
  NOR2_X1 U582 ( .A1(n538), .A2(n519), .ZN(n517) );
  XNOR2_X1 U583 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U585 ( .A(G71GAT), .B(n518), .ZN(G1334GAT) );
  NOR2_X1 U586 ( .A1(n533), .A2(n519), .ZN(n521) );
  XNOR2_X1 U587 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U589 ( .A(G78GAT), .B(n522), .ZN(G1335GAT) );
  NAND2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n532) );
  NOR2_X1 U591 ( .A1(n525), .A2(n532), .ZN(n527) );
  XNOR2_X1 U592 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(G1336GAT) );
  NOR2_X1 U594 ( .A1(n528), .A2(n532), .ZN(n529) );
  XOR2_X1 U595 ( .A(KEYINPUT110), .B(n529), .Z(n530) );
  XNOR2_X1 U596 ( .A(G92GAT), .B(n530), .ZN(G1337GAT) );
  NOR2_X1 U597 ( .A1(n538), .A2(n532), .ZN(n531) );
  XOR2_X1 U598 ( .A(G99GAT), .B(n531), .Z(G1338GAT) );
  NOR2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U600 ( .A(KEYINPUT44), .B(n534), .Z(n535) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(n535), .ZN(G1339GAT) );
  NAND2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n553) );
  NOR2_X1 U603 ( .A1(n538), .A2(n553), .ZN(n539) );
  XOR2_X1 U604 ( .A(KEYINPUT114), .B(n539), .Z(n540) );
  NOR2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n549), .A2(n569), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n542), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n545) );
  NAND2_X1 U609 ( .A1(n549), .A2(n543), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U611 ( .A(G120GAT), .B(n546), .Z(G1341GAT) );
  NAND2_X1 U612 ( .A1(n549), .A2(n581), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n547), .B(KEYINPUT50), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G127GAT), .B(n548), .ZN(G1342GAT) );
  XOR2_X1 U615 ( .A(G134GAT), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U616 ( .A1(n549), .A2(n575), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1343GAT) );
  OR2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n566) );
  NOR2_X1 U619 ( .A1(n554), .A2(n566), .ZN(n555) );
  XOR2_X1 U620 ( .A(n555), .B(KEYINPUT116), .Z(n556) );
  XNOR2_X1 U621 ( .A(G141GAT), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT119), .B(KEYINPUT118), .Z(n558) );
  XNOR2_X1 U623 ( .A(KEYINPUT117), .B(KEYINPUT53), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(n562) );
  NOR2_X1 U625 ( .A1(n454), .A2(n566), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U628 ( .A(n562), .B(n561), .Z(G1345GAT) );
  NOR2_X1 U629 ( .A1(n563), .A2(n566), .ZN(n564) );
  XOR2_X1 U630 ( .A(KEYINPUT120), .B(n564), .Z(n565) );
  XNOR2_X1 U631 ( .A(G155GAT), .B(n565), .ZN(G1346GAT) );
  NOR2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U633 ( .A(G162GAT), .B(n568), .Z(G1347GAT) );
  XOR2_X1 U634 ( .A(G169GAT), .B(KEYINPUT123), .Z(n571) );
  NAND2_X1 U635 ( .A1(n574), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1348GAT) );
  NAND2_X1 U637 ( .A1(n574), .A2(n581), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(KEYINPUT124), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U640 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1351GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n579) );
  NAND2_X1 U644 ( .A1(n582), .A2(n468), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XOR2_X1 U646 ( .A(G204GAT), .B(n580), .Z(G1353GAT) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(n586), .Z(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

