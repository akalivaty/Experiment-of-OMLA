//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT3), .ZN(new_n188));
  OR2_X1    g002(.A1(KEYINPUT77), .A2(G107), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT77), .A2(G107), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n189), .A3(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT78), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G104), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n187), .A2(KEYINPUT78), .A3(G107), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G101), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n193), .A2(G104), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT3), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n191), .A2(new_n196), .A3(new_n197), .A4(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(G104), .B1(new_n189), .B2(new_n190), .ZN(new_n201));
  INV_X1    g015(.A(new_n198), .ZN(new_n202));
  OAI21_X1  g016(.A(G101), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G119), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G116), .ZN(new_n207));
  INV_X1    g021(.A(G116), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G119), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT2), .B(G113), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT66), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G113), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT2), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT2), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G113), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G116), .B(G119), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n212), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT81), .B(KEYINPUT5), .ZN(new_n222));
  INV_X1    g036(.A(new_n207), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n213), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n224), .B1(new_n210), .B2(new_n222), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n205), .A2(new_n221), .A3(new_n225), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n187), .A2(KEYINPUT78), .A3(G107), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT78), .B1(new_n187), .B2(G107), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n199), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n188), .A2(new_n189), .A3(new_n190), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT79), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT79), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n191), .A2(new_n196), .A3(new_n232), .A4(new_n199), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n197), .A2(KEYINPUT4), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n217), .A2(new_n218), .ZN(new_n236));
  AOI211_X1 g050(.A(KEYINPUT67), .B(new_n236), .C1(new_n220), .C2(new_n212), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n210), .A2(new_n211), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n238), .B1(new_n221), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n235), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n231), .A2(G101), .A3(new_n233), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n200), .A2(KEYINPUT4), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n226), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(G110), .B(G122), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n226), .B(new_n246), .C1(new_n241), .C2(new_n244), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(KEYINPUT6), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT6), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n245), .A2(new_n251), .A3(new_n247), .ZN(new_n252));
  INV_X1    g066(.A(G143), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(G146), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n255));
  INV_X1    g069(.A(G146), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(G143), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n253), .A2(KEYINPUT64), .A3(G146), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n254), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G128), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(KEYINPUT1), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT1), .ZN(new_n263));
  OAI21_X1  g077(.A(G128), .B1(new_n254), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n256), .A2(G143), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n253), .A2(G146), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(G125), .ZN(new_n270));
  NAND2_X1  g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(KEYINPUT0), .A2(G128), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n259), .A2(new_n272), .B1(new_n274), .B2(new_n267), .ZN(new_n275));
  INV_X1    g089(.A(G125), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n270), .A2(new_n277), .ZN(new_n278));
  XOR2_X1   g092(.A(KEYINPUT82), .B(G224), .Z(new_n279));
  NOR2_X1   g093(.A1(new_n279), .A2(G953), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n278), .B(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n250), .A2(new_n252), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n278), .B1(KEYINPUT7), .B2(new_n281), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n204), .A2(new_n221), .A3(new_n225), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n246), .B(KEYINPUT8), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT5), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n224), .B1(new_n288), .B2(new_n210), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n204), .B1(new_n221), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT7), .ZN(new_n292));
  NOR4_X1   g106(.A1(new_n270), .A2(new_n277), .A3(new_n292), .A4(new_n280), .ZN(new_n293));
  NOR3_X1   g107(.A1(new_n284), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(G902), .B1(new_n294), .B2(new_n249), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n283), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(G210), .B1(G237), .B2(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n283), .A2(new_n295), .A3(new_n297), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(KEYINPUT83), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(G214), .B1(G237), .B2(G902), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT83), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n296), .A2(new_n303), .A3(new_n298), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n301), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT84), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT84), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n301), .A2(new_n307), .A3(new_n302), .A4(new_n304), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  XOR2_X1   g123(.A(KEYINPUT70), .B(G902), .Z(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT28), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n257), .A2(new_n258), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(new_n272), .A3(new_n265), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n274), .A2(new_n267), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT65), .ZN(new_n317));
  INV_X1    g131(.A(G134), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n317), .B1(new_n318), .B2(G137), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT11), .ZN(new_n320));
  INV_X1    g134(.A(G131), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT11), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n317), .B(new_n322), .C1(new_n318), .C2(G137), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n318), .A2(G137), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n320), .A2(new_n321), .A3(new_n323), .A4(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G137), .ZN(new_n326));
  AOI21_X1  g140(.A(KEYINPUT65), .B1(new_n326), .B2(G134), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n324), .B1(new_n327), .B2(new_n322), .ZN(new_n328));
  INV_X1    g142(.A(new_n323), .ZN(new_n329));
  OAI21_X1  g143(.A(G131), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n316), .B1(new_n325), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n318), .A2(G137), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n326), .A2(G134), .ZN(new_n333));
  OAI21_X1  g147(.A(G131), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n325), .A2(new_n334), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n259), .A2(new_n261), .B1(new_n264), .B2(new_n267), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI22_X1  g151(.A1(new_n331), .A2(new_n337), .B1(new_n237), .B2(new_n240), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n219), .B1(new_n217), .B2(new_n218), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n239), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT67), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n269), .A2(new_n325), .A3(new_n334), .ZN(new_n343));
  INV_X1    g157(.A(new_n325), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n333), .B1(new_n319), .B2(KEYINPUT11), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n321), .B1(new_n345), .B2(new_n323), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n275), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n221), .A2(new_n238), .A3(new_n239), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n342), .A2(new_n343), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n312), .B1(new_n338), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(G237), .A2(G953), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G210), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(KEYINPUT27), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT26), .B(G101), .ZN(new_n354));
  XOR2_X1   g168(.A(new_n353), .B(new_n354), .Z(new_n355));
  NOR2_X1   g169(.A1(new_n237), .A2(new_n240), .ZN(new_n356));
  INV_X1    g170(.A(new_n335), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n330), .A2(new_n325), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n357), .A2(new_n269), .B1(new_n358), .B2(new_n275), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT28), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n350), .A2(new_n355), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n311), .B1(new_n361), .B2(KEYINPUT29), .ZN(new_n362));
  AND4_X1   g176(.A1(new_n348), .A2(new_n342), .A3(new_n347), .A4(new_n343), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n348), .A2(new_n342), .B1(new_n343), .B2(new_n347), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT28), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n353), .B(new_n354), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n349), .A2(new_n312), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n365), .A2(KEYINPUT69), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT29), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT30), .B1(new_n331), .B2(new_n337), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT30), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n343), .A2(new_n347), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n356), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n355), .B1(new_n373), .B2(new_n363), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n368), .A2(new_n369), .A3(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n350), .A2(new_n360), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT69), .B1(new_n376), .B2(new_n366), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n362), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G472), .ZN(new_n379));
  NOR2_X1   g193(.A1(G472), .A2(G902), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n349), .A2(new_n366), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT68), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n370), .A2(new_n372), .ZN(new_n383));
  INV_X1    g197(.A(new_n356), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT31), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT68), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n349), .A2(new_n387), .A3(new_n366), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n382), .A2(new_n385), .A3(new_n386), .A4(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n355), .B1(new_n350), .B2(new_n360), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n355), .B1(new_n356), .B2(new_n359), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n387), .A2(new_n392), .B1(new_n383), .B2(new_n384), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n386), .B1(new_n393), .B2(new_n382), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n380), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT32), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g211(.A(KEYINPUT32), .B(new_n380), .C1(new_n391), .C2(new_n394), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n379), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT22), .B(G137), .ZN(new_n400));
  INV_X1    g214(.A(G953), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(G221), .A3(G234), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n400), .B(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G110), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT71), .ZN(new_n405));
  OAI211_X1 g219(.A(G119), .B(new_n260), .C1(new_n405), .C2(KEYINPUT23), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT23), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n407), .B1(new_n206), .B2(G128), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT71), .B1(new_n206), .B2(G128), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n406), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n404), .B1(new_n410), .B2(KEYINPUT72), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n411), .B1(KEYINPUT72), .B2(new_n410), .ZN(new_n412));
  XOR2_X1   g226(.A(G119), .B(G128), .Z(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT24), .B(G110), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G140), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G125), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n276), .A2(G140), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT73), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n276), .A2(G140), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT73), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n420), .A2(new_n422), .A3(KEYINPUT16), .ZN(new_n423));
  OR2_X1    g237(.A1(new_n421), .A2(KEYINPUT16), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n256), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n256), .B1(new_n423), .B2(new_n424), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n412), .B(new_n415), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n423), .A2(new_n424), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G146), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n413), .A2(new_n414), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n410), .B2(G110), .ZN(new_n432));
  XNOR2_X1  g246(.A(G125), .B(G140), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n256), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n430), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n428), .A2(KEYINPUT74), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT74), .B1(new_n428), .B2(new_n435), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n403), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n403), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n428), .A2(new_n435), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT74), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G217), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(new_n310), .B2(G234), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(G902), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n438), .A2(new_n310), .A3(new_n442), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT25), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n438), .A2(KEYINPUT25), .A3(new_n310), .A4(new_n442), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n448), .B1(new_n453), .B2(new_n445), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n399), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G113), .B(G122), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(new_n187), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n420), .A2(new_n422), .A3(G146), .ZN(new_n459));
  OR2_X1    g273(.A1(new_n459), .A2(KEYINPUT85), .ZN(new_n460));
  NAND2_X1  g274(.A1(KEYINPUT18), .A2(G131), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n351), .A2(G143), .A3(G214), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(G143), .B1(new_n351), .B2(G214), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G237), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n401), .A3(G214), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n253), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n468), .A2(KEYINPUT18), .A3(G131), .A4(new_n462), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n459), .A2(KEYINPUT85), .A3(new_n434), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n460), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n426), .A2(new_n427), .ZN(new_n473));
  OAI211_X1 g287(.A(KEYINPUT17), .B(G131), .C1(new_n463), .C2(new_n464), .ZN(new_n474));
  AOI21_X1  g288(.A(KEYINPUT87), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n430), .A2(KEYINPUT87), .A3(new_n425), .A4(new_n474), .ZN(new_n476));
  OAI21_X1  g290(.A(G131), .B1(new_n463), .B2(new_n464), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n468), .A2(new_n321), .A3(new_n462), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OR2_X1    g293(.A1(new_n479), .A2(KEYINPUT17), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n458), .B(new_n472), .C1(new_n475), .C2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT86), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT19), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n485), .B1(new_n420), .B2(new_n422), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n433), .A2(KEYINPUT19), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n256), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n430), .A2(new_n479), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n472), .ZN(new_n490));
  INV_X1    g304(.A(new_n458), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n484), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI211_X1 g306(.A(KEYINPUT86), .B(new_n458), .C1(new_n489), .C2(new_n472), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n483), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(G475), .A2(G902), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT89), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT20), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT89), .B1(G475), .B2(G902), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT88), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n503), .B1(new_n483), .B2(new_n494), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n482), .B(KEYINPUT88), .C1(new_n492), .C2(new_n493), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n496), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n502), .B1(new_n506), .B2(KEYINPUT20), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n472), .B1(new_n475), .B2(new_n481), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n491), .ZN(new_n509));
  AOI21_X1  g323(.A(G902), .B1(new_n509), .B2(new_n482), .ZN(new_n510));
  XOR2_X1   g324(.A(KEYINPUT90), .B(G475), .Z(new_n511));
  NOR2_X1   g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT93), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n208), .A2(G122), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT92), .B1(new_n514), .B2(KEYINPUT14), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n208), .A2(G122), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(KEYINPUT14), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NOR3_X1   g332(.A1(new_n514), .A2(KEYINPUT92), .A3(KEYINPUT14), .ZN(new_n519));
  OAI21_X1  g333(.A(G107), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n516), .A2(new_n514), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n189), .A2(new_n190), .ZN(new_n522));
  OR2_X1    g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  XOR2_X1   g337(.A(G128), .B(G143), .Z(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(G134), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n524), .A2(G134), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n520), .B(new_n523), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n521), .B(new_n522), .ZN(new_n528));
  OR3_X1    g342(.A1(new_n524), .A2(KEYINPUT91), .A3(G134), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT91), .B1(new_n524), .B2(G134), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT13), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(new_n253), .A3(G128), .ZN(new_n532));
  OAI211_X1 g346(.A(G134), .B(new_n532), .C1(new_n524), .C2(new_n531), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n528), .A2(new_n529), .A3(new_n530), .A4(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT9), .B(G234), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n535), .A2(new_n444), .A3(G953), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n527), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n536), .B1(new_n527), .B2(new_n534), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n513), .B1(new_n539), .B2(new_n311), .ZN(new_n540));
  INV_X1    g354(.A(G478), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n541), .A2(KEYINPUT15), .ZN(new_n542));
  OAI211_X1 g356(.A(KEYINPUT93), .B(new_n310), .C1(new_n537), .C2(new_n538), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  OAI221_X1 g358(.A(new_n310), .B1(KEYINPUT15), .B2(new_n541), .C1(new_n537), .C2(new_n538), .ZN(new_n545));
  INV_X1    g359(.A(G952), .ZN(new_n546));
  AOI211_X1 g360(.A(G953), .B(new_n546), .C1(G234), .C2(G237), .ZN(new_n547));
  AOI211_X1 g361(.A(new_n401), .B(new_n310), .C1(G234), .C2(G237), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT21), .B(G898), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n544), .A2(new_n545), .A3(new_n551), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n507), .A2(new_n512), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G469), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n242), .A2(new_n243), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(new_n275), .A3(new_n235), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n259), .A2(new_n261), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n260), .B1(new_n265), .B2(KEYINPUT1), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n259), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n200), .B(new_n203), .C1(new_n557), .C2(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT80), .B(KEYINPUT10), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT10), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n336), .A2(new_n562), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n560), .A2(new_n561), .B1(new_n205), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n344), .A2(new_n346), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n556), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n401), .A2(G227), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT76), .ZN(new_n568));
  XNOR2_X1  g382(.A(G110), .B(G140), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n568), .B(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n204), .A2(new_n336), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n565), .B1(new_n560), .B2(new_n572), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n573), .A2(KEYINPUT12), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(KEYINPUT12), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n566), .B(new_n571), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n556), .A2(new_n564), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n358), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n571), .B1(new_n579), .B2(new_n566), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n554), .B(new_n310), .C1(new_n577), .C2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n566), .B1(new_n574), .B2(new_n575), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n570), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n579), .A2(new_n571), .A3(new_n566), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(G469), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(G469), .A2(G902), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n581), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(G221), .B1(new_n535), .B2(G902), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n588), .B(KEYINPUT75), .Z(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n553), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n309), .A2(new_n456), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(G101), .ZN(G3));
  INV_X1    g408(.A(KEYINPUT95), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n299), .A2(new_n595), .A3(new_n300), .ZN(new_n596));
  INV_X1    g410(.A(new_n302), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n297), .B1(new_n283), .B2(new_n295), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n597), .B1(new_n598), .B2(KEYINPUT95), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n600), .A2(new_n550), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n507), .A2(new_n512), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n603));
  XOR2_X1   g417(.A(new_n539), .B(KEYINPUT33), .Z(new_n604));
  NAND3_X1  g418(.A1(new_n604), .A2(G478), .A3(new_n310), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n602), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT94), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n389), .A2(new_n390), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n382), .A2(new_n385), .A3(new_n388), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT31), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n311), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(G472), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n608), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n611), .A2(new_n390), .A3(new_n389), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n310), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(KEYINPUT94), .A3(G472), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n614), .A2(new_n395), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n454), .A2(new_n590), .A3(new_n587), .ZN(new_n619));
  OR2_X1    g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n607), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT96), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT34), .B(G104), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  XNOR2_X1  g438(.A(new_n506), .B(KEYINPUT20), .ZN(new_n625));
  INV_X1    g439(.A(new_n512), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n544), .A2(new_n545), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n601), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(new_n620), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT35), .B(G107), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  INV_X1    g446(.A(new_n618), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n453), .A2(new_n445), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n439), .A2(KEYINPUT36), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n440), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n446), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n309), .A2(new_n592), .A3(new_n633), .A4(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT37), .B(G110), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G12));
  AND3_X1   g455(.A1(new_n399), .A2(new_n591), .A3(new_n638), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n547), .B(KEYINPUT97), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(G900), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n644), .B1(new_n645), .B2(new_n548), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  AND4_X1   g461(.A1(new_n626), .A2(new_n625), .A3(new_n627), .A4(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n600), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n642), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G128), .ZN(G30));
  XOR2_X1   g465(.A(new_n646), .B(KEYINPUT39), .Z(new_n652));
  NAND2_X1  g466(.A1(new_n591), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT40), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n301), .A2(new_n304), .ZN(new_n655));
  XOR2_X1   g469(.A(new_n655), .B(KEYINPUT38), .Z(new_n656));
  NOR2_X1   g470(.A1(new_n638), .A2(new_n597), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n506), .A2(KEYINPUT20), .ZN(new_n658));
  INV_X1    g472(.A(new_n502), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n626), .ZN(new_n661));
  INV_X1    g475(.A(G902), .ZN(new_n662));
  INV_X1    g476(.A(new_n610), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n366), .B1(new_n338), .B2(new_n349), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(G472), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n397), .A2(new_n398), .A3(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n657), .A2(new_n661), .A3(new_n627), .A4(new_n667), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n656), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n654), .B1(new_n669), .B2(KEYINPUT98), .ZN(new_n670));
  OR3_X1    g484(.A1(new_n656), .A2(KEYINPUT98), .A3(new_n668), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT99), .B(G143), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G45));
  NAND4_X1  g488(.A1(new_n642), .A2(new_n606), .A3(new_n649), .A4(new_n647), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G146), .ZN(G48));
  NOR2_X1   g490(.A1(new_n577), .A2(new_n580), .ZN(new_n677));
  OAI21_X1  g491(.A(G469), .B1(new_n677), .B2(new_n311), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n678), .A2(new_n590), .A3(new_n581), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n399), .A2(new_n679), .A3(new_n454), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(new_n601), .A3(new_n606), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G15));
  NAND3_X1  g497(.A1(new_n680), .A2(new_n601), .A3(new_n628), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G116), .ZN(G18));
  INV_X1    g499(.A(new_n679), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n600), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n553), .A2(new_n399), .A3(new_n638), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G119), .ZN(G21));
  OAI21_X1  g504(.A(new_n627), .B1(new_n507), .B2(new_n512), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n600), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n616), .A2(G472), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n454), .A2(new_n693), .A3(new_n395), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n678), .A2(new_n551), .A3(new_n590), .A4(new_n581), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G122), .ZN(G24));
  NAND2_X1  g512(.A1(new_n605), .A2(new_n603), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n661), .A2(KEYINPUT100), .A3(new_n699), .A4(new_n647), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n638), .A2(new_n395), .A3(new_n693), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n699), .B(new_n647), .C1(new_n507), .C2(new_n512), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT100), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n687), .A2(new_n700), .A3(new_n702), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G125), .ZN(G27));
  INV_X1    g521(.A(KEYINPUT42), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n398), .A2(KEYINPUT102), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT102), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n615), .A2(new_n710), .A3(KEYINPUT32), .A4(new_n380), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n709), .A2(new_n379), .A3(new_n397), .A4(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n454), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT103), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT103), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n712), .A2(new_n715), .A3(new_n454), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n708), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n597), .B1(new_n301), .B2(new_n304), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n586), .B(KEYINPUT101), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n585), .A2(new_n719), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n556), .A2(new_n564), .A3(new_n565), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n565), .B1(new_n556), .B2(new_n564), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n570), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI211_X1 g537(.A(G469), .B(new_n311), .C1(new_n723), .C2(new_n576), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n590), .B1(new_n720), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  AND4_X1   g540(.A1(new_n705), .A2(new_n700), .A3(new_n718), .A4(new_n726), .ZN(new_n727));
  AOI211_X1 g541(.A(new_n597), .B(new_n725), .C1(new_n301), .C2(new_n304), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(new_n456), .A3(new_n705), .A4(new_n700), .ZN(new_n729));
  AOI22_X1  g543(.A1(new_n717), .A2(new_n727), .B1(new_n729), .B2(new_n708), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n321), .ZN(G33));
  NAND3_X1  g545(.A1(new_n728), .A2(new_n648), .A3(new_n456), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G134), .ZN(G36));
  AND2_X1   g547(.A1(new_n618), .A2(new_n638), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n602), .A2(new_n699), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT105), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT43), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n583), .A2(new_n584), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n743), .A2(KEYINPUT45), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(KEYINPUT45), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(G469), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n719), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT104), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n747), .A2(KEYINPUT104), .A3(new_n748), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n746), .A2(KEYINPUT46), .A3(new_n719), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n751), .A2(new_n581), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n590), .A3(new_n652), .ZN(new_n755));
  INV_X1    g569(.A(new_n718), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n736), .A2(KEYINPUT44), .A3(new_n739), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n742), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G137), .ZN(G39));
  INV_X1    g574(.A(KEYINPUT47), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(KEYINPUT107), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(KEYINPUT107), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n754), .B(new_n590), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  NOR4_X1   g579(.A1(new_n756), .A2(new_n454), .A3(new_n399), .A4(new_n703), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n754), .A2(new_n590), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n765), .B(new_n766), .C1(new_n767), .C2(new_n764), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G140), .ZN(G42));
  XNOR2_X1  g583(.A(new_n655), .B(KEYINPUT38), .ZN(new_n770));
  INV_X1    g584(.A(new_n454), .ZN(new_n771));
  OR4_X1    g585(.A1(new_n771), .A2(new_n737), .A3(new_n597), .A4(new_n589), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n678), .A2(new_n581), .ZN(new_n773));
  AOI22_X1  g587(.A1(new_n772), .A2(KEYINPUT108), .B1(KEYINPUT49), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n774), .B1(KEYINPUT108), .B2(new_n772), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(KEYINPUT109), .Z(new_n776));
  NOR2_X1   g590(.A1(new_n773), .A2(KEYINPUT49), .ZN(new_n777));
  OR4_X1    g591(.A1(new_n770), .A2(new_n776), .A3(new_n667), .A4(new_n777), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n739), .A2(new_n644), .ZN(new_n779));
  INV_X1    g593(.A(new_n694), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n770), .A2(new_n302), .A3(new_n686), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(KEYINPUT50), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n785));
  INV_X1    g599(.A(new_n783), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n785), .B1(new_n781), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n756), .A2(new_n686), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n779), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n547), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n771), .A2(new_n667), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n602), .A2(new_n603), .A3(new_n605), .ZN(new_n794));
  OAI221_X1 g608(.A(new_n788), .B1(new_n701), .B2(new_n790), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n765), .B1(new_n767), .B2(new_n764), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n678), .A2(new_n589), .A3(new_n581), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(KEYINPUT113), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(new_n718), .A3(new_n782), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT113), .B1(new_n796), .B2(new_n797), .ZN(new_n800));
  OAI21_X1  g614(.A(KEYINPUT51), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n795), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n803));
  AOI211_X1 g617(.A(new_n756), .B(new_n781), .C1(new_n796), .C2(new_n797), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n803), .B1(new_n795), .B2(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n714), .A2(new_n716), .ZN(new_n806));
  NOR2_X1   g620(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n807));
  AND2_X1   g621(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n808));
  OR4_X1    g622(.A1(new_n806), .A2(new_n790), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n807), .B1(new_n790), .B2(new_n806), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n789), .A2(new_n606), .A3(new_n792), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(G952), .A3(new_n401), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n812), .B1(new_n782), .B2(new_n687), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n809), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n802), .A2(new_n805), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n618), .A2(new_n619), .A3(new_n550), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n309), .A2(new_n606), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n593), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT110), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n602), .A2(new_n627), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n309), .A2(new_n817), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n639), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n819), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n687), .A2(new_n688), .B1(new_n692), .B2(new_n696), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n680), .B(new_n601), .C1(new_n606), .C2(new_n628), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n627), .A2(new_n646), .ZN(new_n827));
  INV_X1    g641(.A(new_n658), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n506), .A2(KEYINPUT20), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n626), .B(new_n827), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT111), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n625), .A2(KEYINPUT111), .A3(new_n626), .A4(new_n827), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n642), .A2(new_n832), .A3(new_n718), .A4(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n825), .A2(new_n732), .A3(new_n826), .A4(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n730), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n639), .A2(KEYINPUT110), .A3(new_n822), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n727), .A2(KEYINPUT112), .A3(new_n702), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT112), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n728), .A2(new_n705), .A3(new_n700), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n839), .B1(new_n840), .B2(new_n701), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n824), .A2(new_n836), .A3(new_n837), .A4(new_n842), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n638), .A2(new_n646), .A3(new_n725), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n692), .A2(new_n667), .A3(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n706), .A2(new_n675), .A3(new_n650), .A4(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT52), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n816), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n838), .A2(new_n841), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n849), .A2(new_n730), .A3(new_n835), .ZN(new_n850));
  INV_X1    g664(.A(new_n837), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT110), .B1(new_n639), .B2(new_n822), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n851), .A2(new_n852), .A3(new_n819), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT52), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n846), .B(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n850), .A2(new_n853), .A3(new_n855), .A4(KEYINPUT53), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n848), .A2(KEYINPUT54), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT54), .B1(new_n848), .B2(new_n856), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n815), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(G952), .A2(G953), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n778), .B1(new_n860), .B2(new_n861), .ZN(G75));
  NAND2_X1  g676(.A1(new_n546), .A2(G953), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT116), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n848), .A2(new_n856), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n311), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT56), .B1(new_n867), .B2(new_n298), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n250), .A2(new_n252), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(new_n282), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT55), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n864), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n868), .A2(new_n871), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT115), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n868), .A2(KEYINPUT115), .A3(new_n871), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n872), .B1(new_n875), .B2(new_n876), .ZN(G51));
  XNOR2_X1  g691(.A(new_n719), .B(KEYINPUT117), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(KEYINPUT57), .Z(new_n879));
  AOI21_X1  g693(.A(new_n677), .B1(new_n859), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n746), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n865), .A2(new_n311), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT118), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n865), .A2(new_n884), .A3(new_n311), .A4(new_n881), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n864), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI211_X1 g703(.A(KEYINPUT119), .B(new_n864), .C1(new_n880), .C2(new_n886), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(G54));
  NAND3_X1  g705(.A1(new_n867), .A2(KEYINPUT58), .A3(G475), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n504), .A2(new_n505), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n892), .A2(new_n894), .ZN(new_n896));
  INV_X1    g710(.A(new_n864), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G60));
  XNOR2_X1  g712(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n541), .A2(new_n662), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n899), .B(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n859), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n604), .B(KEYINPUT120), .Z(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n864), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n902), .B2(new_n904), .ZN(G63));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n864), .B1(new_n907), .B2(KEYINPUT61), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n848), .A2(new_n856), .ZN(new_n909));
  NAND2_X1  g723(.A1(G217), .A2(G902), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT60), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n908), .B1(new_n912), .B2(new_n636), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n443), .B1(new_n909), .B2(new_n911), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n907), .A2(KEYINPUT61), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n915), .B(new_n916), .ZN(G66));
  NOR2_X1   g731(.A1(new_n279), .A2(new_n549), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(new_n401), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n825), .A2(new_n826), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n853), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n919), .B1(new_n922), .B2(new_n401), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n869), .B1(G898), .B2(new_n401), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n923), .B(new_n924), .Z(G69));
  NOR2_X1   g739(.A1(new_n486), .A2(new_n487), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT123), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n383), .B(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n401), .A2(G900), .ZN(new_n929));
  NOR4_X1   g743(.A1(new_n755), .A2(new_n600), .A3(new_n691), .A4(new_n806), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n706), .A2(new_n675), .A3(new_n650), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n732), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n930), .A2(new_n730), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n934), .A2(new_n759), .A3(new_n768), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n929), .B1(new_n935), .B2(new_n401), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(KEYINPUT125), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT125), .ZN(new_n938));
  AOI211_X1 g752(.A(new_n938), .B(new_n929), .C1(new_n935), .C2(new_n401), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n928), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n931), .B1(new_n670), .B2(new_n671), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n756), .A2(new_n455), .A3(new_n653), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n606), .B2(new_n821), .ZN(new_n945));
  AND4_X1   g759(.A1(new_n759), .A2(new_n943), .A3(new_n768), .A4(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n941), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT124), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT62), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT124), .B1(new_n941), .B2(new_n942), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n946), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n928), .A2(G953), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT126), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n928), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n401), .B1(G227), .B2(G900), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n940), .A2(new_n954), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n958), .B1(new_n940), .B2(new_n954), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(G72));
  NAND2_X1  g775(.A1(G472), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT63), .Z(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(new_n935), .B2(new_n922), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT127), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n373), .A2(new_n363), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n965), .A2(new_n355), .A3(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n922), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n946), .A2(new_n951), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n963), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n966), .A2(new_n355), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n897), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n610), .A2(new_n374), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n865), .A2(new_n963), .A3(new_n973), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n967), .A2(new_n972), .A3(new_n974), .ZN(G57));
endmodule


