//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 0 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT2), .ZN(new_n189));
  INV_X1    g003(.A(G113), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT66), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT2), .A3(G113), .ZN(new_n193));
  AOI22_X1  g007(.A1(new_n191), .A2(new_n193), .B1(new_n189), .B2(new_n190), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT67), .ZN(new_n195));
  INV_X1    g009(.A(G116), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n195), .B1(new_n196), .B2(G119), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT67), .A3(G116), .ZN(new_n199));
  AOI22_X1  g013(.A1(new_n197), .A2(new_n199), .B1(new_n196), .B2(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n194), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT3), .B1(new_n203), .B2(G107), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G104), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n203), .A2(G107), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n204), .A2(new_n207), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n203), .A2(G107), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n206), .A2(G104), .ZN(new_n212));
  OAI21_X1  g026(.A(G101), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n202), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT5), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT68), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n197), .A2(new_n199), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n196), .A2(G119), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n200), .A2(new_n217), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n216), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n198), .A2(G116), .ZN(new_n224));
  OAI21_X1  g038(.A(G113), .B1(new_n224), .B2(KEYINPUT5), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n215), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n204), .A2(new_n207), .A3(new_n209), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT4), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(G101), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n218), .A2(new_n217), .A3(new_n219), .ZN(new_n230));
  NOR3_X1   g044(.A1(new_n230), .A2(new_n220), .A3(new_n194), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n229), .B1(new_n231), .B2(new_n202), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n228), .B1(new_n227), .B2(G101), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT84), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n233), .A2(new_n234), .A3(new_n210), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n234), .B1(new_n233), .B2(new_n210), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n226), .B1(new_n232), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G110), .B(G122), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n226), .B(new_n239), .C1(new_n232), .C2(new_n237), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(KEYINPUT6), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(KEYINPUT1), .ZN(new_n245));
  INV_X1    g059(.A(G146), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G143), .ZN(new_n247));
  INV_X1    g061(.A(G143), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G146), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n245), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(KEYINPUT1), .A3(G146), .ZN(new_n251));
  XNOR2_X1  g065(.A(G143), .B(G146), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n250), .B(new_n251), .C1(G128), .C2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G125), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AND2_X1   g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n247), .A2(new_n249), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT64), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT64), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n252), .A2(new_n260), .A3(new_n257), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n247), .A2(new_n249), .ZN(new_n262));
  NOR2_X1   g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n259), .A2(new_n261), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n256), .B1(new_n255), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G953), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G224), .ZN(new_n268));
  XOR2_X1   g082(.A(new_n266), .B(new_n268), .Z(new_n269));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n238), .A2(new_n270), .A3(new_n240), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n243), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT89), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n268), .A2(new_n273), .A3(KEYINPUT7), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n273), .B1(new_n268), .B2(KEYINPUT7), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n266), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n275), .B1(new_n266), .B2(new_n274), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n239), .B(KEYINPUT8), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n210), .A2(new_n213), .ZN(new_n280));
  INV_X1    g094(.A(new_n225), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n230), .A2(new_n220), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n281), .B1(new_n282), .B2(new_n216), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n280), .B1(new_n283), .B2(new_n201), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT88), .B1(new_n200), .B2(KEYINPUT5), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(new_n225), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n200), .A2(KEYINPUT88), .A3(KEYINPUT5), .ZN(new_n287));
  AOI211_X1 g101(.A(new_n202), .B(new_n214), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n279), .B1(new_n284), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n278), .A2(new_n289), .A3(new_n242), .ZN(new_n290));
  INV_X1    g104(.A(G902), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G210), .B1(G237), .B2(G902), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n272), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT90), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n296), .B1(new_n272), .B2(new_n292), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n290), .A2(new_n291), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n243), .A2(new_n269), .A3(new_n271), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(KEYINPUT90), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n300), .A3(new_n294), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT91), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n295), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n297), .A2(new_n300), .A3(KEYINPUT91), .A4(new_n294), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n188), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT9), .B(G234), .ZN(new_n306));
  OAI21_X1  g120(.A(G221), .B1(new_n306), .B2(G902), .ZN(new_n307));
  XOR2_X1   g121(.A(new_n307), .B(KEYINPUT83), .Z(new_n308));
  INV_X1    g122(.A(G469), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT12), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT11), .ZN(new_n311));
  INV_X1    g125(.A(G134), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n311), .B1(new_n312), .B2(G137), .ZN(new_n313));
  AOI21_X1  g127(.A(G131), .B1(new_n312), .B2(G137), .ZN(new_n314));
  INV_X1    g128(.A(G137), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(KEYINPUT11), .A3(G134), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n313), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT65), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT65), .A4(new_n316), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n313), .A2(new_n316), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n315), .A2(G134), .ZN(new_n323));
  OAI21_X1  g137(.A(G131), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT69), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n321), .A2(KEYINPUT69), .A3(new_n324), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n253), .B(new_n214), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n310), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n325), .ZN(new_n332));
  OR3_X1    g146(.A1(new_n330), .A2(new_n332), .A3(new_n310), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(G110), .B(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n267), .A2(G227), .ZN(new_n336));
  XOR2_X1   g150(.A(new_n335), .B(new_n336), .Z(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT85), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n259), .A2(new_n261), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n262), .A2(new_n264), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(new_n229), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n227), .A2(G101), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(KEYINPUT4), .A3(new_n210), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT84), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n233), .A2(new_n234), .A3(new_n210), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n342), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT10), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n348), .B1(new_n254), .B2(new_n214), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n280), .A2(KEYINPUT10), .A3(new_n253), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n339), .B1(new_n352), .B2(new_n329), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n340), .A2(new_n341), .A3(new_n229), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n235), .B2(new_n236), .ZN(new_n355));
  AND4_X1   g169(.A1(KEYINPUT10), .A2(new_n253), .A3(new_n210), .A4(new_n213), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT10), .B1(new_n280), .B2(new_n253), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n329), .A2(new_n355), .A3(new_n358), .A4(new_n339), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n334), .B(new_n338), .C1(new_n353), .C2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n329), .A2(new_n355), .A3(new_n358), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT85), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n359), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n352), .A2(new_n329), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n338), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n309), .B(new_n291), .C1(new_n362), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT87), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n352), .A2(new_n329), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n370), .B1(new_n364), .B2(new_n359), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n361), .B1(new_n371), .B2(new_n338), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT87), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n372), .A2(new_n373), .A3(new_n309), .A4(new_n291), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n338), .B1(new_n365), .B2(new_n334), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n337), .B1(new_n364), .B2(new_n359), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n370), .B1(new_n377), .B2(KEYINPUT86), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n338), .B1(new_n353), .B2(new_n360), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT86), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n376), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(G469), .B1(new_n382), .B2(G902), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n308), .B1(new_n375), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(G475), .A2(G902), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT71), .B(G237), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(G214), .A3(new_n267), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n248), .ZN(new_n388));
  OR2_X1    g202(.A1(KEYINPUT71), .A2(G237), .ZN(new_n389));
  NAND2_X1  g203(.A1(KEYINPUT71), .A2(G237), .ZN(new_n390));
  AOI21_X1  g204(.A(G953), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(G143), .A3(G214), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G131), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT17), .ZN(new_n395));
  INV_X1    g209(.A(G131), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n388), .A2(new_n396), .A3(new_n392), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT93), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n394), .A2(KEYINPUT93), .A3(new_n395), .A4(new_n397), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT16), .ZN(new_n402));
  XNOR2_X1  g216(.A(G125), .B(G140), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT79), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G140), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(KEYINPUT79), .A3(G125), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n402), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n255), .A2(KEYINPUT16), .A3(G140), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n246), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n409), .ZN(new_n411));
  INV_X1    g225(.A(new_n407), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(new_n404), .B2(new_n403), .ZN(new_n413));
  OAI211_X1 g227(.A(G146), .B(new_n411), .C1(new_n413), .C2(new_n402), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  AOI211_X1 g229(.A(new_n395), .B(new_n396), .C1(new_n388), .C2(new_n392), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n400), .A2(new_n401), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n403), .A2(new_n246), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n405), .A2(new_n407), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n419), .B1(new_n420), .B2(new_n246), .ZN(new_n421));
  NAND2_X1  g235(.A1(KEYINPUT18), .A2(G131), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n388), .A2(new_n392), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n423), .B1(new_n388), .B2(new_n392), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT92), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT92), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n428), .B(new_n421), .C1(new_n424), .C2(new_n425), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(G113), .B(G122), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(new_n203), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n418), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n420), .A2(KEYINPUT19), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(KEYINPUT19), .B2(new_n403), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n246), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n394), .A2(new_n397), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(new_n437), .A3(new_n414), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n432), .B1(new_n430), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n385), .B1(new_n433), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT94), .ZN(new_n441));
  INV_X1    g255(.A(new_n425), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n388), .A2(new_n392), .A3(new_n423), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n428), .B1(new_n444), .B2(new_n421), .ZN(new_n445));
  INV_X1    g259(.A(new_n429), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n438), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n432), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n418), .A2(new_n430), .A3(new_n432), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n441), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n440), .B1(new_n451), .B2(KEYINPUT20), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n449), .A2(new_n450), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT20), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n453), .A2(new_n441), .A3(new_n454), .A4(new_n385), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n432), .B1(new_n418), .B2(new_n430), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n291), .B1(new_n433), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G475), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(G234), .A2(G237), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n461), .A2(G952), .A3(new_n267), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n461), .A2(G902), .A3(G953), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(G898), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G478), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n466), .A2(KEYINPUT15), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n196), .A2(KEYINPUT14), .A3(G122), .ZN(new_n469));
  XNOR2_X1  g283(.A(G116), .B(G122), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  OAI211_X1 g285(.A(G107), .B(new_n469), .C1(new_n471), .C2(KEYINPUT14), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n206), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n248), .A2(G128), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n244), .A2(G143), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(new_n475), .A3(new_n312), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n312), .B1(new_n474), .B2(new_n475), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n472), .B(new_n473), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(KEYINPUT95), .B(KEYINPUT13), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n474), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT96), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n480), .A2(new_n474), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(new_n244), .B2(G143), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n312), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n471), .A2(G107), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n487), .A2(new_n473), .B1(KEYINPUT97), .B2(new_n476), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(KEYINPUT97), .B2(new_n476), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n479), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G217), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n306), .A2(new_n491), .A3(G953), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n492), .B(new_n479), .C1(new_n486), .C2(new_n489), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n468), .B1(new_n496), .B2(new_n291), .ZN(new_n497));
  AOI211_X1 g311(.A(G902), .B(new_n467), .C1(new_n494), .C2(new_n495), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT98), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT98), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n501), .B1(new_n497), .B2(new_n498), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n460), .A2(new_n465), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n305), .A2(new_n384), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(G234), .ZN(new_n506));
  OAI21_X1  g320(.A(G217), .B1(new_n506), .B2(G902), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n267), .A2(G221), .A3(G234), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(KEYINPUT22), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(new_n315), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT81), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n244), .A2(KEYINPUT23), .A3(G119), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n198), .A2(G128), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n244), .A2(G119), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n514), .B(new_n515), .C1(new_n517), .C2(KEYINPUT23), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G110), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT78), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT78), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n518), .A2(new_n521), .A3(G110), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT76), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n244), .B2(G119), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n198), .A2(KEYINPUT76), .A3(G128), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n516), .A3(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT24), .B(G110), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT77), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n525), .A2(new_n516), .ZN(new_n529));
  INV_X1    g343(.A(new_n527), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT77), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n529), .A2(new_n530), .A3(new_n531), .A4(new_n524), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n520), .A2(new_n522), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n419), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n409), .B1(new_n420), .B2(KEYINPUT16), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n534), .B1(new_n535), .B2(G146), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n526), .A2(new_n527), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT80), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n526), .A2(KEYINPUT80), .A3(new_n527), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n539), .B(new_n540), .C1(G110), .C2(new_n518), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n415), .A2(new_n533), .B1(new_n536), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n510), .A2(KEYINPUT81), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n513), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n533), .A2(new_n415), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n536), .A2(new_n541), .ZN(new_n546));
  AND4_X1   g360(.A1(new_n513), .A2(new_n545), .A3(new_n546), .A4(new_n543), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n291), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n507), .B1(new_n548), .B2(KEYINPUT25), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT25), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n550), .B(new_n291), .C1(new_n544), .C2(new_n547), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n544), .A2(new_n547), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n507), .A2(new_n291), .ZN(new_n554));
  OR2_X1    g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n327), .A2(new_n328), .A3(new_n265), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT70), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT70), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n327), .A2(new_n560), .A3(new_n328), .A4(new_n265), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n312), .A2(G137), .ZN(new_n562));
  OAI21_X1  g376(.A(G131), .B1(new_n562), .B2(new_n323), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n321), .A2(new_n563), .A3(new_n253), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n559), .A2(KEYINPUT30), .A3(new_n561), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n221), .A2(new_n222), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n201), .B1(new_n566), .B2(new_n194), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n265), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n564), .B1(new_n332), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT30), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n568), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n565), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n564), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n567), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n559), .A2(new_n561), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n391), .A2(G210), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT27), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT26), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT27), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n391), .A2(new_n580), .A3(G210), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n579), .B1(new_n578), .B2(new_n581), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n208), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n584), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(G101), .A3(new_n582), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n576), .A2(KEYINPUT72), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT72), .B1(new_n576), .B2(new_n589), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n573), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT73), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT73), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n594), .B(new_n573), .C1(new_n590), .C2(new_n591), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n593), .A2(KEYINPUT31), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT31), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n597), .B(new_n573), .C1(new_n590), .C2(new_n591), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n558), .A2(new_n564), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n567), .B1(new_n599), .B2(KEYINPUT74), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT74), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n558), .A2(new_n601), .A3(new_n564), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT28), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT28), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n570), .A2(new_n567), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n604), .B1(new_n576), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n588), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n598), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n596), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(G472), .A2(G902), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT32), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n589), .A2(KEYINPUT29), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT75), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n559), .A2(new_n561), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n559), .A2(new_n561), .A3(new_n564), .ZN(new_n618));
  AOI22_X1  g432(.A1(new_n617), .A2(new_n575), .B1(new_n618), .B2(new_n567), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n616), .B1(new_n619), .B2(new_n604), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n567), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n576), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(KEYINPUT75), .A3(KEYINPUT28), .ZN(new_n623));
  AOI211_X1 g437(.A(new_n603), .B(new_n615), .C1(new_n620), .C2(new_n623), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n321), .A2(KEYINPUT69), .A3(new_n324), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT69), .B1(new_n321), .B2(new_n324), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n625), .A2(new_n626), .A3(new_n569), .ZN(new_n627));
  OAI21_X1  g441(.A(KEYINPUT74), .B1(new_n627), .B2(new_n574), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n628), .A2(new_n568), .A3(new_n602), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n604), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n576), .A2(new_n605), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n630), .B(new_n589), .C1(new_n631), .C2(new_n604), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n573), .A2(new_n576), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n588), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT29), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n632), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n291), .ZN(new_n637));
  OAI21_X1  g451(.A(G472), .B1(new_n624), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n614), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n611), .B1(new_n596), .B2(new_n608), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(KEYINPUT32), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n557), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT82), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n614), .B(new_n638), .C1(KEYINPUT32), .C2(new_n640), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT82), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(new_n645), .A3(new_n557), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n505), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT99), .B(G101), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT100), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n647), .B(new_n649), .ZN(G3));
  NAND2_X1  g464(.A1(new_n609), .A2(new_n291), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n651), .A2(KEYINPUT101), .A3(G472), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n653));
  AOI21_X1  g467(.A(G902), .B1(new_n596), .B2(new_n608), .ZN(new_n654));
  INV_X1    g468(.A(G472), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n609), .A2(new_n610), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n652), .A2(new_n656), .A3(new_n657), .A4(new_n384), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n658), .A2(new_n556), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n496), .B(KEYINPUT33), .Z(new_n660));
  NOR2_X1   g474(.A1(new_n466), .A2(G902), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(G902), .B1(new_n494), .B2(new_n495), .ZN(new_n663));
  OAI22_X1  g477(.A1(new_n660), .A2(new_n662), .B1(G478), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n460), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n293), .B1(new_n298), .B2(new_n299), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n187), .B1(new_n295), .B2(new_n666), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n665), .A2(new_n465), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n659), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT34), .B(G104), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT102), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n670), .B(new_n672), .ZN(G6));
  AOI21_X1  g487(.A(new_n454), .B1(new_n453), .B2(new_n385), .ZN(new_n674));
  INV_X1    g488(.A(new_n385), .ZN(new_n675));
  AOI211_X1 g489(.A(KEYINPUT20), .B(new_n675), .C1(new_n449), .C2(new_n450), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n503), .B(new_n459), .C1(new_n674), .C2(new_n676), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n677), .A2(new_n667), .A3(new_n465), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n659), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n680), .B(KEYINPUT103), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT35), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G107), .ZN(G9));
  NOR2_X1   g497(.A1(new_n510), .A2(KEYINPUT36), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n545), .A2(new_n546), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(KEYINPUT104), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n542), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n685), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n686), .A2(KEYINPUT104), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n542), .A2(new_n688), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n691), .A2(new_n692), .A3(new_n684), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n554), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n694), .B1(new_n549), .B2(new_n551), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n504), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n305), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n658), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT37), .B(G110), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G12));
  INV_X1    g515(.A(G900), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n462), .B1(new_n463), .B2(new_n702), .ZN(new_n703));
  NOR4_X1   g517(.A1(new_n677), .A2(new_n667), .A3(new_n695), .A4(new_n703), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n704), .B(new_n384), .C1(new_n639), .C2(new_n641), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G128), .ZN(G30));
  NAND2_X1  g520(.A1(new_n303), .A2(new_n304), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT38), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT38), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n303), .A2(new_n709), .A3(new_n304), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  AOI22_X1  g525(.A1(new_n452), .A2(new_n455), .B1(G475), .B2(new_n458), .ZN(new_n712));
  INV_X1    g526(.A(new_n503), .ZN(new_n713));
  NOR4_X1   g527(.A1(new_n712), .A2(new_n713), .A3(new_n696), .A4(new_n188), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(new_n703), .B(KEYINPUT39), .Z(new_n716));
  NAND2_X1  g530(.A1(new_n384), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT40), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n622), .A2(new_n588), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n593), .A2(new_n595), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n291), .ZN(new_n722));
  AOI22_X1  g536(.A1(G472), .A2(new_n722), .B1(new_n609), .B2(new_n613), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n657), .A2(new_n612), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n725), .B1(new_n723), .B2(new_n724), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n719), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n722), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n614), .B1(new_n729), .B2(new_n655), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT105), .B1(new_n730), .B2(new_n641), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(new_n732), .A3(KEYINPUT106), .ZN(new_n733));
  AOI211_X1 g547(.A(new_n715), .B(new_n718), .C1(new_n728), .C2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n248), .ZN(G45));
  INV_X1    g549(.A(new_n703), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n460), .A2(new_n664), .A3(new_n736), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n696), .B(new_n187), .C1(new_n295), .C2(new_n666), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n739), .B(new_n384), .C1(new_n639), .C2(new_n641), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G146), .ZN(G48));
  NOR3_X1   g555(.A1(new_n619), .A2(new_n616), .A3(new_n604), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT75), .B1(new_n622), .B2(KEYINPUT28), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n630), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n291), .B(new_n636), .C1(new_n744), .C2(new_n615), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n745), .A2(G472), .B1(new_n609), .B2(new_n613), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n556), .B1(new_n746), .B2(new_n724), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT107), .ZN(new_n748));
  INV_X1    g562(.A(new_n308), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n309), .B1(new_n372), .B2(new_n291), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  AND4_X1   g565(.A1(new_n748), .A2(new_n375), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n750), .B1(new_n369), .B2(new_n374), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n748), .B1(new_n753), .B2(new_n749), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n747), .A2(new_n668), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(KEYINPUT41), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G113), .ZN(G15));
  NAND4_X1  g572(.A1(new_n755), .A2(new_n644), .A3(new_n557), .A4(new_n678), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G116), .ZN(G18));
  INV_X1    g574(.A(new_n667), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n755), .A2(new_n644), .A3(new_n697), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G119), .ZN(G21));
  AOI21_X1  g577(.A(new_n603), .B1(new_n620), .B2(new_n623), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n596), .B(new_n598), .C1(new_n589), .C2(new_n764), .ZN(new_n765));
  AOI22_X1  g579(.A1(new_n651), .A2(G472), .B1(new_n765), .B2(new_n610), .ZN(new_n766));
  NOR4_X1   g580(.A1(new_n667), .A2(new_n712), .A3(new_n713), .A4(new_n465), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n755), .A2(new_n557), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G122), .ZN(G24));
  NAND2_X1  g583(.A1(new_n651), .A2(G472), .ZN(new_n770));
  INV_X1    g584(.A(new_n737), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n765), .A2(new_n610), .ZN(new_n772));
  AND4_X1   g586(.A1(new_n770), .A2(new_n696), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n375), .A2(new_n749), .A3(new_n751), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT107), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n753), .A2(new_n748), .A3(new_n749), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n761), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G125), .ZN(G27));
  NAND3_X1  g594(.A1(new_n303), .A2(new_n187), .A3(new_n304), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n366), .B1(new_n353), .B2(new_n360), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n337), .ZN(new_n783));
  AOI21_X1  g597(.A(G902), .B1(new_n783), .B2(new_n361), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n373), .B1(new_n784), .B2(new_n309), .ZN(new_n785));
  INV_X1    g599(.A(new_n374), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n383), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n749), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT108), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT108), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n384), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n781), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT42), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT109), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n792), .A2(new_n747), .A3(new_n771), .A4(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n781), .ZN(new_n796));
  AOI211_X1 g610(.A(KEYINPUT108), .B(new_n308), .C1(new_n375), .C2(new_n383), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n790), .B1(new_n787), .B2(new_n749), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n799), .A2(new_n642), .A3(new_n737), .ZN(new_n800));
  XNOR2_X1  g614(.A(KEYINPUT109), .B(KEYINPUT42), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n795), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G131), .ZN(G33));
  NOR2_X1   g617(.A1(new_n677), .A2(new_n703), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n792), .A2(new_n747), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G134), .ZN(G36));
  NAND2_X1  g620(.A1(new_n712), .A2(new_n664), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT43), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT43), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n712), .A2(new_n809), .A3(new_n664), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n652), .A2(new_n657), .A3(new_n656), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n811), .A2(new_n812), .A3(new_n696), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n812), .B1(new_n811), .B2(new_n696), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n808), .B(new_n810), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT44), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  NAND2_X1  g632(.A1(G469), .A2(G902), .ZN(new_n819));
  OAI21_X1  g633(.A(G469), .B1(new_n382), .B2(KEYINPUT45), .ZN(new_n820));
  INV_X1    g634(.A(new_n376), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n366), .B1(new_n379), .B2(new_n380), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n377), .A2(KEYINPUT86), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT45), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT110), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n820), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n309), .B1(new_n824), .B2(new_n825), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n382), .A2(KEYINPUT45), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT110), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n819), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT46), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n827), .B1(new_n820), .B2(new_n826), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n829), .A2(KEYINPUT110), .A3(new_n830), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n835), .A2(new_n836), .B1(G469), .B2(G902), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT46), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n834), .A2(new_n838), .A3(new_n375), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n839), .A2(new_n749), .A3(new_n716), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n781), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n817), .A2(new_n818), .A3(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(G137), .ZN(G39));
  OAI21_X1  g657(.A(new_n375), .B1(new_n837), .B2(KEYINPUT46), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n832), .A2(new_n833), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n749), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT47), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT47), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n839), .A2(new_n848), .A3(new_n749), .ZN(new_n849));
  NOR4_X1   g663(.A1(new_n644), .A2(new_n557), .A3(new_n781), .A4(new_n737), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(G140), .ZN(G42));
  NAND2_X1  g666(.A1(new_n775), .A2(new_n776), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n711), .A2(new_n187), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n770), .A2(new_n557), .A3(new_n772), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n808), .A2(new_n462), .A3(new_n810), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT113), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT113), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n808), .A2(new_n858), .A3(new_n462), .A4(new_n810), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n855), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(KEYINPUT114), .A2(KEYINPUT50), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(KEYINPUT114), .A2(KEYINPUT50), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n862), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n854), .B2(new_n860), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n863), .A2(KEYINPUT115), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT115), .ZN(new_n868));
  INV_X1    g682(.A(new_n866), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n854), .B(new_n860), .C1(KEYINPUT114), .C2(KEYINPUT50), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n853), .A2(new_n781), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n873), .A2(new_n557), .A3(new_n462), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n460), .A2(new_n664), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n874), .A2(new_n728), .A3(new_n733), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n857), .A2(new_n859), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n877), .A2(new_n873), .A3(new_n696), .A4(new_n766), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n847), .A2(new_n849), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n753), .B(KEYINPUT112), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n308), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n860), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n884), .A2(new_n781), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n879), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT51), .B1(new_n872), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n877), .A2(new_n747), .A3(new_n873), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT48), .ZN(new_n889));
  INV_X1    g703(.A(new_n665), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n874), .A2(new_n728), .A3(new_n890), .A4(new_n733), .ZN(new_n891));
  INV_X1    g705(.A(G952), .ZN(new_n892));
  AOI211_X1 g706(.A(new_n892), .B(G953), .C1(new_n860), .C2(new_n778), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n889), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  AOI22_X1  g708(.A1(new_n847), .A2(new_n849), .B1(new_n308), .B2(new_n881), .ZN(new_n895));
  INV_X1    g709(.A(new_n885), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n878), .B(new_n876), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT51), .B1(new_n863), .B2(new_n866), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n887), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT52), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n770), .A2(new_n771), .A3(new_n772), .A4(new_n696), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n705), .B(new_n740), .C1(new_n903), .C2(new_n777), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n667), .A2(new_n712), .A3(new_n713), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n384), .A2(new_n905), .A3(new_n695), .A4(new_n736), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n731), .B2(new_n732), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n902), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n906), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(new_n726), .B2(new_n727), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n644), .B(new_n384), .C1(new_n704), .C2(new_n739), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n910), .A2(KEYINPUT52), .A3(new_n779), .A4(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n773), .A2(new_n792), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n459), .B1(new_n674), .B2(new_n676), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n499), .A2(new_n736), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n915), .A2(new_n695), .A3(new_n916), .ZN(new_n917));
  AND4_X1   g731(.A1(new_n187), .A2(new_n303), .A3(new_n917), .A4(new_n304), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n644), .A2(new_n918), .A3(new_n384), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n805), .A2(new_n914), .A3(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n756), .A2(new_n759), .A3(new_n762), .A4(new_n768), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n665), .B1(new_n460), .B2(new_n499), .ZN(new_n923));
  INV_X1    g737(.A(new_n465), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n305), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n658), .A2(new_n925), .A3(new_n556), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n647), .A2(new_n699), .A3(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n913), .A2(new_n922), .A3(new_n802), .A4(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT53), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n644), .A2(new_n668), .A3(new_n557), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n644), .A2(new_n557), .A3(new_n678), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n853), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n697), .A2(new_n644), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n767), .A2(new_n775), .A3(new_n776), .ZN(new_n935));
  OAI22_X1  g749(.A1(new_n934), .A2(new_n777), .B1(new_n935), .B2(new_n855), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n804), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n799), .A2(new_n642), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n919), .B1(new_n799), .B2(new_n903), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n802), .A2(new_n937), .A3(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n942), .A2(KEYINPUT53), .A3(new_n913), .A4(new_n927), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n901), .B1(new_n930), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n930), .A2(new_n901), .A3(new_n943), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n900), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT116), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT116), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n900), .A2(new_n949), .A3(new_n945), .A4(new_n946), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n892), .A2(new_n267), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n948), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n881), .B(KEYINPUT49), .ZN(new_n953));
  NOR4_X1   g767(.A1(new_n807), .A2(new_n556), .A3(new_n188), .A4(new_n308), .ZN(new_n954));
  AND4_X1   g768(.A1(new_n708), .A2(new_n953), .A3(new_n710), .A4(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n955), .A2(new_n728), .A3(new_n733), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n952), .A2(new_n956), .ZN(G75));
  NOR2_X1   g771(.A1(new_n267), .A2(G952), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n291), .B1(new_n930), .B2(new_n943), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT56), .B1(new_n960), .B2(G210), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n243), .A2(new_n271), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(new_n269), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT55), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n959), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT56), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n930), .A2(new_n943), .ZN(new_n968));
  AOI21_X1  g782(.A(KEYINPUT117), .B1(new_n968), .B2(G902), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT117), .ZN(new_n970));
  AOI211_X1 g784(.A(new_n970), .B(new_n291), .C1(new_n930), .C2(new_n943), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n294), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT118), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n967), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n960), .B(KEYINPUT117), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n975), .A2(KEYINPUT118), .A3(new_n294), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n965), .B1(new_n974), .B2(new_n976), .ZN(G51));
  XOR2_X1   g791(.A(new_n819), .B(KEYINPUT57), .Z(new_n978));
  AND3_X1   g792(.A1(new_n930), .A2(new_n901), .A3(new_n943), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n978), .B1(new_n979), .B2(new_n944), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT119), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g796(.A(KEYINPUT119), .B(new_n978), .C1(new_n979), .C2(new_n944), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n982), .A2(new_n372), .A3(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n975), .A2(new_n835), .A3(new_n836), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n958), .B1(new_n984), .B2(new_n985), .ZN(G54));
  NAND2_X1  g800(.A1(KEYINPUT58), .A2(G475), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT120), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n453), .B1(new_n975), .B2(new_n988), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n453), .B(new_n988), .C1(new_n969), .C2(new_n971), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n959), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n989), .A2(new_n991), .ZN(G60));
  INV_X1    g806(.A(new_n660), .ZN(new_n993));
  NAND2_X1  g807(.A1(G478), .A2(G902), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT59), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n993), .B(new_n995), .C1(new_n979), .C2(new_n944), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n996), .A2(KEYINPUT121), .A3(new_n959), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n995), .B1(new_n979), .B2(new_n944), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n660), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(KEYINPUT121), .B1(new_n996), .B2(new_n959), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n1000), .A2(new_n1001), .ZN(G63));
  AND2_X1   g816(.A1(new_n930), .A2(new_n943), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n690), .A2(new_n693), .ZN(new_n1004));
  NAND2_X1  g818(.A1(G217), .A2(G902), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT122), .Z(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT60), .ZN(new_n1007));
  OR3_X1    g821(.A1(new_n1003), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n553), .B1(new_n1003), .B2(new_n1007), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1008), .A2(new_n959), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT61), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1008), .A2(KEYINPUT61), .A3(new_n959), .A4(new_n1009), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1012), .A2(new_n1013), .ZN(G66));
  INV_X1    g828(.A(G224), .ZN(new_n1015));
  OAI21_X1  g829(.A(G953), .B1(new_n464), .B2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1016), .B(KEYINPUT123), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n927), .A2(new_n937), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1017), .B1(new_n1018), .B2(G953), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n962), .B1(G898), .B2(new_n267), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1019), .B(new_n1020), .ZN(G69));
  OR3_X1    g835(.A1(new_n734), .A2(KEYINPUT62), .A3(new_n904), .ZN(new_n1022));
  OAI21_X1  g836(.A(KEYINPUT62), .B1(new_n734), .B2(new_n904), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n923), .B(KEYINPUT124), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n1024), .A2(new_n717), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n643), .A2(new_n646), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1025), .A2(new_n1026), .A3(new_n796), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n1022), .A2(new_n1023), .A3(new_n851), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(new_n842), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n267), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n570), .A2(new_n571), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n565), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1032), .B(new_n435), .ZN(new_n1033));
  AND2_X1   g847(.A1(new_n747), .A2(new_n905), .ZN(new_n1034));
  NAND4_X1  g848(.A1(new_n839), .A2(new_n1034), .A3(new_n749), .A4(new_n716), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1035), .B(KEYINPUT126), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n904), .A2(new_n939), .ZN(new_n1037));
  AND3_X1   g851(.A1(new_n851), .A2(new_n802), .A3(new_n1037), .ZN(new_n1038));
  NAND4_X1  g852(.A1(new_n842), .A2(new_n267), .A3(new_n1036), .A4(new_n1038), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1033), .B1(G900), .B2(G953), .ZN(new_n1040));
  AOI22_X1  g854(.A1(new_n1030), .A2(new_n1033), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g855(.A(KEYINPUT125), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n267), .B1(G227), .B2(G900), .ZN(new_n1043));
  NOR2_X1   g857(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g858(.A(new_n1041), .B(new_n1044), .ZN(G72));
  NAND2_X1  g859(.A1(G472), .A2(G902), .ZN(new_n1046));
  XOR2_X1   g860(.A(new_n1046), .B(KEYINPUT63), .Z(new_n1047));
  INV_X1    g861(.A(new_n1047), .ZN(new_n1048));
  AND2_X1   g862(.A1(new_n593), .A2(new_n595), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1048), .B1(new_n1049), .B2(new_n634), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n958), .B1(new_n968), .B2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g865(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n1048), .B1(new_n1052), .B2(new_n1018), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n633), .A2(new_n589), .ZN(new_n1054));
  OAI21_X1  g868(.A(new_n1051), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g869(.A1(new_n842), .A2(new_n1018), .A3(new_n1036), .A4(new_n1038), .ZN(new_n1056));
  INV_X1    g870(.A(KEYINPUT127), .ZN(new_n1057));
  NAND3_X1  g871(.A1(new_n1056), .A2(new_n1057), .A3(new_n1047), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n1057), .B1(new_n1056), .B2(new_n1047), .ZN(new_n1059));
  NOR3_X1   g873(.A1(new_n1059), .A2(new_n589), .A3(new_n633), .ZN(new_n1060));
  AOI21_X1  g874(.A(new_n1055), .B1(new_n1058), .B2(new_n1060), .ZN(G57));
endmodule


