//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n606, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218, new_n1219;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT67), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OR2_X1    g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n469), .B1(new_n463), .B2(new_n464), .ZN(new_n470));
  AND2_X1   g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  AND2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n468), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n478), .B(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G2104), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  AOI22_X1  g060(.A1(new_n481), .A2(G136), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n480), .A2(new_n486), .ZN(G162));
  OAI21_X1  g062(.A(G2104), .B1(new_n468), .B2(G114), .ZN(new_n488));
  NOR2_X1   g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT69), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n491), .A2(new_n493), .A3(new_n494), .A4(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n468), .C1(new_n474), .C2(new_n475), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(G126), .B(G2105), .C1(new_n474), .C2(new_n475), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT4), .A2(G138), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n468), .B(new_n501), .C1(new_n474), .C2(new_n475), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n496), .A2(new_n499), .A3(new_n500), .A4(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT70), .B1(new_n505), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n505), .A2(G543), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n510), .A2(G88), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(G543), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n510), .A2(G62), .A3(new_n511), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n516), .A2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  AND2_X1   g097(.A1(new_n510), .A2(new_n511), .ZN(new_n523));
  AND2_X1   g098(.A1(G76), .A2(G543), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n523), .A2(G63), .B1(KEYINPUT7), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n517), .ZN(new_n526));
  AOI21_X1  g101(.A(KEYINPUT7), .B1(new_n524), .B2(G651), .ZN(new_n527));
  INV_X1    g102(.A(new_n515), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n527), .B1(new_n528), .B2(G51), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n523), .A2(new_n512), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT71), .B(G89), .Z(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n526), .A2(new_n532), .ZN(G168));
  AOI22_X1  g108(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n517), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n528), .A2(G52), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n530), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n535), .A2(new_n538), .ZN(G171));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n510), .A2(new_n511), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G651), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n510), .A2(G81), .A3(new_n511), .A4(new_n512), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT72), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n512), .A2(G43), .A3(G543), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n546), .B1(new_n545), .B2(new_n547), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n544), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(new_n517), .A2(KEYINPUT6), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT6), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G651), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n557), .A2(new_n559), .A3(G53), .A4(G543), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT9), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n512), .A2(new_n562), .A3(G53), .A4(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n510), .A2(G91), .A3(new_n511), .A4(new_n512), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n510), .A2(G65), .A3(new_n511), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n517), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  NAND2_X1  g148(.A1(new_n528), .A2(G49), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n510), .A2(G87), .A3(new_n511), .A4(new_n512), .ZN(new_n575));
  AOI21_X1  g150(.A(G74), .B1(new_n510), .B2(new_n511), .ZN(new_n576));
  OAI211_X1 g151(.A(new_n574), .B(new_n575), .C1(new_n517), .C2(new_n576), .ZN(G288));
  NAND3_X1  g152(.A1(new_n510), .A2(G61), .A3(new_n511), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n510), .A2(G86), .A3(new_n511), .A4(new_n512), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n512), .A2(G48), .A3(G543), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n581), .A2(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(new_n528), .A2(G47), .ZN(new_n586));
  INV_X1    g161(.A(G85), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OAI221_X1 g163(.A(new_n586), .B1(new_n530), .B2(new_n587), .C1(new_n588), .C2(new_n517), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n523), .A2(G92), .A3(new_n512), .ZN(new_n591));
  XOR2_X1   g166(.A(new_n591), .B(KEYINPUT10), .Z(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n541), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(G54), .B2(new_n528), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n590), .B1(G868), .B2(new_n597), .ZN(G284));
  OAI21_X1  g173(.A(new_n590), .B1(G868), .B2(new_n597), .ZN(G321));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(G299), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(G168), .B2(new_n600), .ZN(G297));
  OAI21_X1  g177(.A(new_n601), .B1(G168), .B2(new_n600), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n597), .B1(new_n604), .B2(G860), .ZN(G148));
  NAND2_X1  g180(.A1(new_n550), .A2(new_n600), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n592), .A2(new_n596), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n606), .B1(new_n608), .B2(new_n600), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n481), .A2(G2104), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT73), .Z(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT13), .ZN(new_n614));
  INV_X1    g189(.A(G2100), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT74), .Z(new_n617));
  NAND2_X1  g192(.A1(new_n477), .A2(G123), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n481), .A2(G135), .ZN(new_n619));
  NOR2_X1   g194(.A1(G99), .A2(G2105), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(new_n468), .B2(G111), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2096), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n623), .B1(new_n614), .B2(new_n615), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n617), .A2(new_n624), .ZN(G156));
  XOR2_X1   g200(.A(G1341), .B(G1348), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT77), .ZN(new_n627));
  XOR2_X1   g202(.A(G2451), .B(G2454), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n627), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT76), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2438), .Z(new_n636));
  XOR2_X1   g211(.A(G2427), .B(G2430), .Z(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(KEYINPUT75), .B(KEYINPUT14), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n636), .A2(new_n637), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n633), .A2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(G14), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n633), .A2(new_n641), .ZN(new_n644));
  NOR3_X1   g219(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(G401));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2072), .B(G2078), .Z(new_n649));
  NOR2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT18), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n649), .B(KEYINPUT17), .ZN(new_n652));
  INV_X1    g227(.A(new_n646), .ZN(new_n653));
  INV_X1    g228(.A(new_n647), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n653), .A2(new_n649), .A3(new_n654), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(new_n648), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n651), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2096), .B(G2100), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT78), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  AND2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT20), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n664), .A2(new_n665), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n663), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n663), .B2(new_n669), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1981), .B(G1986), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT79), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n672), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1991), .B(G1996), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(G229));
  INV_X1    g256(.A(G1986), .ZN(new_n682));
  NAND2_X1  g257(.A1(G290), .A2(G16), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT80), .ZN(new_n684));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G24), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n683), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n684), .B1(new_n683), .B2(new_n686), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n682), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n689), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n691), .A2(G1986), .A3(new_n687), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT81), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n690), .A2(new_n692), .A3(KEYINPUT81), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n477), .A2(G119), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n481), .A2(G131), .ZN(new_n698));
  NOR2_X1   g273(.A1(G95), .A2(G2105), .ZN(new_n699));
  OAI21_X1  g274(.A(G2104), .B1(new_n468), .B2(G107), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n697), .B(new_n698), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(G25), .B(new_n701), .S(G29), .Z(new_n702));
  XOR2_X1   g277(.A(KEYINPUT35), .B(G1991), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n695), .A2(new_n696), .A3(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT33), .B(G1976), .Z(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n685), .A2(G23), .ZN(new_n708));
  INV_X1    g283(.A(G288), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n685), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(KEYINPUT83), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n710), .A2(KEYINPUT83), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n707), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n713), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n715), .A2(new_n706), .A3(new_n711), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(KEYINPUT84), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(KEYINPUT84), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n685), .A2(G22), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT85), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G166), .B2(new_n685), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G1971), .ZN(new_n723));
  INV_X1    g298(.A(G305), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G16), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G6), .B2(G16), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(KEYINPUT32), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n726), .A2(KEYINPUT32), .ZN(new_n729));
  OAI21_X1  g304(.A(G1981), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n726), .A2(KEYINPUT32), .ZN(new_n731));
  INV_X1    g306(.A(G1981), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n731), .A2(new_n732), .A3(new_n727), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n723), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  AND3_X1   g309(.A1(new_n718), .A2(new_n719), .A3(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT82), .B(KEYINPUT34), .Z(new_n736));
  AOI21_X1  g311(.A(new_n705), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(KEYINPUT87), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n718), .A2(new_n734), .A3(new_n719), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT86), .ZN(new_n741));
  INV_X1    g316(.A(new_n736), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n741), .B1(new_n740), .B2(new_n742), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n737), .B(new_n739), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G29), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n747), .A2(G33), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT25), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n751), .A2(new_n752), .B1(new_n481), .B2(G139), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT88), .ZN(new_n754));
  NAND2_X1  g329(.A1(G115), .A2(G2104), .ZN(new_n755));
  INV_X1    g330(.A(G127), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n476), .B2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT89), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n468), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n758), .B2(new_n757), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n754), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n748), .B1(new_n761), .B2(G29), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G2072), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT90), .Z(new_n765));
  NOR2_X1   g340(.A1(G5), .A2(G16), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT96), .Z(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G171), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT97), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n765), .B1(G1961), .B2(new_n769), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(G1961), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT92), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT93), .B(KEYINPUT26), .ZN(new_n774));
  NAND3_X1  g349(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n773), .B(new_n776), .C1(G129), .C2(new_n477), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n481), .A2(G141), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT91), .Z(new_n779));
  NAND2_X1  g354(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(new_n747), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT94), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G29), .B2(G32), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT27), .B(G1996), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n783), .A2(new_n785), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n770), .B(new_n771), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G162), .A2(new_n747), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n747), .A2(G35), .ZN(new_n790));
  OR3_X1    g365(.A1(new_n789), .A2(KEYINPUT29), .A3(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G2090), .ZN(new_n792));
  OAI21_X1  g367(.A(KEYINPUT29), .B1(new_n789), .B2(new_n790), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT98), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n685), .A2(G4), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n597), .B2(new_n685), .ZN(new_n797));
  INV_X1    g372(.A(G1348), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n791), .A2(new_n793), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n795), .B(new_n799), .C1(new_n792), .C2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(G28), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(KEYINPUT30), .ZN(new_n803));
  AOI21_X1  g378(.A(G29), .B1(new_n802), .B2(KEYINPUT30), .ZN(new_n804));
  OR2_X1    g379(.A1(KEYINPUT31), .A2(G11), .ZN(new_n805));
  NAND2_X1  g380(.A1(KEYINPUT31), .A2(G11), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n803), .A2(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n622), .B2(new_n747), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n747), .B1(KEYINPUT24), .B2(G34), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(KEYINPUT24), .B2(G34), .ZN(new_n810));
  INV_X1    g385(.A(G160), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(G29), .ZN(new_n812));
  INV_X1    g387(.A(G2084), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n808), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n813), .B2(new_n812), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n685), .A2(G21), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G168), .B2(new_n685), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT95), .B(G1966), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OAI22_X1  g394(.A1(new_n763), .A2(G2072), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  AOI211_X1 g395(.A(new_n815), .B(new_n820), .C1(new_n817), .C2(new_n819), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n685), .A2(G20), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT23), .Z(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(G299), .B2(G16), .ZN(new_n824));
  INV_X1    g399(.A(G1956), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(G164), .A2(new_n747), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(G27), .B2(new_n747), .ZN(new_n828));
  INV_X1    g403(.A(G2078), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n477), .A2(G128), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n481), .A2(G140), .ZN(new_n833));
  NOR2_X1   g408(.A1(G104), .A2(G2105), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(new_n468), .B2(G116), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n832), .B(new_n833), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G29), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n747), .A2(G26), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT28), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G2067), .ZN(new_n841));
  NOR4_X1   g416(.A1(new_n826), .A2(new_n830), .A3(new_n831), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n685), .A2(G19), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n551), .B2(new_n685), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(G1341), .Z(new_n845));
  NAND3_X1  g420(.A1(new_n821), .A2(new_n842), .A3(new_n845), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n788), .A2(new_n801), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n746), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(KEYINPUT87), .B(KEYINPUT36), .Z(new_n849));
  OAI21_X1  g424(.A(KEYINPUT86), .B1(new_n735), .B2(new_n736), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(new_n743), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n849), .B1(new_n851), .B2(new_n737), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n848), .A2(new_n852), .ZN(G311));
  NOR2_X1   g428(.A1(new_n740), .A2(new_n742), .ZN(new_n854));
  AOI211_X1 g429(.A(new_n854), .B(new_n705), .C1(new_n850), .C2(new_n743), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n746), .B(new_n847), .C1(new_n855), .C2(new_n849), .ZN(G150));
  NAND3_X1  g431(.A1(new_n523), .A2(G93), .A3(new_n512), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n528), .A2(G55), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(G80), .A2(G543), .ZN(new_n860));
  INV_X1    g435(.A(G67), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n541), .B2(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n862), .A2(KEYINPUT99), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n517), .B1(new_n862), .B2(KEYINPUT99), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n859), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G860), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT37), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT39), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n550), .A2(KEYINPUT100), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n544), .B(new_n871), .C1(new_n548), .C2(new_n549), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n865), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n865), .B1(new_n870), .B2(new_n872), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT38), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n870), .A2(new_n872), .ZN(new_n879));
  INV_X1    g454(.A(new_n865), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n873), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  NOR3_X1   g459(.A1(new_n884), .A2(new_n604), .A3(new_n607), .ZN(new_n885));
  AOI22_X1  g460(.A1(new_n878), .A2(new_n883), .B1(G559), .B2(new_n597), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n869), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n866), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n885), .A2(new_n869), .A3(new_n886), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n868), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n890), .B(new_n891), .ZN(G145));
  XOR2_X1   g467(.A(KEYINPUT104), .B(G37), .Z(new_n893));
  AOI22_X1  g468(.A1(new_n477), .A2(G130), .B1(G142), .B2(new_n481), .ZN(new_n894));
  OAI21_X1  g469(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n895));
  INV_X1    g470(.A(G118), .ZN(new_n896));
  AOI22_X1  g471(.A1(new_n895), .A2(KEYINPUT102), .B1(new_n896), .B2(G2105), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(KEYINPUT102), .B2(new_n895), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n612), .B(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n701), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n761), .B(new_n836), .Z(new_n903));
  XNOR2_X1  g478(.A(new_n780), .B(G164), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n904), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT105), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n811), .B(new_n622), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(G162), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n905), .A2(new_n902), .A3(new_n906), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n908), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n907), .A2(KEYINPUT105), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n893), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n905), .A2(new_n906), .ZN(new_n915));
  OR3_X1    g490(.A1(new_n915), .A2(KEYINPUT103), .A3(new_n901), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n911), .B1(new_n907), .B2(KEYINPUT103), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n910), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT40), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n919), .B(new_n920), .ZN(G395));
  OR2_X1    g496(.A1(new_n882), .A2(KEYINPUT106), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n882), .A2(KEYINPUT106), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n922), .A2(new_n608), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n608), .B1(new_n922), .B2(new_n923), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n592), .A2(G299), .A3(new_n596), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(G299), .B1(new_n592), .B2(new_n596), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT107), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n926), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT41), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(new_n928), .B2(new_n929), .ZN(new_n934));
  INV_X1    g509(.A(new_n929), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n935), .A2(KEYINPUT41), .A3(new_n927), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n934), .A2(new_n936), .A3(KEYINPUT108), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n930), .A2(new_n938), .A3(KEYINPUT41), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(new_n924), .B2(new_n925), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n588), .A2(new_n517), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n586), .B1(new_n530), .B2(new_n587), .ZN(new_n943));
  OR3_X1    g518(.A1(new_n942), .A2(new_n943), .A3(G288), .ZN(new_n944));
  NAND2_X1  g519(.A1(G290), .A2(G288), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(G303), .B(G305), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n946), .B1(new_n944), .B2(new_n945), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n948), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n954), .B(KEYINPUT42), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n932), .A2(new_n941), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n955), .B1(new_n932), .B2(new_n941), .ZN(new_n957));
  OAI21_X1  g532(.A(G868), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(G868), .B2(new_n865), .ZN(G295));
  OAI21_X1  g534(.A(new_n958), .B1(G868), .B2(new_n865), .ZN(G331));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n961));
  INV_X1    g536(.A(new_n930), .ZN(new_n962));
  OAI21_X1  g537(.A(G168), .B1(new_n874), .B2(new_n875), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n881), .A2(G286), .A3(new_n873), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(new_n964), .A3(G171), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(G171), .B1(new_n963), .B2(new_n964), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n962), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n874), .A2(new_n875), .A3(G168), .ZN(new_n969));
  AOI21_X1  g544(.A(G286), .B1(new_n881), .B2(new_n873), .ZN(new_n970));
  OAI21_X1  g545(.A(G301), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n971), .A2(new_n937), .A3(new_n939), .A4(new_n965), .ZN(new_n972));
  INV_X1    g547(.A(new_n954), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n968), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G37), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n973), .B1(new_n968), .B2(new_n972), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n961), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n931), .B1(new_n966), .B2(new_n967), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n971), .A2(new_n936), .A3(new_n934), .A4(new_n965), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(new_n980), .A3(new_n954), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n981), .A2(new_n974), .A3(KEYINPUT43), .A4(new_n893), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n978), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT44), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT43), .B1(new_n976), .B2(new_n977), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n981), .A2(new_n974), .A3(new_n961), .A4(new_n893), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n984), .A2(new_n989), .ZN(G397));
  INV_X1    g565(.A(G1384), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n503), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT50), .ZN(new_n993));
  XNOR2_X1  g568(.A(KEYINPUT110), .B(G40), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n467), .A2(new_n472), .A3(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n995), .B1(new_n503), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n993), .A2(new_n997), .A3(new_n813), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n467), .A2(new_n472), .A3(new_n994), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT4), .B1(new_n481), .B2(G138), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n500), .A2(new_n502), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1384), .B1(new_n1005), .B2(new_n496), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1001), .B(new_n1002), .C1(new_n1006), .C2(KEYINPUT45), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT45), .B1(new_n503), .B2(new_n991), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT114), .B1(new_n1008), .B2(new_n995), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(G1384), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n499), .A2(new_n500), .A3(new_n502), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n490), .A2(new_n495), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1007), .A2(new_n1009), .A3(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1015), .A2(KEYINPUT115), .A3(new_n818), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT115), .B1(new_n1015), .B2(new_n818), .ZN(new_n1017));
  OAI211_X1 g592(.A(G168), .B(new_n1000), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT123), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(new_n1019), .A3(G8), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n1020), .A2(KEYINPUT51), .ZN(new_n1021));
  NOR2_X1   g596(.A1(KEYINPUT123), .A2(KEYINPUT51), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1000), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1022), .B1(new_n1023), .B2(G286), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1018), .A2(G8), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT62), .B1(new_n1021), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1020), .A2(KEYINPUT51), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT62), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1028), .B(new_n1029), .C1(new_n1025), .C2(new_n1024), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1002), .A2(new_n991), .A3(new_n503), .ZN(new_n1031));
  OAI21_X1  g606(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1032), .A2(G1976), .A3(new_n575), .A4(new_n574), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n1033), .A3(G8), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT52), .ZN(new_n1035));
  INV_X1    g610(.A(G1976), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT52), .B1(G288), .B2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1037), .A2(G8), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n581), .A2(new_n584), .A3(new_n732), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n517), .B1(new_n578), .B2(new_n579), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n582), .A2(new_n583), .ZN(new_n1043));
  OAI21_X1  g618(.A(G1981), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT49), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1040), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1041), .A2(new_n1044), .A3(KEYINPUT113), .A4(KEYINPUT49), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1031), .A2(G8), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1050), .B1(new_n1046), .B2(new_n1045), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1039), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n1053));
  NAND3_X1  g628(.A1(G303), .A2(new_n1053), .A3(G8), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1053), .B1(G303), .B2(G8), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G8), .ZN(new_n1058));
  INV_X1    g633(.A(G1971), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1014), .A2(new_n1002), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1059), .B1(new_n1060), .B2(new_n1008), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n993), .A2(new_n997), .A3(new_n792), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1058), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OR2_X1    g638(.A1(new_n1057), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(KEYINPUT112), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT112), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n993), .A2(new_n997), .A3(new_n1066), .A4(new_n792), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1065), .A2(new_n1067), .A3(new_n1061), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1068), .A2(G8), .A3(new_n1057), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1052), .A2(new_n1064), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT125), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n992), .A2(new_n1010), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n995), .B1(new_n503), .B2(new_n1011), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1072), .A2(new_n1073), .A3(new_n829), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n993), .A2(new_n997), .ZN(new_n1076));
  INV_X1    g651(.A(G1961), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1074), .A2(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1075), .A2(G2078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1007), .A2(new_n1009), .A3(new_n1014), .A4(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT125), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1052), .A2(new_n1064), .A3(new_n1069), .A4(new_n1082), .ZN(new_n1083));
  AND4_X1   g658(.A1(G171), .A2(new_n1071), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1027), .A2(new_n1030), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n503), .A2(new_n996), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n1002), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT50), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1089), .B1(new_n503), .B2(new_n991), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n798), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G2067), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1006), .A2(new_n1092), .A3(new_n1002), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1091), .A2(KEYINPUT60), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT60), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1094), .B1(new_n1095), .B2(new_n607), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n597), .A2(KEYINPUT60), .A3(new_n1093), .A4(new_n1091), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1060), .A2(new_n1008), .A3(G1996), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT58), .B(G1341), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1100), .B1(new_n1006), .B2(new_n1002), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n551), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n551), .B(new_n1103), .C1(new_n1099), .C2(new_n1101), .ZN(new_n1106));
  NAND2_X1  g681(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n570), .B2(KEYINPUT118), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1111), .B(KEYINPUT57), .C1(new_n566), .C2(new_n569), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT56), .B(G2072), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1060), .A2(new_n1008), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(G1956), .B1(new_n993), .B2(new_n997), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1113), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n825), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1072), .A2(new_n1073), .A3(new_n1114), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1119), .A2(new_n1120), .A3(new_n1110), .A4(new_n1112), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1118), .A2(KEYINPUT61), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1098), .A2(new_n1108), .A3(new_n1122), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1119), .A2(new_n1120), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT61), .B1(new_n1124), .B2(KEYINPUT120), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT120), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1118), .A2(new_n1126), .A3(new_n1121), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1125), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1128), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1123), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1118), .B1(new_n1132), .B2(new_n607), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n1121), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1086), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1028), .B1(new_n1025), .B2(new_n1024), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1130), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1125), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g715(.A(KEYINPUT122), .B(new_n1134), .C1(new_n1140), .C2(new_n1123), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1081), .A2(G171), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1079), .A2(G40), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1072), .A2(G160), .A3(new_n1014), .A4(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1143), .A2(new_n1144), .A3(G301), .A4(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT124), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1078), .A2(new_n1149), .A3(G301), .A4(new_n1146), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1142), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT54), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1143), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT126), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1078), .A2(KEYINPUT126), .A3(new_n1146), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(G171), .A3(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1078), .A2(G301), .A3(new_n1080), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1158), .A2(KEYINPUT54), .A3(new_n1159), .ZN(new_n1160));
  AND4_X1   g735(.A1(new_n1071), .A2(new_n1153), .A3(new_n1083), .A4(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1136), .A2(new_n1137), .A3(new_n1141), .A4(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1163));
  NOR2_X1   g738(.A1(G288), .A2(G1976), .ZN(new_n1164));
  AOI22_X1  g739(.A1(new_n1163), .A2(new_n1164), .B1(new_n732), .B2(new_n724), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1039), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  OAI22_X1  g742(.A1(new_n1165), .A2(new_n1050), .B1(new_n1069), .B2(new_n1167), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n1052), .A2(new_n1069), .A3(KEYINPUT63), .ZN(new_n1169));
  NOR2_X1   g744(.A1(G286), .A2(new_n1058), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1068), .A2(G8), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1171), .B1(new_n1056), .B2(new_n1055), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1169), .A2(new_n1023), .A3(new_n1170), .A4(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT117), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1057), .A2(new_n1063), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1167), .A2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1176), .A2(new_n1023), .A3(new_n1069), .A4(new_n1170), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT63), .ZN(new_n1178));
  AOI22_X1  g753(.A1(new_n1173), .A2(new_n1174), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n1023), .A2(new_n1170), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1180), .A2(KEYINPUT117), .A3(new_n1172), .A4(new_n1169), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1168), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1085), .A2(new_n1162), .A3(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1072), .A2(new_n995), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1184), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1185), .A2(G1986), .A3(G290), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1184), .A2(G1986), .A3(G290), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1189), .B(KEYINPUT111), .Z(new_n1190));
  XNOR2_X1  g765(.A(new_n836), .B(G2067), .ZN(new_n1191));
  INV_X1    g766(.A(G1996), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n780), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n777), .A2(G1996), .A3(new_n779), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1191), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n701), .B(new_n703), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1185), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1190), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1183), .A2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g774(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1197), .B1(new_n1187), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1201), .B1(new_n1187), .B2(new_n1200), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT46), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1203), .B1(new_n1185), .B2(G1996), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1184), .A2(KEYINPUT46), .A3(new_n1192), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1184), .B1(new_n1191), .B2(new_n780), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1207), .B(KEYINPUT47), .ZN(new_n1208));
  INV_X1    g783(.A(new_n703), .ZN(new_n1209));
  NOR2_X1   g784(.A1(new_n701), .A2(new_n1209), .ZN(new_n1210));
  AND2_X1   g785(.A1(new_n1195), .A2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n836), .A2(G2067), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1184), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  AND3_X1   g788(.A1(new_n1202), .A2(new_n1208), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1199), .A2(new_n1214), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g790(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1217));
  AND3_X1   g791(.A1(new_n1217), .A2(new_n679), .A3(new_n680), .ZN(new_n1218));
  OAI21_X1  g792(.A(new_n1218), .B1(new_n914), .B2(new_n918), .ZN(new_n1219));
  AOI21_X1  g793(.A(new_n1219), .B1(new_n985), .B2(new_n986), .ZN(G308));
  OAI211_X1 g794(.A(new_n987), .B(new_n1218), .C1(new_n918), .C2(new_n914), .ZN(G225));
endmodule


