//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n810, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g002(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT27), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT27), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n206), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n207));
  INV_X1    g006(.A(G190gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT67), .ZN(new_n210));
  AOI21_X1  g009(.A(G190gat), .B1(new_n204), .B2(KEYINPUT27), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT67), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(new_n212), .A3(new_n207), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT28), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT28), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT27), .B(G183gat), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(new_n208), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT68), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n211), .A2(new_n212), .A3(new_n207), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n212), .B1(new_n211), .B2(new_n207), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n215), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT68), .ZN(new_n222));
  INV_X1    g021(.A(new_n217), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NOR3_X1   g027(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n225), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n230), .B(KEYINPUT69), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n218), .A2(new_n224), .A3(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n233));
  NOR2_X1   g032(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n234));
  OAI22_X1  g033(.A1(new_n233), .A2(new_n234), .B1(G169gat), .B2(G176gat), .ZN(new_n235));
  INV_X1    g034(.A(G169gat), .ZN(new_n236));
  INV_X1    g035(.A(G176gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n235), .B(new_n227), .C1(new_n238), .C2(new_n234), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT25), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT24), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G183gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(new_n208), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n246), .B1(new_n242), .B2(new_n225), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n241), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n243), .A2(KEYINPUT64), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n243), .A2(KEYINPUT64), .ZN(new_n250));
  NOR3_X1   g049(.A1(new_n249), .A2(new_n250), .A3(new_n247), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n240), .B1(new_n251), .B2(new_n239), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G113gat), .B(G120gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT71), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G113gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n257), .A2(G120gat), .ZN(new_n258));
  INV_X1    g057(.A(G120gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n259), .A2(G113gat), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT71), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G134gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G127gat), .ZN(new_n263));
  INV_X1    g062(.A(G127gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G134gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT1), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n263), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n256), .A2(new_n261), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT70), .B1(new_n264), .B2(G134gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n265), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n263), .A2(KEYINPUT70), .ZN(new_n271));
  OAI22_X1  g070(.A1(new_n270), .A2(new_n271), .B1(new_n254), .B2(KEYINPUT1), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n232), .A2(new_n253), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n273), .B1(new_n232), .B2(new_n253), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n203), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT32), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT33), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G15gat), .B(G43gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(G71gat), .B(G99gat), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n280), .B(new_n281), .Z(new_n282));
  NAND3_X1  g081(.A1(new_n277), .A2(new_n279), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n282), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n276), .B(KEYINPUT32), .C1(new_n278), .C2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n232), .A2(new_n253), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n268), .A2(new_n272), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n232), .A2(new_n253), .A3(new_n273), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT34), .B1(new_n291), .B2(new_n203), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n274), .A2(new_n275), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT34), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n293), .A2(new_n294), .A3(new_n295), .A4(new_n202), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n289), .A2(new_n295), .A3(new_n202), .A4(new_n290), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT73), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n292), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT74), .B1(new_n286), .B2(new_n299), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n292), .A2(new_n296), .A3(new_n298), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n301), .A2(new_n302), .A3(new_n285), .A4(new_n283), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n305));
  XNOR2_X1  g104(.A(G197gat), .B(G204gat), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n307), .A2(KEYINPUT75), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(KEYINPUT75), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n306), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(G211gat), .B(G218gat), .Z(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n305), .B1(new_n313), .B2(KEYINPUT29), .ZN(new_n314));
  NAND2_X1  g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315));
  INV_X1    g114(.A(G155gat), .ZN(new_n316));
  INV_X1    g115(.A(G162gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n315), .B1(new_n318), .B2(KEYINPUT2), .ZN(new_n319));
  INV_X1    g118(.A(G148gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G141gat), .ZN(new_n321));
  INV_X1    g120(.A(G141gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(G148gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  OR2_X1    g124(.A1(KEYINPUT81), .A2(KEYINPUT2), .ZN(new_n326));
  NAND2_X1  g125(.A1(KEYINPUT81), .A2(KEYINPUT2), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n321), .A2(new_n323), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n318), .A2(new_n315), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n326), .A2(new_n327), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n324), .ZN(new_n333));
  INV_X1    g132(.A(new_n329), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n333), .A2(new_n334), .B1(new_n319), .B2(new_n324), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT29), .B1(new_n335), .B2(new_n305), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n312), .A2(new_n336), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n337), .A2(KEYINPUT87), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(KEYINPUT87), .ZN(new_n339));
  NAND2_X1  g138(.A1(G228gat), .A2(G233gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n331), .A2(new_n338), .A3(new_n339), .A4(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT29), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n310), .A2(KEYINPUT86), .A3(new_n311), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n343), .B(new_n344), .C1(new_n312), .C2(KEYINPUT86), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(new_n305), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n337), .B1(new_n346), .B2(new_n330), .ZN(new_n347));
  XOR2_X1   g146(.A(new_n340), .B(KEYINPUT85), .Z(new_n348));
  OAI21_X1  g147(.A(new_n342), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G78gat), .B(G106gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n350), .B(G22gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT31), .B(G50gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n349), .B(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT72), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n286), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n283), .A2(KEYINPUT72), .A3(new_n285), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n299), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n304), .A2(new_n355), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT76), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n363), .B1(new_n287), .B2(new_n343), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n361), .B1(new_n232), .B2(new_n253), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n313), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n287), .A2(new_n363), .ZN(new_n367));
  INV_X1    g166(.A(new_n361), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT29), .B1(new_n232), .B2(new_n253), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n367), .B(new_n312), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G8gat), .B(G36gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(G92gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT77), .B(G64gat), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n373), .B(new_n374), .Z(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n371), .A2(KEYINPUT78), .A3(KEYINPUT30), .A4(new_n376), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n366), .A2(KEYINPUT30), .A3(new_n370), .A4(new_n376), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n376), .B1(new_n366), .B2(new_n370), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT78), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT79), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n377), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n366), .A2(new_n370), .A3(new_n376), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT30), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT80), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT80), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n386), .A2(new_n390), .A3(new_n387), .ZN(new_n391));
  XOR2_X1   g190(.A(G57gat), .B(G85gat), .Z(new_n392));
  XNOR2_X1  g191(.A(G1gat), .B(G29gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT5), .ZN(new_n398));
  NAND2_X1  g197(.A1(G225gat), .A2(G233gat), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n399), .B(KEYINPUT82), .Z(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n335), .A2(new_n305), .B1(new_n268), .B2(new_n272), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n330), .A2(KEYINPUT3), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT4), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n273), .B2(new_n335), .ZN(new_n406));
  NOR3_X1   g205(.A1(new_n288), .A2(new_n330), .A3(KEYINPUT4), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n401), .B(new_n404), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n273), .A2(new_n335), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n288), .A2(new_n330), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n400), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n398), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n273), .A2(new_n405), .A3(new_n335), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT4), .B1(new_n288), .B2(new_n330), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n413), .A2(new_n414), .B1(new_n402), .B2(new_n403), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT5), .B1(new_n415), .B2(new_n401), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n397), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT84), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n412), .A2(new_n416), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n396), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT6), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT84), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n422), .B(new_n397), .C1(new_n412), .C2(new_n416), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n418), .A2(new_n420), .A3(new_n421), .A4(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n419), .A2(KEYINPUT6), .A3(new_n396), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n389), .A2(new_n391), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n383), .A2(new_n385), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT35), .B1(new_n360), .B2(new_n427), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n386), .A2(new_n390), .A3(new_n387), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n390), .B1(new_n386), .B2(new_n387), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n381), .B(new_n377), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n425), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n418), .A2(new_n421), .A3(new_n423), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n419), .A2(KEYINPUT88), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT88), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n412), .A2(new_n416), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n396), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n432), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT89), .B(KEYINPUT35), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n431), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n300), .A2(new_n303), .B1(new_n286), .B2(new_n299), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n355), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n428), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n354), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n304), .A2(new_n359), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT36), .ZN(new_n446));
  OR3_X1    g245(.A1(new_n409), .A2(new_n400), .A3(new_n410), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n447), .B(KEYINPUT39), .C1(new_n401), .C2(new_n415), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n415), .A2(new_n401), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n448), .B(new_n397), .C1(KEYINPUT39), .C2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT40), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OR2_X1    g251(.A1(new_n450), .A2(new_n451), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n437), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n431), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n366), .A2(new_n370), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT37), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT37), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n366), .A2(new_n458), .A3(new_n370), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT38), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n376), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n457), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n312), .B1(new_n364), .B2(new_n365), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n367), .B(new_n313), .C1(new_n368), .C2(new_n369), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(KEYINPUT37), .A3(new_n464), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n459), .A2(new_n465), .A3(new_n375), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n386), .A2(new_n460), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n438), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n455), .A2(new_n469), .A3(new_n355), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT36), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n441), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n444), .A2(new_n446), .A3(new_n470), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n443), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT90), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT90), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n443), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(G43gat), .B(G50gat), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT15), .ZN(new_n480));
  INV_X1    g279(.A(G29gat), .ZN(new_n481));
  INV_X1    g280(.A(G36gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT14), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n485), .A2(new_n481), .A3(new_n482), .ZN(new_n486));
  AOI211_X1 g285(.A(new_n480), .B(new_n483), .C1(new_n484), .C2(new_n486), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n486), .A2(new_n484), .B1(G29gat), .B2(G36gat), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n479), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n491));
  INV_X1    g290(.A(new_n479), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT17), .ZN(new_n495));
  XNOR2_X1  g294(.A(G15gat), .B(G22gat), .ZN(new_n496));
  INV_X1    g295(.A(G1gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT16), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(G1gat), .B2(new_n496), .ZN(new_n500));
  XOR2_X1   g299(.A(new_n500), .B(G8gat), .Z(new_n501));
  INV_X1    g300(.A(KEYINPUT17), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n490), .A2(new_n502), .A3(new_n493), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n495), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n501), .A2(new_n494), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT92), .ZN(new_n507));
  NAND2_X1  g306(.A1(G229gat), .A2(G233gat), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT18), .A4(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT91), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT18), .A4(new_n508), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT92), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n501), .A2(new_n494), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n505), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n508), .B(KEYINPUT13), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n509), .A2(new_n510), .A3(new_n512), .A4(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G113gat), .B(G141gat), .ZN(new_n519));
  INV_X1    g318(.A(G197gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT11), .B(G169gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT12), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n518), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n504), .A2(new_n505), .A3(new_n508), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT18), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n509), .A2(new_n529), .A3(new_n512), .A4(new_n517), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n518), .A3(new_n525), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT97), .ZN(new_n535));
  XNOR2_X1  g334(.A(G134gat), .B(G162gat), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n536), .B(new_n537), .Z(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(G99gat), .A2(G106gat), .ZN(new_n541));
  INV_X1    g340(.A(G85gat), .ZN(new_n542));
  INV_X1    g341(.A(G92gat), .ZN(new_n543));
  AOI22_X1  g342(.A1(KEYINPUT8), .A2(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT7), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(new_n542), .B2(new_n543), .ZN(new_n546));
  NAND3_X1  g345(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G99gat), .B(G106gat), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n548), .B(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n540), .B1(new_n494), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT96), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n495), .A2(new_n503), .A3(new_n551), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G190gat), .B(G218gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT95), .ZN(new_n558));
  AOI211_X1 g357(.A(new_n535), .B(new_n539), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n558), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT97), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n538), .B1(new_n557), .B2(new_n535), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n559), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OR2_X1    g362(.A1(G57gat), .A2(G64gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(G57gat), .A2(G64gat), .ZN(new_n565));
  AND2_X1   g364(.A1(G71gat), .A2(G78gat), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n564), .B(new_n565), .C1(new_n566), .C2(KEYINPUT9), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n566), .A2(KEYINPUT93), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(G71gat), .A2(G78gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n567), .B(new_n568), .C1(new_n566), .C2(new_n570), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT21), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n501), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G127gat), .B(G155gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT20), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n578), .B(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n574), .A2(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(new_n245), .ZN(new_n584));
  INV_X1    g383(.A(G211gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n582), .B(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n581), .B(new_n587), .Z(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n563), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n551), .A2(new_n572), .A3(new_n573), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n548), .B(new_n549), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(new_n574), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT98), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(G230gat), .ZN(new_n596));
  INV_X1    g395(.A(G233gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n551), .A2(KEYINPUT98), .A3(new_n572), .A4(new_n573), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n595), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n600), .A2(KEYINPUT100), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT101), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT10), .B1(new_n595), .B2(new_n599), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT10), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n593), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT99), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  OR2_X1    g405(.A1(new_n605), .A2(KEYINPUT99), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n598), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n600), .A2(KEYINPUT100), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n601), .B(new_n602), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G120gat), .B(G148gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(G176gat), .B(G204gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n610), .A2(new_n614), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n590), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n478), .A2(new_n534), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n424), .A2(new_n425), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(new_n497), .ZN(G1324gat));
  INV_X1    g422(.A(new_n431), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT102), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT102), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n627), .B1(new_n620), .B2(new_n624), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT16), .B(G8gat), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT42), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n629), .A2(G8gat), .B1(new_n625), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n631), .B1(new_n629), .B2(new_n630), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(G1325gat));
  INV_X1    g434(.A(G15gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n446), .A2(new_n472), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n620), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n478), .A2(new_n534), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n640), .A2(new_n441), .A3(new_n619), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n639), .B1(new_n641), .B2(new_n636), .ZN(G1326gat));
  NOR2_X1   g441(.A1(new_n620), .A2(new_n355), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT43), .B(G22gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(G1327gat));
  INV_X1    g444(.A(new_n617), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n646), .A2(new_n588), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n563), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n478), .A2(new_n534), .A3(new_n650), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n651), .A2(G29gat), .A3(new_n621), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n652), .B(KEYINPUT45), .Z(new_n653));
  NAND3_X1  g452(.A1(new_n475), .A2(new_n477), .A3(new_n563), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT44), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n428), .A2(KEYINPUT104), .A3(new_n442), .ZN(new_n656));
  AOI21_X1  g455(.A(KEYINPUT104), .B1(new_n428), .B2(new_n442), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n473), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n563), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT103), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n530), .A2(new_n518), .A3(new_n525), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n530), .B1(new_n518), .B2(new_n525), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n532), .A2(KEYINPUT103), .A3(new_n533), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n648), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n661), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(G29gat), .B1(new_n669), .B2(new_n621), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n653), .A2(new_n670), .ZN(G1328gat));
  NOR2_X1   g470(.A1(new_n624), .A2(G36gat), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n640), .A2(KEYINPUT106), .A3(new_n650), .A4(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT46), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n675));
  INV_X1    g474(.A(new_n672), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n675), .B1(new_n651), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n673), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(G36gat), .B1(new_n669), .B2(new_n624), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n673), .A2(new_n677), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n680), .B1(new_n681), .B2(KEYINPUT46), .ZN(new_n682));
  AOI211_X1 g481(.A(KEYINPUT107), .B(new_n674), .C1(new_n673), .C2(new_n677), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n678), .B(new_n679), .C1(new_n682), .C2(new_n683), .ZN(G1329gat));
  OAI21_X1  g483(.A(G43gat), .B1(new_n669), .B2(new_n638), .ZN(new_n685));
  INV_X1    g484(.A(new_n441), .ZN(new_n686));
  OR3_X1    g485(.A1(new_n651), .A2(G43gat), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT47), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n685), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n688), .B1(new_n685), .B2(new_n687), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(G1330gat));
  NAND2_X1  g490(.A1(new_n354), .A2(G50gat), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n651), .A2(new_n355), .ZN(new_n693));
  OAI22_X1  g492(.A1(new_n669), .A2(new_n692), .B1(new_n693), .B2(G50gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1331gat));
  NAND3_X1  g495(.A1(new_n590), .A2(new_n646), .A3(new_n667), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n658), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n621), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g502(.A1(new_n699), .A2(new_n624), .ZN(new_n704));
  NOR2_X1   g503(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n705));
  AND2_X1   g504(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(new_n704), .B2(new_n705), .ZN(G1333gat));
  INV_X1    g507(.A(G71gat), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n700), .B2(new_n637), .ZN(new_n710));
  OR3_X1    g509(.A1(new_n699), .A2(KEYINPUT109), .A3(new_n686), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT109), .B1(new_n699), .B2(new_n686), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n710), .B1(new_n713), .B2(new_n709), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n354), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(G78gat), .ZN(G1335gat));
  INV_X1    g516(.A(new_n667), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(new_n588), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n658), .A2(new_n563), .A3(new_n719), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n720), .A2(KEYINPUT51), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n617), .B1(new_n720), .B2(KEYINPUT51), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n724), .A2(new_n542), .A3(new_n701), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n719), .A2(new_n646), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n726), .B1(new_n655), .B2(new_n660), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(KEYINPUT110), .A3(new_n701), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G85gat), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT110), .B1(new_n727), .B2(new_n701), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n725), .B1(new_n729), .B2(new_n730), .ZN(G1336gat));
  INV_X1    g530(.A(new_n726), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n661), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT111), .B1(new_n733), .B2(new_n624), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT111), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n727), .A2(new_n735), .A3(new_n431), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n734), .A2(G92gat), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n624), .A2(G92gat), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT52), .B1(new_n724), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n723), .A2(G92gat), .A3(new_n624), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n543), .B1(new_n727), .B2(new_n431), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT52), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n743), .ZN(G1337gat));
  AOI21_X1  g543(.A(G99gat), .B1(new_n724), .B2(new_n441), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n727), .A2(G99gat), .A3(new_n637), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(G1338gat));
  INV_X1    g546(.A(G106gat), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n721), .A2(new_n722), .A3(new_n748), .A4(new_n354), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n748), .B1(new_n727), .B2(new_n354), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT112), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AOI211_X1 g551(.A(KEYINPUT112), .B(new_n748), .C1(new_n727), .C2(new_n354), .ZN(new_n753));
  OAI21_X1  g552(.A(KEYINPUT53), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n749), .A2(KEYINPUT113), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n750), .A2(KEYINPUT53), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n749), .A2(KEYINPUT113), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n754), .A2(new_n758), .ZN(G1339gat));
  NAND3_X1  g558(.A1(new_n590), .A2(new_n617), .A3(new_n667), .ZN(new_n760));
  INV_X1    g559(.A(new_n559), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n561), .A2(new_n562), .ZN(new_n762));
  OR3_X1    g561(.A1(new_n506), .A2(KEYINPUT115), .A3(new_n508), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n505), .A2(new_n513), .A3(new_n515), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT116), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT115), .B1(new_n506), .B2(new_n508), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n763), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n531), .A2(new_n524), .B1(new_n767), .B2(new_n523), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n761), .A2(new_n762), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n606), .A2(new_n607), .ZN(new_n770));
  INV_X1    g569(.A(new_n598), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n606), .A2(new_n598), .A3(new_n607), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n772), .A2(KEYINPUT54), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n614), .B1(new_n608), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n774), .A2(KEYINPUT55), .A3(new_n776), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n601), .B1(new_n608), .B2(new_n609), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n614), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n779), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n769), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n768), .B1(new_n615), .B2(new_n616), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n667), .B2(new_n783), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n563), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n785), .B(KEYINPUT117), .C1(new_n667), .C2(new_n783), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n784), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n760), .B1(new_n790), .B2(new_n588), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n431), .A2(new_n621), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n686), .A2(new_n354), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n534), .ZN(new_n796));
  OAI21_X1  g595(.A(G113gat), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n360), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n718), .A2(new_n257), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n797), .B1(new_n799), .B2(new_n800), .ZN(G1340gat));
  INV_X1    g600(.A(new_n799), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(new_n259), .A3(new_n646), .ZN(new_n803));
  OAI21_X1  g602(.A(G120gat), .B1(new_n795), .B2(new_n617), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n803), .A2(KEYINPUT118), .A3(new_n804), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(G1341gat));
  NOR3_X1   g608(.A1(new_n795), .A2(new_n264), .A3(new_n589), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n802), .A2(new_n588), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n810), .B1(new_n264), .B2(new_n811), .ZN(G1342gat));
  NAND2_X1  g611(.A1(new_n563), .A2(new_n262), .ZN(new_n813));
  OR3_X1    g612(.A1(new_n799), .A2(KEYINPUT56), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n786), .A2(new_n787), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n815), .A2(new_n649), .A3(new_n789), .ZN(new_n816));
  INV_X1    g615(.A(new_n784), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n588), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n760), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR4_X1   g619(.A1(new_n820), .A2(new_n621), .A3(new_n431), .A4(new_n649), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n794), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G134gat), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT56), .B1(new_n799), .B2(new_n813), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n814), .A2(new_n823), .A3(new_n824), .ZN(G1343gat));
  NOR2_X1   g624(.A1(new_n820), .A2(new_n355), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n638), .A2(new_n792), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  AND4_X1   g627(.A1(new_n322), .A2(new_n826), .A3(new_n534), .A4(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(KEYINPUT58), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n791), .A2(new_n831), .A3(new_n354), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n534), .A2(new_n779), .A3(new_n780), .A4(new_n782), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n563), .B1(new_n785), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n589), .B1(new_n834), .B2(new_n784), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n760), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n354), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n827), .B1(new_n837), .B2(KEYINPUT57), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n832), .A2(new_n838), .A3(new_n534), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n839), .A2(KEYINPUT120), .ZN(new_n840));
  OAI21_X1  g639(.A(G141gat), .B1(new_n839), .B2(KEYINPUT120), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n830), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n832), .A2(new_n838), .A3(new_n718), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n843), .A2(KEYINPUT119), .A3(G141gat), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT119), .B1(new_n843), .B2(G141gat), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n844), .A2(new_n845), .A3(new_n829), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n842), .B1(new_n846), .B2(new_n847), .ZN(G1344gat));
  NAND2_X1  g647(.A1(new_n826), .A2(new_n828), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n320), .A3(new_n646), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n852));
  OAI211_X1 g651(.A(KEYINPUT57), .B(new_n354), .C1(new_n818), .C2(new_n819), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n791), .A2(KEYINPUT121), .A3(KEYINPUT57), .A4(new_n354), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n835), .B1(new_n534), .B2(new_n618), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT57), .B1(new_n857), .B2(new_n354), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n855), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n646), .A3(new_n828), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n852), .B1(new_n861), .B2(G148gat), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n832), .A2(new_n838), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n617), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n864), .A2(KEYINPUT59), .A3(new_n320), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n851), .B1(new_n862), .B2(new_n865), .ZN(G1345gat));
  NOR3_X1   g665(.A1(new_n863), .A2(new_n316), .A3(new_n589), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n588), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n868), .B2(new_n316), .ZN(G1346gat));
  NAND4_X1  g668(.A1(new_n821), .A2(new_n317), .A3(new_n354), .A4(new_n638), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n870), .A2(KEYINPUT122), .ZN(new_n871));
  OAI21_X1  g670(.A(G162gat), .B1(new_n863), .B2(new_n649), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(KEYINPUT122), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(G1347gat));
  NAND2_X1  g673(.A1(new_n798), .A2(new_n431), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n621), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n877), .B1(new_n876), .B2(new_n875), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n791), .A2(new_n236), .A3(new_n718), .A4(new_n878), .ZN(new_n879));
  XOR2_X1   g678(.A(new_n879), .B(KEYINPUT124), .Z(new_n880));
  NAND2_X1  g679(.A1(new_n431), .A2(new_n621), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n881), .B(KEYINPUT125), .Z(new_n882));
  AND2_X1   g681(.A1(new_n882), .A2(new_n794), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n791), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(G169gat), .B1(new_n884), .B2(new_n796), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT126), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n880), .A2(new_n885), .A3(KEYINPUT126), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(G1348gat));
  AND2_X1   g689(.A1(new_n791), .A2(new_n878), .ZN(new_n891));
  AOI21_X1  g690(.A(G176gat), .B1(new_n891), .B2(new_n646), .ZN(new_n892));
  INV_X1    g691(.A(new_n884), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n617), .A2(new_n237), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(G1349gat));
  NAND3_X1  g694(.A1(new_n891), .A2(new_n216), .A3(new_n588), .ZN(new_n896));
  OAI21_X1  g695(.A(G183gat), .B1(new_n884), .B2(new_n589), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g698(.A1(new_n891), .A2(new_n208), .A3(new_n563), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n791), .A2(new_n883), .A3(new_n563), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n901), .A2(new_n902), .A3(G190gat), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n901), .B2(G190gat), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT127), .ZN(G1351gat));
  NOR4_X1   g705(.A1(new_n820), .A2(new_n355), .A3(new_n637), .A4(new_n881), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n520), .A3(new_n718), .ZN(new_n908));
  INV_X1    g707(.A(new_n882), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(new_n637), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n858), .B1(new_n853), .B2(new_n854), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(new_n912), .B2(new_n856), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n913), .A2(new_n534), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n908), .B1(new_n914), .B2(new_n520), .ZN(G1352gat));
  INV_X1    g714(.A(G204gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n907), .A2(new_n916), .A3(new_n646), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n917), .A2(KEYINPUT62), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(KEYINPUT62), .ZN(new_n919));
  AOI211_X1 g718(.A(new_n617), .B(new_n911), .C1(new_n912), .C2(new_n856), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n918), .B(new_n919), .C1(new_n916), .C2(new_n920), .ZN(G1353gat));
  NAND3_X1  g720(.A1(new_n907), .A2(new_n585), .A3(new_n588), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n860), .A2(new_n588), .A3(new_n910), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n923), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT63), .B1(new_n923), .B2(G211gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(G1354gat));
  AOI21_X1  g725(.A(G218gat), .B1(new_n907), .B2(new_n563), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n563), .A2(G218gat), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n927), .B1(new_n913), .B2(new_n928), .ZN(G1355gat));
endmodule


