//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985;
  NOR2_X1   g000(.A1(G475), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G237), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  AND4_X1   g004(.A1(G143), .A2(new_n189), .A3(new_n190), .A4(G214), .ZN(new_n191));
  NOR2_X1   g005(.A1(G237), .A2(G953), .ZN(new_n192));
  AOI21_X1  g006(.A(G143), .B1(new_n192), .B2(G214), .ZN(new_n193));
  OAI21_X1  g007(.A(G131), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n189), .A2(new_n190), .A3(G214), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n192), .A2(G143), .A3(G214), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G125), .ZN(new_n201));
  NOR3_X1   g015(.A1(new_n201), .A2(KEYINPUT16), .A3(G140), .ZN(new_n202));
  XNOR2_X1  g016(.A(G125), .B(G140), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(KEYINPUT16), .ZN(new_n204));
  AOI22_X1  g018(.A1(new_n194), .A2(new_n200), .B1(new_n204), .B2(G146), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  INV_X1    g020(.A(G140), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n201), .A2(G140), .ZN(new_n209));
  AND3_X1   g023(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT19), .ZN(new_n210));
  AOI21_X1  g024(.A(KEYINPUT19), .B1(new_n208), .B2(new_n209), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n206), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT87), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT87), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n214), .B(new_n206), .C1(new_n210), .C2(new_n211), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n205), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n203), .B(new_n206), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT18), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n197), .B(new_n199), .C1(new_n218), .C2(new_n198), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n217), .B(new_n219), .C1(new_n218), .C2(new_n194), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT88), .ZN(new_n222));
  XNOR2_X1  g036(.A(G113), .B(G122), .ZN(new_n223));
  INV_X1    g037(.A(G104), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n223), .B(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT88), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n216), .A2(new_n220), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n222), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  OR2_X1    g043(.A1(new_n204), .A2(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n204), .A2(G146), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n194), .A2(new_n200), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n230), .B(new_n231), .C1(KEYINPUT17), .C2(new_n232), .ZN(new_n233));
  OAI211_X1 g047(.A(KEYINPUT17), .B(G131), .C1(new_n191), .C2(new_n193), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n234), .B(KEYINPUT89), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n225), .B(new_n220), .C1(new_n233), .C2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n188), .B1(new_n229), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT20), .ZN(new_n238));
  OAI21_X1  g052(.A(KEYINPUT90), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n228), .A2(new_n226), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n227), .B1(new_n216), .B2(new_n220), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n236), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n187), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT90), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(new_n244), .A3(KEYINPUT20), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n237), .A2(new_n238), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n239), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G902), .ZN(new_n248));
  OR2_X1    g062(.A1(new_n233), .A2(new_n235), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n225), .B1(new_n249), .B2(new_n220), .ZN(new_n250));
  INV_X1    g064(.A(new_n236), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G475), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n247), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G478), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(KEYINPUT15), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n196), .A2(G128), .ZN(new_n258));
  INV_X1    g072(.A(G128), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G143), .ZN(new_n260));
  INV_X1    g074(.A(G134), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G116), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G122), .ZN(new_n264));
  INV_X1    g078(.A(G122), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G116), .ZN(new_n266));
  INV_X1    g080(.A(G107), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n267), .B1(new_n264), .B2(new_n266), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n262), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n196), .A2(G128), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT13), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n258), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n259), .A2(G143), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT13), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n261), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(G134), .B1(new_n274), .B2(new_n271), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n268), .B1(new_n262), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT91), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n281), .B(KEYINPUT14), .C1(new_n265), .C2(G116), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT14), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(new_n263), .A3(G122), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n266), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n281), .B1(new_n264), .B2(KEYINPUT14), .ZN(new_n286));
  OAI21_X1  g100(.A(G107), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n280), .A2(new_n287), .A3(KEYINPUT92), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT92), .B1(new_n280), .B2(new_n287), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n278), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  XOR2_X1   g105(.A(KEYINPUT9), .B(G234), .Z(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(G217), .A3(new_n190), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n280), .A2(new_n287), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT92), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n288), .ZN(new_n298));
  INV_X1    g112(.A(new_n293), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n278), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n248), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n257), .B1(new_n302), .B2(KEYINPUT93), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(KEYINPUT93), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n303), .B(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  XOR2_X1   g120(.A(KEYINPUT21), .B(G898), .Z(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(KEYINPUT94), .ZN(new_n308));
  AOI211_X1 g122(.A(new_n248), .B(new_n190), .C1(G234), .C2(G237), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G952), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n312), .A2(G953), .ZN(new_n313));
  INV_X1    g127(.A(G234), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n313), .B1(new_n314), .B2(new_n189), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(KEYINPUT95), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n255), .A2(new_n306), .A3(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(G214), .B1(G237), .B2(G902), .ZN(new_n320));
  XNOR2_X1  g134(.A(G110), .B(G122), .ZN(new_n321));
  INV_X1    g135(.A(G119), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT67), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT67), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G119), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT5), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n323), .A2(new_n325), .A3(new_n326), .A4(G116), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT82), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT67), .B(G119), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT82), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n329), .A2(new_n330), .A3(new_n326), .A4(G116), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G113), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n322), .A2(G116), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n334), .B1(new_n329), .B2(G116), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n333), .B1(new_n335), .B2(KEYINPUT5), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n323), .A2(new_n325), .A3(G116), .ZN(new_n337));
  INV_X1    g151(.A(new_n334), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n333), .A2(KEYINPUT2), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT2), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G113), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n337), .A2(new_n338), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT68), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT68), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n337), .A2(new_n342), .A3(new_n345), .A4(new_n338), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n332), .A2(new_n336), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT3), .B1(new_n224), .B2(G107), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT3), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n267), .A3(G104), .ZN(new_n350));
  INV_X1    g164(.A(G101), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n224), .A2(G107), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n348), .A2(new_n350), .A3(new_n351), .A4(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n224), .A2(G107), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n267), .A2(G104), .ZN(new_n355));
  OAI21_X1  g169(.A(G101), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT80), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n353), .A2(new_n356), .A3(KEYINPUT80), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n347), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n344), .A2(new_n346), .ZN(new_n363));
  INV_X1    g177(.A(new_n335), .ZN(new_n364));
  INV_X1    g178(.A(new_n342), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n348), .A2(new_n350), .A3(new_n352), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n368), .A2(new_n369), .A3(G101), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n369), .B1(new_n368), .B2(G101), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n370), .B1(new_n353), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n321), .B1(new_n362), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(KEYINPUT6), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n337), .A2(KEYINPUT5), .A3(new_n338), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n377), .A2(new_n328), .A3(new_n331), .A4(G113), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n363), .A2(new_n378), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n353), .A2(new_n356), .A3(KEYINPUT80), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT80), .B1(new_n353), .B2(new_n356), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n344), .A2(new_n346), .B1(new_n364), .B2(new_n365), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n368), .A2(G101), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(KEYINPUT4), .A3(new_n353), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n368), .A2(new_n369), .A3(G101), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI22_X1  g201(.A1(new_n379), .A2(new_n382), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n321), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT83), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT83), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n362), .A2(new_n373), .A3(new_n391), .A4(new_n321), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n374), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT6), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n376), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT64), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT0), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(new_n259), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n206), .A2(G143), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n196), .A2(G146), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(KEYINPUT0), .A2(G128), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n400), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT65), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT65), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n400), .A2(new_n407), .A3(new_n403), .A4(new_n404), .ZN(new_n408));
  OR2_X1    g222(.A1(new_n403), .A2(new_n404), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n406), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G125), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n401), .A2(KEYINPUT1), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n403), .A2(new_n412), .A3(G128), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n401), .B(new_n402), .C1(KEYINPUT1), .C2(new_n259), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n201), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n190), .A2(G224), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n417), .B(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n395), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(G210), .B1(G237), .B2(G902), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n411), .A2(KEYINPUT7), .A3(new_n418), .A4(new_n416), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT86), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n416), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n415), .A2(KEYINPUT86), .A3(new_n201), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n425), .A2(new_n426), .B1(new_n410), .B2(G125), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n418), .A2(KEYINPUT7), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n423), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(new_n392), .B2(new_n390), .ZN(new_n430));
  XNOR2_X1  g244(.A(KEYINPUT84), .B(KEYINPUT8), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n321), .B(new_n431), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n379), .A2(new_n357), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT85), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n362), .B1(new_n433), .B2(new_n434), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n432), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(G902), .B1(new_n430), .B2(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n421), .A2(new_n422), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n422), .B1(new_n421), .B2(new_n438), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n320), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n319), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT26), .B(G101), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n192), .A2(G210), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n443), .B(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n446));
  XOR2_X1   g260(.A(new_n445), .B(new_n446), .Z(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n408), .A2(new_n409), .ZN(new_n449));
  NAND2_X1  g263(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n261), .A2(G137), .ZN(new_n452));
  OR2_X1    g266(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n261), .A2(G137), .ZN(new_n455));
  INV_X1    g269(.A(G137), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G134), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n455), .B1(new_n457), .B2(new_n450), .ZN(new_n458));
  OAI21_X1  g272(.A(G131), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n456), .A2(G134), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n460), .B1(new_n452), .B2(new_n451), .ZN(new_n461));
  NOR2_X1   g275(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n450), .B1(new_n457), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n461), .A2(new_n198), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n449), .A2(new_n465), .A3(new_n406), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n413), .A2(new_n414), .ZN(new_n467));
  OAI21_X1  g281(.A(G131), .B1(new_n452), .B2(new_n460), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n464), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n466), .A2(new_n383), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n383), .B1(new_n466), .B2(new_n469), .ZN(new_n472));
  OAI211_X1 g286(.A(KEYINPUT70), .B(KEYINPUT28), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT28), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n459), .A2(new_n464), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n469), .B1(new_n410), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n367), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n470), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT70), .B1(new_n480), .B2(KEYINPUT28), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n448), .B1(new_n476), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n478), .A2(KEYINPUT30), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT30), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n466), .A2(new_n484), .A3(new_n469), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n471), .B1(new_n486), .B2(new_n367), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT31), .B1(new_n487), .B2(new_n447), .ZN(new_n488));
  INV_X1    g302(.A(new_n485), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n484), .B1(new_n466), .B2(new_n469), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n367), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AND4_X1   g305(.A1(KEYINPUT31), .A2(new_n491), .A3(new_n447), .A4(new_n470), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n482), .B1(new_n488), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G472), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n494), .A3(new_n248), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT32), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n491), .A2(new_n447), .A3(new_n470), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT31), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n487), .A2(KEYINPUT31), .A3(new_n447), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(G902), .B1(new_n501), .B2(new_n482), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT32), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n503), .A3(new_n494), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n479), .A2(KEYINPUT71), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT71), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n472), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n471), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n475), .B1(new_n509), .B2(new_n474), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT29), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n448), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  OR2_X1    g327(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n476), .A2(new_n481), .A3(new_n448), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n487), .A2(new_n447), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n511), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n514), .B(new_n248), .C1(new_n515), .C2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G472), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n505), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT76), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT74), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n329), .B2(G128), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n323), .A2(new_n325), .A3(G128), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT23), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n323), .A2(new_n325), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(KEYINPUT74), .A3(new_n259), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n523), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G110), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n322), .A2(G128), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT23), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n528), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT73), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n524), .B1(new_n533), .B2(new_n530), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n329), .A2(KEYINPUT73), .A3(G128), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g350(.A(KEYINPUT24), .B(G110), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n532), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT75), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n203), .A2(new_n206), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n231), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n539), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  AND2_X1   g358(.A1(new_n534), .A2(new_n535), .ZN(new_n545));
  INV_X1    g359(.A(new_n537), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n545), .A2(new_n546), .B1(new_n230), .B2(new_n231), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n528), .A2(new_n531), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G110), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n542), .B1(new_n532), .B2(new_n538), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(new_n540), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n521), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT77), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT22), .B(G137), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n552), .A2(new_n540), .B1(new_n547), .B2(new_n549), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n539), .A2(new_n543), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT75), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n560), .A2(new_n562), .A3(KEYINPUT76), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n554), .A2(new_n559), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n560), .A2(new_n562), .A3(new_n558), .ZN(new_n565));
  OAI21_X1  g379(.A(G217), .B1(new_n314), .B2(G902), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n564), .A2(new_n248), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT78), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n566), .B(KEYINPUT72), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n564), .A2(new_n248), .A3(new_n565), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n570), .B1(new_n571), .B2(KEYINPUT25), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT25), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n564), .A2(new_n573), .A3(new_n248), .A4(new_n565), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n292), .ZN(new_n578));
  OAI21_X1  g392(.A(G221), .B1(new_n578), .B2(G902), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n372), .A2(new_n406), .A3(new_n449), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT10), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n582), .B1(new_n361), .B2(new_n467), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n415), .A2(new_n357), .A3(KEYINPUT10), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n581), .B(new_n477), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(G110), .B(G140), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n190), .A2(G227), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n415), .A2(new_n357), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n589), .B1(new_n382), .B2(new_n415), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT12), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n590), .A2(new_n591), .A3(new_n477), .ZN(new_n592));
  INV_X1    g406(.A(new_n589), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n359), .A2(new_n415), .A3(new_n360), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT12), .B1(new_n595), .B2(new_n465), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n585), .B(new_n588), .C1(new_n592), .C2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT81), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n591), .B1(new_n590), .B2(new_n477), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n595), .A2(KEYINPUT12), .A3(new_n465), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT81), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n601), .A2(new_n602), .A3(new_n585), .A4(new_n588), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n465), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n588), .B1(new_n606), .B2(new_n585), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(G469), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n610), .A3(new_n248), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n606), .A2(new_n585), .ZN(new_n612));
  INV_X1    g426(.A(new_n588), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n588), .B(KEYINPUT79), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(new_n601), .B2(new_n585), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n248), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(G469), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n580), .B1(new_n611), .B2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n442), .A2(new_n520), .A3(new_n577), .A4(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G101), .ZN(G3));
  INV_X1    g435(.A(new_n318), .ZN(new_n622));
  AOI21_X1  g436(.A(G478), .B1(new_n301), .B2(new_n248), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT33), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n624), .A2(KEYINPUT33), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n299), .B1(new_n298), .B2(new_n278), .ZN(new_n628));
  AOI211_X1 g442(.A(new_n293), .B(new_n277), .C1(new_n297), .C2(new_n288), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n625), .B(new_n627), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT33), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n294), .A2(new_n300), .A3(KEYINPUT97), .A4(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n256), .A2(G902), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n623), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n254), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT96), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n441), .A2(new_n638), .ZN(new_n639));
  OAI211_X1 g453(.A(KEYINPUT96), .B(new_n320), .C1(new_n439), .C2(new_n440), .ZN(new_n640));
  AOI211_X1 g454(.A(new_n622), .B(new_n637), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n493), .A2(new_n248), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(G472), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n495), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n576), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n641), .A2(new_n619), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  NAND2_X1  g462(.A1(new_n247), .A2(KEYINPUT98), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT98), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n239), .A2(new_n245), .A3(new_n650), .A4(new_n246), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n649), .A2(new_n305), .A3(new_n253), .A4(new_n651), .ZN(new_n652));
  AOI211_X1 g466(.A(new_n622), .B(new_n652), .C1(new_n639), .C2(new_n640), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n619), .A3(new_n645), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT99), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT35), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G107), .ZN(G9));
  NOR2_X1   g471(.A1(new_n559), .A2(KEYINPUT36), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT100), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n554), .A2(new_n659), .A3(new_n563), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n659), .B1(new_n554), .B2(new_n563), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n658), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n551), .A2(new_n521), .A3(new_n553), .ZN(new_n664));
  AOI21_X1  g478(.A(KEYINPUT76), .B1(new_n560), .B2(new_n562), .ZN(new_n665));
  OAI21_X1  g479(.A(KEYINPUT100), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n658), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n666), .A2(new_n667), .A3(new_n660), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(G902), .B1(new_n314), .B2(G217), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n669), .A2(new_n670), .B1(new_n572), .B2(new_n574), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n644), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n442), .A2(new_n672), .A3(new_n619), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  NAND2_X1  g489(.A1(new_n639), .A2(new_n640), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n310), .A2(G900), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n315), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n671), .A2(new_n652), .A3(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n676), .A2(new_n680), .A3(new_n520), .A4(new_n619), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G128), .ZN(G30));
  NOR2_X1   g496(.A1(new_n439), .A2(new_n440), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT101), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n683), .B(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n320), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n254), .A2(new_n305), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n607), .B1(new_n598), .B2(new_n603), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n690), .A2(G469), .A3(G902), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n601), .A2(new_n585), .ZN(new_n692));
  OAI22_X1  g506(.A1(new_n692), .A2(new_n615), .B1(new_n612), .B2(new_n613), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n610), .B1(new_n693), .B2(new_n248), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n579), .B1(new_n691), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n678), .B(KEYINPUT39), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n699), .A2(KEYINPUT40), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(KEYINPUT40), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n666), .A2(new_n667), .A3(new_n660), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n667), .B1(new_n666), .B2(new_n660), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n670), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n575), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n497), .B1(new_n509), .B2(new_n447), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n248), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(G472), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n705), .B1(new_n505), .B2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n689), .A2(new_n700), .A3(new_n701), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G143), .ZN(G45));
  AOI211_X1 g525(.A(new_n635), .B(new_n679), .C1(new_n247), .C2(new_n253), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n705), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n676), .A2(new_n520), .A3(new_n619), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G146), .ZN(G48));
  INV_X1    g529(.A(KEYINPUT103), .ZN(new_n716));
  OAI21_X1  g530(.A(G469), .B1(new_n690), .B2(G902), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n611), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  OAI211_X1 g532(.A(KEYINPUT103), .B(G469), .C1(new_n690), .C2(G902), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT104), .B1(new_n720), .B2(new_n579), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT104), .ZN(new_n722));
  AOI211_X1 g536(.A(new_n722), .B(new_n580), .C1(new_n718), .C2(new_n719), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  AOI22_X1  g538(.A1(new_n496), .A2(new_n504), .B1(new_n518), .B2(G472), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n576), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n641), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT41), .B(G113), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G15));
  NAND3_X1  g543(.A1(new_n653), .A2(new_n724), .A3(new_n726), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT105), .B(G116), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G18));
  AOI21_X1  g546(.A(new_n725), .B1(new_n639), .B2(new_n640), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n580), .B1(new_n718), .B2(new_n719), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n319), .A2(new_n671), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G119), .ZN(G21));
  AOI211_X1 g551(.A(new_n622), .B(new_n688), .C1(new_n639), .C2(new_n640), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT106), .B(G472), .ZN(new_n739));
  AOI22_X1  g553(.A1(new_n448), .A2(new_n510), .B1(new_n499), .B2(new_n500), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n494), .A2(new_n248), .ZN(new_n741));
  OAI22_X1  g555(.A1(new_n502), .A2(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n576), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n569), .A2(KEYINPUT107), .A3(new_n575), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n742), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n738), .A2(new_n724), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  NAND2_X1  g562(.A1(new_n510), .A2(new_n448), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n741), .B1(new_n749), .B2(new_n501), .ZN(new_n750));
  INV_X1    g564(.A(new_n739), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n750), .B1(new_n642), .B2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n676), .A2(new_n713), .A3(new_n734), .A4(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G125), .ZN(G27));
  INV_X1    g568(.A(KEYINPUT108), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n505), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n496), .A2(new_n504), .A3(KEYINPUT108), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n519), .A3(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n683), .A2(new_n619), .A3(new_n712), .A4(new_n320), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT42), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n744), .A2(new_n745), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n758), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n374), .ZN(new_n764));
  AOI22_X1  g578(.A1(new_n361), .A2(new_n347), .B1(new_n367), .B2(new_n372), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n391), .B1(new_n765), .B2(new_n321), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n388), .A2(KEYINPUT83), .A3(new_n389), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n764), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n375), .B1(new_n768), .B2(KEYINPUT6), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n438), .B1(new_n769), .B2(new_n419), .ZN(new_n770));
  INV_X1    g584(.A(new_n422), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n421), .A2(new_n422), .A3(new_n438), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n320), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n695), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n520), .A2(new_n775), .A3(new_n577), .A4(new_n712), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n760), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n763), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G131), .ZN(G33));
  NOR2_X1   g593(.A1(new_n652), .A2(new_n679), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n520), .A2(new_n780), .A3(new_n775), .A4(new_n577), .ZN(new_n781));
  XOR2_X1   g595(.A(KEYINPUT109), .B(G134), .Z(new_n782));
  XNOR2_X1  g596(.A(new_n781), .B(new_n782), .ZN(G36));
  NAND2_X1  g597(.A1(new_n255), .A2(new_n636), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT43), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n644), .A3(new_n705), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT44), .ZN(new_n789));
  OR3_X1    g603(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n774), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n788), .B1(new_n787), .B2(new_n789), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT113), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n693), .B(KEYINPUT45), .ZN(new_n795));
  OAI21_X1  g609(.A(G469), .B1(new_n795), .B2(G902), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(KEYINPUT46), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(KEYINPUT46), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(KEYINPUT110), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT110), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n796), .A2(new_n800), .A3(KEYINPUT46), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n799), .A2(new_n611), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n797), .B1(new_n802), .B2(KEYINPUT111), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(KEYINPUT111), .B2(new_n802), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n804), .A2(new_n579), .A3(new_n696), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n787), .A2(new_n789), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n790), .A2(new_n807), .A3(new_n791), .A4(new_n792), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n794), .A2(new_n805), .A3(new_n806), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G137), .ZN(G39));
  NAND4_X1  g624(.A1(new_n725), .A2(new_n576), .A3(new_n712), .A4(new_n791), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n804), .A2(KEYINPUT47), .A3(new_n579), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT47), .B1(new_n804), .B2(new_n579), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G140), .ZN(G42));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n817));
  INV_X1    g631(.A(new_n688), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n678), .B(KEYINPUT116), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n695), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n709), .A2(new_n676), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(new_n681), .A3(new_n714), .A4(new_n753), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n733), .B(new_n619), .C1(new_n680), .C2(new_n713), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n825), .A2(KEYINPUT52), .A3(new_n753), .A4(new_n821), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n705), .A2(new_n752), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT114), .B1(new_n759), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n671), .A2(new_n742), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n830), .A2(new_n775), .A3(new_n831), .A4(new_n712), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n649), .A2(new_n253), .A3(new_n651), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n835), .A2(new_n305), .A3(new_n679), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n520), .A2(new_n705), .A3(new_n836), .A4(new_n775), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n833), .A2(new_n834), .A3(new_n781), .A4(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n637), .B1(new_n306), .B2(new_n254), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n441), .A2(new_n622), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n645), .A2(new_n619), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n620), .A2(new_n841), .A3(new_n673), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n838), .A2(new_n778), .A3(new_n842), .ZN(new_n843));
  AND4_X1   g657(.A1(new_n727), .A2(new_n730), .A3(new_n747), .A4(new_n736), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n833), .A2(new_n781), .A3(new_n837), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT115), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n827), .A2(new_n843), .A3(new_n844), .A4(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n848));
  OR2_X1    g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n847), .A2(KEYINPUT119), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT119), .B1(new_n847), .B2(new_n850), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n817), .B(new_n849), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n847), .A2(KEYINPUT118), .A3(new_n850), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n847), .A2(new_n848), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n847), .A2(new_n850), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n853), .B1(new_n859), .B2(new_n817), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n758), .A2(new_n762), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n786), .A2(new_n316), .ZN(new_n863));
  INV_X1    g677(.A(new_n734), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n774), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT48), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n863), .A2(new_n746), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n676), .A2(new_n734), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n313), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n505), .A2(new_n708), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n871), .A2(new_n576), .A3(new_n315), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n865), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n873), .A2(new_n637), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n867), .A2(new_n875), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n876), .B(KEYINPUT121), .Z(new_n877));
  NAND3_X1  g691(.A1(new_n863), .A2(new_n830), .A3(new_n865), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n255), .A2(new_n635), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n878), .B1(new_n873), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT120), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n881), .A2(KEYINPUT50), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n686), .A2(new_n687), .A3(new_n734), .ZN(new_n883));
  OR3_X1    g697(.A1(new_n868), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n882), .B1(new_n868), .B2(new_n883), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n880), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n579), .B1(new_n718), .B2(new_n719), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n813), .A2(new_n814), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n863), .A2(new_n746), .A3(new_n791), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT51), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g706(.A(KEYINPUT51), .B(new_n886), .C1(new_n888), .C2(new_n889), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n877), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  OAI22_X1  g708(.A1(new_n860), .A2(new_n894), .B1(G952), .B2(G953), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n720), .B(KEYINPUT49), .Z(new_n896));
  NOR4_X1   g710(.A1(new_n871), .A2(new_n580), .A3(new_n687), .A4(new_n784), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(new_n686), .A3(new_n762), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n895), .B1(new_n896), .B2(new_n898), .ZN(G75));
  OAI21_X1  g713(.A(new_n849), .B1(new_n851), .B2(new_n852), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n900), .A2(G210), .A3(G902), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT56), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n395), .B(new_n419), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT55), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n904), .B1(new_n901), .B2(new_n902), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n190), .A2(G952), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT122), .Z(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n905), .A2(new_n906), .A3(new_n909), .ZN(G51));
  NAND2_X1  g724(.A1(G469), .A2(G902), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT123), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT57), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n847), .A2(new_n850), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n847), .A2(KEYINPUT119), .A3(new_n850), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n817), .B1(new_n918), .B2(new_n849), .ZN(new_n919));
  INV_X1    g733(.A(new_n853), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n913), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n609), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n248), .B1(new_n918), .B2(new_n849), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n923), .A2(G469), .A3(new_n795), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n907), .B1(new_n922), .B2(new_n924), .ZN(G54));
  NAND2_X1  g739(.A1(KEYINPUT58), .A2(G475), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT124), .Z(new_n927));
  AND3_X1   g741(.A1(new_n923), .A2(new_n242), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n242), .B1(new_n923), .B2(new_n927), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n928), .A2(new_n929), .A3(new_n907), .ZN(G60));
  NOR2_X1   g744(.A1(new_n919), .A2(new_n920), .ZN(new_n931));
  NAND2_X1  g745(.A1(G478), .A2(G902), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT59), .Z(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n633), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n908), .B1(new_n931), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n633), .B1(new_n860), .B2(new_n934), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(G63));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT60), .Z(new_n940));
  NAND3_X1  g754(.A1(new_n900), .A2(new_n669), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n940), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n918), .B2(new_n849), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n564), .A2(new_n565), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n941), .B(new_n908), .C1(new_n943), .C2(new_n945), .ZN(new_n946));
  OAI211_X1 g760(.A(KEYINPUT125), .B(new_n908), .C1(new_n943), .C2(new_n945), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n900), .A2(new_n940), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n909), .B1(new_n950), .B2(new_n944), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n951), .B(new_n941), .C1(KEYINPUT125), .C2(KEYINPUT61), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n949), .A2(new_n952), .ZN(G66));
  AOI21_X1  g767(.A(new_n190), .B1(new_n308), .B2(G224), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n844), .A2(new_n842), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n954), .B1(new_n955), .B2(new_n190), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n769), .B1(G898), .B2(new_n190), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n956), .B(new_n957), .Z(G69));
  NOR2_X1   g772(.A1(new_n210), .A2(new_n211), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n486), .B(new_n959), .Z(new_n960));
  NAND2_X1  g774(.A1(G900), .A2(G953), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n805), .A2(new_n676), .A3(new_n818), .A4(new_n862), .ZN(new_n962));
  AND4_X1   g776(.A1(new_n753), .A2(new_n778), .A3(new_n781), .A4(new_n825), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n809), .A2(new_n815), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n960), .B(new_n961), .C1(new_n964), .C2(G953), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n710), .A2(new_n753), .A3(new_n825), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT62), .Z(new_n967));
  NAND4_X1  g781(.A1(new_n726), .A2(new_n698), .A3(new_n791), .A4(new_n839), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n967), .A2(new_n809), .A3(new_n815), .A4(new_n968), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n969), .A2(new_n190), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n965), .B1(new_n970), .B2(new_n960), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(G72));
  NAND2_X1  g787(.A1(G472), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT63), .Z(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(new_n969), .B2(new_n955), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n487), .B(KEYINPUT126), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n976), .A2(new_n447), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n975), .B1(new_n964), .B2(new_n955), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n977), .A2(new_n447), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT127), .Z(new_n981));
  AND2_X1   g795(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n516), .A2(new_n497), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n975), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n859), .A2(new_n984), .ZN(new_n985));
  NOR4_X1   g799(.A1(new_n978), .A2(new_n982), .A3(new_n907), .A4(new_n985), .ZN(G57));
endmodule


