

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574;

  XNOR2_X1 U317 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U318 ( .A(n460), .B(n459), .ZN(n506) );
  XNOR2_X1 U319 ( .A(n458), .B(KEYINPUT103), .ZN(n459) );
  XNOR2_X1 U320 ( .A(n382), .B(n381), .ZN(n544) );
  OR2_X1 U321 ( .A1(n538), .A2(n561), .ZN(n368) );
  XNOR2_X1 U322 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n386) );
  XNOR2_X1 U323 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U324 ( .A(G134GAT), .B(KEYINPUT78), .Z(n410) );
  XNOR2_X1 U325 ( .A(n405), .B(n404), .ZN(n409) );
  INV_X1 U326 ( .A(n412), .ZN(n335) );
  XNOR2_X1 U327 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U328 ( .A(n336), .B(n335), .ZN(n343) );
  XNOR2_X1 U329 ( .A(n392), .B(KEYINPUT48), .ZN(n393) );
  XNOR2_X1 U330 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U331 ( .A(n343), .B(n342), .ZN(n345) );
  OR2_X1 U332 ( .A1(n438), .A2(n491), .ZN(n439) );
  XOR2_X1 U333 ( .A(n564), .B(KEYINPUT41), .Z(n538) );
  XNOR2_X1 U334 ( .A(n439), .B(KEYINPUT119), .ZN(n553) );
  INV_X1 U335 ( .A(n443), .ZN(n508) );
  XNOR2_X1 U336 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n440) );
  XNOR2_X1 U337 ( .A(n463), .B(KEYINPUT106), .ZN(n464) );
  XNOR2_X1 U338 ( .A(n441), .B(n440), .ZN(G1351GAT) );
  XNOR2_X1 U339 ( .A(n465), .B(n464), .ZN(G1331GAT) );
  XOR2_X1 U340 ( .A(G218GAT), .B(G162GAT), .Z(n378) );
  XOR2_X1 U341 ( .A(G22GAT), .B(G155GAT), .Z(n322) );
  XNOR2_X1 U342 ( .A(n378), .B(n322), .ZN(n287) );
  XOR2_X1 U343 ( .A(KEYINPUT2), .B(KEYINPUT88), .Z(n286) );
  XNOR2_X1 U344 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n285) );
  XNOR2_X1 U345 ( .A(n286), .B(n285), .ZN(n411) );
  XNOR2_X1 U346 ( .A(n287), .B(n411), .ZN(n292) );
  XNOR2_X1 U347 ( .A(G197GAT), .B(KEYINPUT87), .ZN(n288) );
  XNOR2_X1 U348 ( .A(n288), .B(KEYINPUT21), .ZN(n311) );
  XOR2_X1 U349 ( .A(G78GAT), .B(n311), .Z(n290) );
  NAND2_X1 U350 ( .A1(G228GAT), .A2(G233GAT), .ZN(n289) );
  XNOR2_X1 U351 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U352 ( .A(n292), .B(n291), .Z(n300) );
  XOR2_X1 U353 ( .A(KEYINPUT22), .B(G211GAT), .Z(n294) );
  XNOR2_X1 U354 ( .A(G50GAT), .B(G106GAT), .ZN(n293) );
  XNOR2_X1 U355 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U356 ( .A(G148GAT), .B(G204GAT), .Z(n296) );
  XNOR2_X1 U357 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n295) );
  XNOR2_X1 U358 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U359 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U360 ( .A(n300), .B(n299), .ZN(n449) );
  XOR2_X1 U361 ( .A(KEYINPUT19), .B(G190GAT), .Z(n302) );
  XNOR2_X1 U362 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n301) );
  XNOR2_X1 U363 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U364 ( .A(G169GAT), .B(n303), .Z(n433) );
  XOR2_X1 U365 ( .A(G64GAT), .B(KEYINPUT76), .Z(n305) );
  XNOR2_X1 U366 ( .A(G176GAT), .B(G204GAT), .ZN(n304) );
  XNOR2_X1 U367 ( .A(n305), .B(n304), .ZN(n341) );
  XNOR2_X1 U368 ( .A(n433), .B(n341), .ZN(n315) );
  XOR2_X1 U369 ( .A(G92GAT), .B(G218GAT), .Z(n307) );
  NAND2_X1 U370 ( .A1(G226GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U371 ( .A(n307), .B(n306), .ZN(n310) );
  XOR2_X1 U372 ( .A(KEYINPUT80), .B(G211GAT), .Z(n309) );
  XNOR2_X1 U373 ( .A(G8GAT), .B(G183GAT), .ZN(n308) );
  XNOR2_X1 U374 ( .A(n309), .B(n308), .ZN(n326) );
  XOR2_X1 U375 ( .A(n310), .B(n326), .Z(n313) );
  XNOR2_X1 U376 ( .A(G36GAT), .B(n311), .ZN(n312) );
  XNOR2_X1 U377 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U378 ( .A(n315), .B(n314), .ZN(n489) );
  XNOR2_X1 U379 ( .A(G15GAT), .B(G1GAT), .ZN(n316) );
  XNOR2_X1 U380 ( .A(n316), .B(KEYINPUT71), .ZN(n356) );
  XOR2_X1 U381 ( .A(KEYINPUT13), .B(G57GAT), .Z(n318) );
  XNOR2_X1 U382 ( .A(G71GAT), .B(G78GAT), .ZN(n317) );
  XNOR2_X1 U383 ( .A(n318), .B(n317), .ZN(n333) );
  XNOR2_X1 U384 ( .A(n356), .B(n333), .ZN(n330) );
  XOR2_X1 U385 ( .A(KEYINPUT81), .B(KEYINPUT14), .Z(n320) );
  XNOR2_X1 U386 ( .A(G127GAT), .B(G64GAT), .ZN(n319) );
  XNOR2_X1 U387 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U388 ( .A(n322), .B(n321), .Z(n324) );
  NAND2_X1 U389 ( .A1(G231GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U390 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U391 ( .A(n325), .B(KEYINPUT15), .Z(n328) );
  XNOR2_X1 U392 ( .A(n326), .B(KEYINPUT12), .ZN(n327) );
  XNOR2_X1 U393 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U394 ( .A(n330), .B(n329), .ZN(n567) );
  XNOR2_X1 U395 ( .A(n567), .B(KEYINPUT111), .ZN(n524) );
  XOR2_X1 U396 ( .A(KEYINPUT33), .B(KEYINPUT74), .Z(n332) );
  XNOR2_X1 U397 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n331) );
  XNOR2_X1 U398 ( .A(n332), .B(n331), .ZN(n334) );
  XOR2_X1 U399 ( .A(n334), .B(n333), .Z(n336) );
  XOR2_X1 U400 ( .A(G120GAT), .B(G148GAT), .Z(n412) );
  INV_X1 U401 ( .A(G106GAT), .ZN(n340) );
  XOR2_X1 U402 ( .A(KEYINPUT75), .B(G92GAT), .Z(n338) );
  XNOR2_X1 U403 ( .A(G99GAT), .B(G85GAT), .ZN(n337) );
  XNOR2_X1 U404 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U405 ( .A(n340), .B(n339), .ZN(n377) );
  XNOR2_X1 U406 ( .A(n341), .B(n377), .ZN(n342) );
  NAND2_X1 U407 ( .A1(G230GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n564) );
  XOR2_X1 U409 ( .A(G43GAT), .B(G29GAT), .Z(n347) );
  XNOR2_X1 U410 ( .A(KEYINPUT70), .B(G50GAT), .ZN(n346) );
  XNOR2_X1 U411 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U412 ( .A(n348), .B(KEYINPUT8), .Z(n350) );
  XNOR2_X1 U413 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n349) );
  XNOR2_X1 U414 ( .A(n350), .B(n349), .ZN(n382) );
  XOR2_X1 U415 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n352) );
  XNOR2_X1 U416 ( .A(KEYINPUT29), .B(KEYINPUT67), .ZN(n351) );
  XNOR2_X1 U417 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U418 ( .A(n382), .B(n353), .ZN(n366) );
  XOR2_X1 U419 ( .A(G197GAT), .B(G22GAT), .Z(n355) );
  XNOR2_X1 U420 ( .A(G169GAT), .B(G113GAT), .ZN(n354) );
  XNOR2_X1 U421 ( .A(n355), .B(n354), .ZN(n364) );
  XOR2_X1 U422 ( .A(n356), .B(KEYINPUT72), .Z(n358) );
  NAND2_X1 U423 ( .A1(G229GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U424 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U425 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n360) );
  XNOR2_X1 U426 ( .A(G141GAT), .B(G8GAT), .ZN(n359) );
  XNOR2_X1 U427 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U428 ( .A(n362), .B(n361), .Z(n363) );
  XNOR2_X1 U429 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n561) );
  INV_X1 U431 ( .A(KEYINPUT46), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n368), .B(n367), .ZN(n369) );
  NOR2_X1 U433 ( .A1(n524), .A2(n369), .ZN(n370) );
  XNOR2_X1 U434 ( .A(n370), .B(KEYINPUT112), .ZN(n383) );
  XOR2_X1 U435 ( .A(KEYINPUT77), .B(n410), .Z(n372) );
  NAND2_X1 U436 ( .A1(G232GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U437 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U438 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n374) );
  XNOR2_X1 U439 ( .A(G190GAT), .B(KEYINPUT9), .ZN(n373) );
  XNOR2_X1 U440 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U441 ( .A(n376), .B(n375), .Z(n380) );
  XNOR2_X1 U442 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U443 ( .A(n380), .B(n379), .ZN(n381) );
  NAND2_X1 U444 ( .A1(n383), .A2(n544), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n384), .B(KEYINPUT47), .ZN(n391) );
  XNOR2_X1 U446 ( .A(KEYINPUT79), .B(n544), .ZN(n528) );
  XNOR2_X1 U447 ( .A(KEYINPUT36), .B(KEYINPUT101), .ZN(n385) );
  XNOR2_X1 U448 ( .A(n528), .B(n385), .ZN(n571) );
  NOR2_X1 U449 ( .A1(n567), .A2(n571), .ZN(n387) );
  NAND2_X1 U450 ( .A1(n388), .A2(n564), .ZN(n389) );
  XNOR2_X1 U451 ( .A(KEYINPUT73), .B(n561), .ZN(n547) );
  NOR2_X1 U452 ( .A1(n389), .A2(n547), .ZN(n390) );
  NOR2_X1 U453 ( .A1(n391), .A2(n390), .ZN(n394) );
  INV_X1 U454 ( .A(KEYINPUT113), .ZN(n392) );
  XNOR2_X1 U455 ( .A(n394), .B(n393), .ZN(n533) );
  NOR2_X1 U456 ( .A1(n489), .A2(n533), .ZN(n395) );
  XNOR2_X1 U457 ( .A(n395), .B(KEYINPUT54), .ZN(n418) );
  XOR2_X1 U458 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n397) );
  XNOR2_X1 U459 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n396) );
  XNOR2_X1 U460 ( .A(n397), .B(n396), .ZN(n417) );
  XOR2_X1 U461 ( .A(G127GAT), .B(KEYINPUT0), .Z(n399) );
  XNOR2_X1 U462 ( .A(G113GAT), .B(KEYINPUT82), .ZN(n398) );
  XNOR2_X1 U463 ( .A(n399), .B(n398), .ZN(n429) );
  XOR2_X1 U464 ( .A(n429), .B(G57GAT), .Z(n405) );
  XOR2_X1 U465 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n401) );
  XNOR2_X1 U466 ( .A(KEYINPUT1), .B(KEYINPUT91), .ZN(n400) );
  XNOR2_X1 U467 ( .A(n401), .B(n400), .ZN(n403) );
  NAND2_X1 U468 ( .A1(G225GAT), .A2(G233GAT), .ZN(n402) );
  XOR2_X1 U469 ( .A(G85GAT), .B(G155GAT), .Z(n407) );
  XNOR2_X1 U470 ( .A(G29GAT), .B(G162GAT), .ZN(n406) );
  XNOR2_X1 U471 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U472 ( .A(n409), .B(n408), .ZN(n415) );
  XOR2_X1 U473 ( .A(n411), .B(n410), .Z(n413) );
  XNOR2_X1 U474 ( .A(n417), .B(n416), .ZN(n443) );
  NAND2_X1 U475 ( .A1(n418), .A2(n443), .ZN(n558) );
  NOR2_X1 U476 ( .A1(n449), .A2(n558), .ZN(n420) );
  XNOR2_X1 U477 ( .A(KEYINPUT118), .B(KEYINPUT55), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n420), .B(n419), .ZN(n438) );
  XOR2_X1 U479 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n422) );
  XNOR2_X1 U480 ( .A(KEYINPUT86), .B(KEYINPUT85), .ZN(n421) );
  XNOR2_X1 U481 ( .A(n422), .B(n421), .ZN(n437) );
  XOR2_X1 U482 ( .A(G120GAT), .B(G134GAT), .Z(n424) );
  XNOR2_X1 U483 ( .A(G43GAT), .B(G99GAT), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U485 ( .A(KEYINPUT20), .B(G183GAT), .Z(n426) );
  XNOR2_X1 U486 ( .A(G15GAT), .B(G71GAT), .ZN(n425) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U488 ( .A(n428), .B(n427), .Z(n435) );
  XOR2_X1 U489 ( .A(n429), .B(G176GAT), .Z(n431) );
  NAND2_X1 U490 ( .A1(G227GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U491 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U492 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U494 ( .A(n437), .B(n436), .ZN(n491) );
  NAND2_X1 U495 ( .A1(n553), .A2(n528), .ZN(n441) );
  XOR2_X1 U496 ( .A(n449), .B(KEYINPUT65), .Z(n442) );
  XNOR2_X1 U497 ( .A(KEYINPUT28), .B(n442), .ZN(n515) );
  INV_X1 U498 ( .A(n515), .ZN(n462) );
  INV_X1 U499 ( .A(n491), .ZN(n519) );
  XNOR2_X1 U500 ( .A(n489), .B(KEYINPUT27), .ZN(n447) );
  NAND2_X1 U501 ( .A1(n508), .A2(n462), .ZN(n444) );
  NOR2_X1 U502 ( .A1(n447), .A2(n444), .ZN(n518) );
  XOR2_X1 U503 ( .A(KEYINPUT92), .B(n518), .Z(n445) );
  NOR2_X1 U504 ( .A1(n519), .A2(n445), .ZN(n454) );
  NAND2_X1 U505 ( .A1(n491), .A2(n449), .ZN(n446) );
  XNOR2_X1 U506 ( .A(n446), .B(KEYINPUT26), .ZN(n559) );
  NOR2_X1 U507 ( .A1(n559), .A2(n447), .ZN(n535) );
  NOR2_X1 U508 ( .A1(n489), .A2(n491), .ZN(n448) );
  NOR2_X1 U509 ( .A1(n449), .A2(n448), .ZN(n450) );
  XOR2_X1 U510 ( .A(KEYINPUT25), .B(n450), .Z(n451) );
  NOR2_X1 U511 ( .A1(n535), .A2(n451), .ZN(n452) );
  NOR2_X1 U512 ( .A1(n508), .A2(n452), .ZN(n453) );
  NOR2_X1 U513 ( .A1(n454), .A2(n453), .ZN(n455) );
  XNOR2_X1 U514 ( .A(KEYINPUT93), .B(n455), .ZN(n469) );
  NAND2_X1 U515 ( .A1(n469), .A2(n567), .ZN(n456) );
  XNOR2_X1 U516 ( .A(n456), .B(KEYINPUT102), .ZN(n457) );
  NOR2_X1 U517 ( .A1(n571), .A2(n457), .ZN(n460) );
  INV_X1 U518 ( .A(KEYINPUT37), .ZN(n458) );
  NAND2_X1 U519 ( .A1(n547), .A2(n564), .ZN(n472) );
  NOR2_X1 U520 ( .A1(n506), .A2(n472), .ZN(n461) );
  XOR2_X1 U521 ( .A(KEYINPUT38), .B(n461), .Z(n492) );
  NOR2_X1 U522 ( .A1(n462), .A2(n492), .ZN(n465) );
  INV_X1 U523 ( .A(G50GAT), .ZN(n463) );
  NAND2_X1 U524 ( .A1(n524), .A2(n553), .ZN(n467) );
  XNOR2_X1 U525 ( .A(G183GAT), .B(KEYINPUT122), .ZN(n466) );
  XNOR2_X1 U526 ( .A(n467), .B(n466), .ZN(G1350GAT) );
  XNOR2_X1 U527 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n477) );
  XOR2_X1 U528 ( .A(G1GAT), .B(KEYINPUT34), .Z(n475) );
  NOR2_X1 U529 ( .A1(n528), .A2(n567), .ZN(n468) );
  XNOR2_X1 U530 ( .A(KEYINPUT16), .B(n468), .ZN(n470) );
  NAND2_X1 U531 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n471), .B(KEYINPUT94), .ZN(n497) );
  NOR2_X1 U533 ( .A1(n497), .A2(n472), .ZN(n473) );
  XOR2_X1 U534 ( .A(KEYINPUT95), .B(n473), .Z(n482) );
  NAND2_X1 U535 ( .A1(n482), .A2(n508), .ZN(n474) );
  XNOR2_X1 U536 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U537 ( .A(n477), .B(n476), .ZN(G1324GAT) );
  INV_X1 U538 ( .A(n489), .ZN(n510) );
  NAND2_X1 U539 ( .A1(n510), .A2(n482), .ZN(n478) );
  XNOR2_X1 U540 ( .A(n478), .B(KEYINPUT98), .ZN(n479) );
  XNOR2_X1 U541 ( .A(G8GAT), .B(n479), .ZN(G1325GAT) );
  XOR2_X1 U542 ( .A(G15GAT), .B(KEYINPUT35), .Z(n481) );
  NAND2_X1 U543 ( .A1(n482), .A2(n519), .ZN(n480) );
  XNOR2_X1 U544 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n484) );
  NAND2_X1 U546 ( .A1(n482), .A2(n515), .ZN(n483) );
  XNOR2_X1 U547 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U548 ( .A(G22GAT), .B(n485), .ZN(G1327GAT) );
  NOR2_X1 U549 ( .A1(n492), .A2(n443), .ZN(n487) );
  XNOR2_X1 U550 ( .A(KEYINPUT104), .B(KEYINPUT39), .ZN(n486) );
  XNOR2_X1 U551 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(n488), .ZN(G1328GAT) );
  NOR2_X1 U553 ( .A1(n489), .A2(n492), .ZN(n490) );
  XOR2_X1 U554 ( .A(G36GAT), .B(n490), .Z(G1329GAT) );
  NOR2_X1 U555 ( .A1(n492), .A2(n491), .ZN(n494) );
  XNOR2_X1 U556 ( .A(KEYINPUT40), .B(KEYINPUT105), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U558 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  XNOR2_X1 U559 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n500) );
  XNOR2_X1 U560 ( .A(n538), .B(KEYINPUT107), .ZN(n552) );
  NAND2_X1 U561 ( .A1(n552), .A2(n561), .ZN(n496) );
  XNOR2_X1 U562 ( .A(n496), .B(KEYINPUT108), .ZN(n507) );
  NOR2_X1 U563 ( .A1(n507), .A2(n497), .ZN(n498) );
  XOR2_X1 U564 ( .A(KEYINPUT109), .B(n498), .Z(n503) );
  NAND2_X1 U565 ( .A1(n508), .A2(n503), .ZN(n499) );
  XNOR2_X1 U566 ( .A(n500), .B(n499), .ZN(G1332GAT) );
  NAND2_X1 U567 ( .A1(n510), .A2(n503), .ZN(n501) );
  XNOR2_X1 U568 ( .A(n501), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U569 ( .A1(n503), .A2(n519), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n502), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(G78GAT), .B(KEYINPUT43), .Z(n505) );
  NAND2_X1 U572 ( .A1(n503), .A2(n515), .ZN(n504) );
  XNOR2_X1 U573 ( .A(n505), .B(n504), .ZN(G1335GAT) );
  NOR2_X1 U574 ( .A1(n507), .A2(n506), .ZN(n514) );
  NAND2_X1 U575 ( .A1(n508), .A2(n514), .ZN(n509) );
  XNOR2_X1 U576 ( .A(G85GAT), .B(n509), .ZN(G1336GAT) );
  XNOR2_X1 U577 ( .A(G92GAT), .B(KEYINPUT110), .ZN(n512) );
  NAND2_X1 U578 ( .A1(n514), .A2(n510), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n512), .B(n511), .ZN(G1337GAT) );
  NAND2_X1 U580 ( .A1(n514), .A2(n519), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n513), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U582 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n516), .B(KEYINPUT44), .ZN(n517) );
  XNOR2_X1 U584 ( .A(G106GAT), .B(n517), .ZN(G1339GAT) );
  NAND2_X1 U585 ( .A1(n519), .A2(n518), .ZN(n520) );
  NOR2_X1 U586 ( .A1(n533), .A2(n520), .ZN(n529) );
  NAND2_X1 U587 ( .A1(n547), .A2(n529), .ZN(n521) );
  XNOR2_X1 U588 ( .A(G113GAT), .B(n521), .ZN(G1340GAT) );
  XOR2_X1 U589 ( .A(G120GAT), .B(KEYINPUT49), .Z(n523) );
  NAND2_X1 U590 ( .A1(n529), .A2(n552), .ZN(n522) );
  XNOR2_X1 U591 ( .A(n523), .B(n522), .ZN(G1341GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n526) );
  NAND2_X1 U593 ( .A1(n529), .A2(n524), .ZN(n525) );
  XNOR2_X1 U594 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U595 ( .A(G127GAT), .B(n527), .Z(G1342GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n531) );
  NAND2_X1 U597 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U599 ( .A(G134GAT), .B(n532), .Z(G1343GAT) );
  NOR2_X1 U600 ( .A1(n443), .A2(n533), .ZN(n534) );
  NAND2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U602 ( .A(KEYINPUT116), .B(n536), .ZN(n545) );
  NOR2_X1 U603 ( .A1(n545), .A2(n561), .ZN(n537) );
  XOR2_X1 U604 ( .A(G141GAT), .B(n537), .Z(G1344GAT) );
  XNOR2_X1 U605 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n540) );
  NOR2_X1 U606 ( .A1(n538), .A2(n545), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(n541), .ZN(G1345GAT) );
  XNOR2_X1 U609 ( .A(G155GAT), .B(KEYINPUT117), .ZN(n543) );
  NOR2_X1 U610 ( .A1(n567), .A2(n545), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(G1346GAT) );
  NOR2_X1 U612 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U613 ( .A(G162GAT), .B(n546), .Z(G1347GAT) );
  NAND2_X1 U614 ( .A1(n547), .A2(n553), .ZN(n548) );
  XNOR2_X1 U615 ( .A(G169GAT), .B(n548), .ZN(G1348GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n550) );
  XNOR2_X1 U617 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U619 ( .A(KEYINPUT56), .B(n551), .Z(n555) );
  NAND2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1349GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n557) );
  XNOR2_X1 U623 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n563) );
  NOR2_X1 U625 ( .A1(n558), .A2(n559), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(KEYINPUT123), .ZN(n570) );
  NOR2_X1 U627 ( .A1(n561), .A2(n570), .ZN(n562) );
  XOR2_X1 U628 ( .A(n563), .B(n562), .Z(G1352GAT) );
  NOR2_X1 U629 ( .A1(n564), .A2(n570), .ZN(n566) );
  XNOR2_X1 U630 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(G1353GAT) );
  NOR2_X1 U632 ( .A1(n567), .A2(n570), .ZN(n569) );
  XNOR2_X1 U633 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1354GAT) );
  NOR2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n573) );
  XNOR2_X1 U636 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U638 ( .A(G218GAT), .B(n574), .Z(G1355GAT) );
endmodule

