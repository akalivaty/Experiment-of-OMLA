//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 0 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  XOR2_X1   g000(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT88), .B(G143), .ZN(new_n189));
  NOR2_X1   g003(.A1(G237), .A2(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G214), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT88), .ZN(new_n193));
  AOI22_X1  g007(.A1(new_n190), .A2(G214), .B1(new_n193), .B2(G143), .ZN(new_n194));
  OAI21_X1  g008(.A(G131), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n194), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n196), .B(new_n197), .C1(new_n191), .C2(new_n189), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT17), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n195), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  INV_X1    g015(.A(G140), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G125), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G140), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT73), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(KEYINPUT73), .A3(G140), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(KEYINPUT16), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n203), .A2(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n201), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n209), .A2(new_n201), .A3(new_n211), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n196), .B1(new_n191), .B2(new_n189), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT17), .A3(G131), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n200), .A2(new_n213), .A3(new_n214), .A4(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G113), .B(G122), .ZN(new_n218));
  INV_X1    g032(.A(G104), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n218), .B(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n203), .A2(new_n205), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n201), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n207), .A2(new_n208), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n223), .B1(new_n224), .B2(new_n201), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT18), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(new_n197), .ZN(new_n227));
  OAI221_X1 g041(.A(new_n225), .B1(new_n215), .B2(new_n227), .C1(new_n195), .C2(new_n226), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n217), .A2(new_n220), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n224), .A2(KEYINPUT19), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT19), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n221), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(G146), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT89), .B1(new_n233), .B2(new_n212), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n195), .A2(new_n198), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n231), .B1(new_n207), .B2(new_n208), .ZN(new_n236));
  INV_X1    g050(.A(new_n232), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n201), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT89), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n213), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n234), .A2(new_n235), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n228), .ZN(new_n242));
  INV_X1    g056(.A(new_n220), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n229), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(G475), .A2(G902), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n188), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(KEYINPUT20), .B1(new_n246), .B2(KEYINPUT90), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n220), .B1(new_n241), .B2(new_n228), .ZN(new_n249));
  OAI221_X1 g063(.A(new_n248), .B1(KEYINPUT90), .B2(new_n246), .C1(new_n249), .C2(new_n229), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G902), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n220), .B1(new_n217), .B2(new_n228), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n252), .B1(new_n229), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G475), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G953), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n257), .A2(G952), .ZN(new_n258));
  INV_X1    g072(.A(G234), .ZN(new_n259));
  INV_X1    g073(.A(G237), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AOI211_X1 g076(.A(new_n252), .B(new_n257), .C1(G234), .C2(G237), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT21), .B(G898), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G478), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(KEYINPUT15), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G143), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G128), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(G128), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT13), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G128), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(G143), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT13), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n273), .A2(KEYINPUT91), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT91), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n278), .B(new_n270), .C1(new_n271), .C2(new_n272), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G134), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT92), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n273), .A2(KEYINPUT91), .A3(new_n276), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT92), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n282), .A2(new_n283), .A3(G134), .A4(new_n279), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n275), .A2(new_n271), .A3(G134), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(G116), .B(G122), .ZN(new_n288));
  INV_X1    g102(.A(G107), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n288), .A2(new_n289), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n287), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n285), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n275), .A2(new_n271), .ZN(new_n296));
  INV_X1    g110(.A(G134), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n290), .B1(new_n298), .B2(new_n286), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT93), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT14), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n288), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G116), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G122), .ZN(new_n304));
  OAI21_X1  g118(.A(G107), .B1(new_n304), .B2(new_n301), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n300), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n305), .B1(new_n301), .B2(new_n288), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT93), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n299), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT9), .B(G234), .ZN(new_n311));
  INV_X1    g125(.A(G217), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n311), .A2(new_n312), .A3(G953), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n295), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n313), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n293), .B1(new_n281), .B2(new_n284), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n315), .B1(new_n316), .B2(new_n309), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n268), .B1(new_n318), .B2(new_n252), .ZN(new_n319));
  AOI211_X1 g133(.A(G902), .B(new_n267), .C1(new_n314), .C2(new_n317), .ZN(new_n320));
  OR2_X1    g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n256), .A2(new_n265), .A3(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(KEYINPUT94), .ZN(new_n323));
  OAI21_X1  g137(.A(G221), .B1(new_n311), .B2(G902), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n201), .A2(G143), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n269), .A2(G146), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n201), .A2(G143), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n328), .A2(new_n274), .B1(KEYINPUT1), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n274), .A2(KEYINPUT1), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n326), .A3(new_n327), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT80), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT80), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n331), .A2(new_n326), .A3(new_n327), .A4(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n330), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(KEYINPUT3), .B1(new_n219), .B2(G107), .ZN(new_n337));
  AOI21_X1  g151(.A(G101), .B1(new_n219), .B2(G107), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n289), .A3(G104), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n337), .A2(new_n338), .A3(new_n340), .A4(KEYINPUT78), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n289), .A2(G104), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n219), .A2(G107), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G101), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n336), .A2(new_n345), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n330), .A2(new_n332), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n343), .A2(new_n344), .B1(G101), .B2(new_n348), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT11), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(new_n297), .B2(G137), .ZN(new_n356));
  INV_X1    g170(.A(G137), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(KEYINPUT11), .A3(G134), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n297), .A2(G137), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G131), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n356), .A2(new_n358), .A3(new_n197), .A4(new_n359), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n353), .A2(new_n354), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT12), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT12), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n353), .A2(new_n354), .A3(new_n366), .A4(new_n363), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(KEYINPUT0), .A2(G128), .ZN(new_n369));
  OR2_X1    g183(.A1(KEYINPUT0), .A2(G128), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n269), .A2(G146), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n369), .B(new_n370), .C1(new_n371), .C2(new_n329), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT0), .A4(G128), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n337), .A2(new_n340), .A3(new_n347), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT4), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(G101), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT79), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n376), .B1(new_n375), .B2(G101), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n345), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n380), .B1(new_n345), .B2(new_n381), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n379), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n363), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT10), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n386), .B1(new_n330), .B2(new_n332), .ZN(new_n387));
  AOI22_X1  g201(.A1(new_n350), .A2(new_n386), .B1(new_n352), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n384), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(G110), .B(G140), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n257), .A2(G227), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n391), .B(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n368), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n345), .A2(new_n381), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT79), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n345), .A2(new_n380), .A3(new_n381), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n378), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n350), .A2(new_n386), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n352), .A2(new_n387), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n363), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT83), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n384), .A2(new_n388), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(KEYINPUT83), .A3(new_n363), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n390), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n393), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n395), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G469), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(new_n252), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT84), .ZN(new_n413));
  AOI21_X1  g227(.A(KEYINPUT83), .B1(new_n406), .B2(new_n363), .ZN(new_n414));
  AOI211_X1 g228(.A(new_n404), .B(new_n385), .C1(new_n384), .C2(new_n388), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n389), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n393), .ZN(new_n417));
  AOI21_X1  g231(.A(G902), .B1(new_n417), .B2(new_n395), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT84), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(new_n411), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n413), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n365), .A2(new_n389), .A3(new_n367), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT82), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n365), .A2(new_n389), .A3(new_n367), .A4(KEYINPUT82), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n409), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI211_X1 g240(.A(new_n393), .B(new_n390), .C1(new_n405), .C2(new_n407), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G469), .B1(new_n428), .B2(G902), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n325), .B1(new_n421), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G214), .B1(G237), .B2(G902), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n431), .B(KEYINPUT85), .Z(new_n432));
  INV_X1    g246(.A(G119), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G116), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n303), .A2(G119), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(KEYINPUT2), .B(G113), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT65), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G113), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT2), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT2), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G113), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G116), .B(G119), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT65), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n438), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(KEYINPUT5), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n448), .B(G113), .C1(KEYINPUT5), .C2(new_n434), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n352), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT66), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n436), .A2(new_n437), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n447), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n451), .B1(new_n447), .B2(new_n452), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n377), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n382), .A2(new_n383), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n450), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G110), .B(G122), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n450), .B(new_n458), .C1(new_n455), .C2(new_n456), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(KEYINPUT6), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n457), .A2(new_n463), .A3(new_n459), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n374), .A2(new_n204), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n351), .A2(G125), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n257), .A2(G224), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n467), .B(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n462), .A2(new_n464), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(KEYINPUT7), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n471), .B1(new_n465), .B2(new_n466), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT86), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g288(.A(KEYINPUT86), .B(new_n471), .C1(new_n465), .C2(new_n466), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n458), .B(KEYINPUT8), .ZN(new_n477));
  INV_X1    g291(.A(new_n450), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n352), .B1(new_n447), .B2(new_n449), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n467), .A2(KEYINPUT7), .A3(new_n468), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n476), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(G902), .B1(new_n482), .B2(new_n461), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n470), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(G210), .B1(G237), .B2(G902), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n470), .A2(new_n483), .A3(new_n485), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n432), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n323), .A2(new_n430), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT95), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT95), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n323), .A2(new_n430), .A3(new_n492), .A4(new_n489), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n312), .B1(G234), .B2(new_n252), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n257), .A2(G221), .A3(G234), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(KEYINPUT75), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT22), .B(G137), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n498), .B(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n274), .A2(G119), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n433), .A2(G128), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT24), .B(G110), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT72), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT23), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT72), .B(KEYINPUT23), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n508), .B(new_n502), .C1(new_n509), .C2(new_n501), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n505), .B1(new_n510), .B2(G110), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n209), .A2(new_n201), .A3(new_n211), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n511), .B1(new_n512), .B2(new_n212), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT74), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT74), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n515), .B(new_n511), .C1(new_n512), .C2(new_n212), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n503), .A2(new_n504), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n433), .A2(G128), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT23), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(KEYINPUT72), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n502), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(KEYINPUT72), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n501), .B1(new_n507), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G110), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n518), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n223), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n527), .A2(new_n212), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n500), .B1(new_n517), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n500), .ZN(new_n532));
  AOI211_X1 g346(.A(new_n532), .B(new_n529), .C1(new_n514), .C2(new_n516), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT25), .B1(new_n534), .B2(new_n252), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT25), .ZN(new_n536));
  NOR4_X1   g350(.A1(new_n531), .A2(new_n533), .A3(new_n536), .A4(G902), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n496), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT76), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(KEYINPUT76), .B(new_n496), .C1(new_n535), .C2(new_n537), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n496), .A2(G902), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n534), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT77), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n540), .A2(KEYINPUT77), .A3(new_n541), .A4(new_n543), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(G472), .A2(G902), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n190), .A2(G210), .ZN(new_n550));
  XOR2_X1   g364(.A(new_n550), .B(KEYINPUT27), .Z(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT26), .B(G101), .ZN(new_n552));
  XOR2_X1   g366(.A(new_n551), .B(new_n552), .Z(new_n553));
  INV_X1    g367(.A(KEYINPUT68), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n554), .B1(new_n453), .B2(new_n454), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n436), .A2(new_n437), .A3(KEYINPUT65), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n445), .B1(new_n443), .B2(new_n444), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n452), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT66), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n447), .A2(new_n451), .A3(new_n452), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(KEYINPUT68), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT67), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n374), .A2(new_n363), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n374), .A2(new_n363), .ZN(new_n564));
  INV_X1    g378(.A(new_n359), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n297), .A2(G137), .ZN(new_n566));
  OAI21_X1  g380(.A(G131), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n567), .A2(new_n362), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n564), .A2(KEYINPUT67), .B1(new_n351), .B2(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n555), .A2(new_n561), .A3(new_n563), .A4(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT69), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n564), .A2(KEYINPUT67), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n568), .A2(new_n351), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n573), .A2(new_n563), .A3(new_n574), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n575), .A2(KEYINPUT69), .A3(new_n561), .A4(new_n555), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT64), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n564), .A2(new_n578), .B1(new_n351), .B2(new_n568), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n374), .A2(new_n363), .A3(KEYINPUT64), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n453), .A2(new_n454), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT28), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n555), .A2(new_n561), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n564), .A2(new_n574), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT28), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n553), .B1(new_n586), .B2(new_n590), .ZN(new_n591));
  AND4_X1   g405(.A1(KEYINPUT30), .A2(new_n573), .A3(new_n563), .A4(new_n574), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT30), .B1(new_n579), .B2(new_n580), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n559), .A2(new_n560), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n577), .A2(new_n596), .A3(new_n553), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT31), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n572), .A2(new_n576), .B1(new_n594), .B2(new_n595), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT31), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n600), .A3(new_n553), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n591), .A2(new_n602), .A3(KEYINPUT70), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT70), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n600), .B1(new_n599), .B2(new_n553), .ZN(new_n605));
  AND4_X1   g419(.A1(new_n600), .A2(new_n577), .A3(new_n596), .A4(new_n553), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n553), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n583), .B1(new_n572), .B2(new_n576), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT28), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n608), .B1(new_n611), .B2(new_n589), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n604), .B1(new_n607), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n549), .B1(new_n603), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT32), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(KEYINPUT70), .B1(new_n591), .B2(new_n602), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n612), .A2(new_n604), .A3(new_n598), .A4(new_n601), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n549), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n615), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT71), .ZN(new_n622));
  OAI22_X1  g436(.A1(new_n577), .A2(new_n622), .B1(new_n587), .B2(new_n575), .ZN(new_n623));
  AOI21_X1  g437(.A(KEYINPUT71), .B1(new_n572), .B2(new_n576), .ZN(new_n624));
  OAI21_X1  g438(.A(KEYINPUT28), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n553), .A2(KEYINPUT29), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(new_n590), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n577), .A2(new_n596), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT29), .B1(new_n628), .B2(new_n608), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n590), .B(new_n553), .C1(new_n609), .C2(new_n610), .ZN(new_n630));
  AOI21_X1  g444(.A(G902), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n619), .A2(new_n621), .B1(G472), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n548), .B1(new_n616), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n495), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G101), .ZN(G3));
  AOI21_X1  g450(.A(new_n620), .B1(new_n617), .B2(new_n618), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n252), .B1(new_n603), .B2(new_n613), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n637), .B1(new_n638), .B2(G472), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT96), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n546), .A2(new_n547), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n639), .A2(new_n640), .A3(new_n641), .A4(new_n430), .ZN(new_n642));
  AOI21_X1  g456(.A(G902), .B1(new_n617), .B2(new_n618), .ZN(new_n643));
  INV_X1    g457(.A(G472), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n614), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n419), .B1(new_n418), .B2(new_n411), .ZN(new_n646));
  AOI22_X1  g460(.A1(new_n416), .A2(new_n393), .B1(new_n368), .B2(new_n394), .ZN(new_n647));
  NOR4_X1   g461(.A1(new_n647), .A2(KEYINPUT84), .A3(G469), .A4(G902), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n429), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n546), .A2(new_n649), .A3(new_n547), .A4(new_n324), .ZN(new_n650));
  OAI21_X1  g464(.A(KEYINPUT96), .B1(new_n645), .B2(new_n650), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n642), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n431), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n487), .B2(new_n488), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n318), .A2(new_n266), .A3(new_n252), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n266), .A2(new_n252), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n316), .A2(new_n309), .ZN(new_n659));
  OAI21_X1  g473(.A(KEYINPUT33), .B1(new_n659), .B2(KEYINPUT97), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n318), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n318), .A2(new_n660), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n658), .B1(new_n663), .B2(G478), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n256), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n265), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n652), .A2(new_n654), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT98), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT34), .B(G104), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G6));
  INV_X1    g484(.A(new_n265), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n245), .B(new_n187), .C1(new_n249), .C2(new_n229), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n247), .A2(new_n672), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n673), .A2(new_n321), .A3(new_n255), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n654), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n652), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT35), .B(G107), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G9));
  NAND2_X1  g493(.A1(new_n517), .A2(new_n530), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n532), .A2(KEYINPUT36), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n542), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n540), .A2(new_n541), .A3(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT99), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n540), .A2(KEYINPUT99), .A3(new_n541), .A4(new_n683), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n645), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n495), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT37), .B(G110), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G12));
  NAND2_X1  g507(.A1(new_n649), .A2(new_n324), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n694), .B1(new_n686), .B2(new_n687), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n621), .B1(new_n603), .B2(new_n613), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n632), .A2(G472), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n696), .B(new_n697), .C1(KEYINPUT32), .C2(new_n637), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT100), .B(G900), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n263), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g514(.A1(new_n700), .A2(KEYINPUT101), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(KEYINPUT101), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n701), .A2(new_n261), .A3(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n674), .A2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n695), .A2(new_n698), .A3(new_n654), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G128), .ZN(G30));
  XOR2_X1   g522(.A(new_n703), .B(KEYINPUT39), .Z(new_n709));
  NAND2_X1  g523(.A1(new_n430), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT104), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n711), .A2(KEYINPUT40), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(KEYINPUT40), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n431), .B1(new_n319), .B2(new_n320), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(new_n251), .B2(new_n255), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n689), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT103), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n608), .B1(new_n623), .B2(new_n624), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(KEYINPUT102), .A3(new_n597), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n252), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT102), .B1(new_n718), .B2(new_n597), .ZN(new_n721));
  OAI21_X1  g535(.A(G472), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n696), .B(new_n722), .C1(KEYINPUT32), .C2(new_n637), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n487), .A2(new_n488), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT38), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n712), .A2(new_n713), .A3(new_n717), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT105), .B(G143), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G45));
  NOR2_X1   g545(.A1(new_n665), .A2(new_n703), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n616), .B2(new_n633), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n688), .A2(new_n430), .A3(new_n654), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G146), .ZN(G48));
  AOI21_X1  g551(.A(new_n411), .B1(new_n410), .B2(new_n252), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n421), .A2(new_n324), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n666), .A2(new_n654), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n634), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(KEYINPUT41), .B(G113), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(G15));
  NOR2_X1   g559(.A1(new_n740), .A2(new_n675), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n634), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G116), .ZN(G18));
  NAND4_X1  g562(.A1(new_n421), .A2(new_n324), .A3(new_n654), .A4(new_n739), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n698), .A2(new_n323), .A3(new_n750), .A4(new_n688), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G119), .ZN(G21));
  NAND3_X1  g566(.A1(new_n638), .A2(KEYINPUT106), .A3(G472), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT106), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n754), .B1(new_n643), .B2(new_n644), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  AOI211_X1 g570(.A(new_n325), .B(new_n738), .C1(new_n413), .C2(new_n420), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n470), .A2(new_n483), .A3(new_n485), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n485), .B1(new_n470), .B2(new_n483), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n715), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT107), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT107), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n725), .A2(new_n762), .A3(new_n715), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n757), .A2(new_n764), .A3(new_n671), .ZN(new_n765));
  INV_X1    g579(.A(new_n544), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n553), .B1(new_n625), .B2(new_n590), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n549), .B1(new_n767), .B2(new_n602), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n756), .A2(new_n765), .A3(new_n766), .A4(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G122), .ZN(G24));
  AOI21_X1  g584(.A(new_n749), .B1(new_n686), .B2(new_n687), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n756), .A2(new_n771), .A3(new_n732), .A4(new_n768), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G125), .ZN(G27));
  INV_X1    g587(.A(KEYINPUT42), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n696), .A2(new_n697), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT32), .B1(new_n619), .B2(new_n549), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n641), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n487), .A2(new_n488), .A3(new_n431), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT108), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT108), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n487), .A2(new_n780), .A3(new_n488), .A4(new_n431), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n430), .A3(new_n732), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n774), .B1(new_n777), .B2(new_n784), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n694), .A2(new_n782), .A3(new_n733), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n786), .A2(KEYINPUT42), .A3(new_n698), .A4(new_n766), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G131), .ZN(G33));
  NOR2_X1   g603(.A1(new_n694), .A2(new_n782), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n634), .A2(new_n706), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G134), .ZN(G36));
  OR2_X1    g606(.A1(new_n428), .A2(KEYINPUT45), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n428), .A2(KEYINPUT45), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(G469), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(G469), .A2(G902), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT46), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n421), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n795), .A2(KEYINPUT46), .A3(new_n796), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n325), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n709), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n256), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n664), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT43), .Z(new_n806));
  NAND3_X1  g620(.A1(new_n645), .A2(new_n806), .A3(new_n688), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT44), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n782), .B(KEYINPUT109), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n803), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G137), .ZN(G39));
  XOR2_X1   g625(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n812));
  AND2_X1   g626(.A1(new_n801), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT110), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(KEYINPUT47), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n801), .A2(new_n815), .ZN(new_n816));
  OR4_X1    g630(.A1(new_n698), .A2(new_n641), .A3(new_n733), .A4(new_n782), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n813), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(new_n202), .ZN(G42));
  NOR2_X1   g633(.A1(new_n798), .A2(new_n738), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(KEYINPUT49), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(KEYINPUT111), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n805), .A2(new_n325), .A3(new_n432), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n727), .A2(new_n824), .A3(new_n766), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n825), .B1(KEYINPUT49), .B2(new_n821), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n823), .A2(new_n724), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n783), .A2(new_n757), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT119), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(new_n641), .A3(new_n262), .A4(new_n724), .ZN(new_n830));
  OR3_X1    g644(.A1(new_n830), .A2(new_n256), .A3(new_n664), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n756), .A2(new_n768), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n806), .A2(new_n262), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n829), .A2(new_n688), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(KEYINPUT120), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n832), .A2(new_n766), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n833), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n740), .A2(new_n431), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n839), .A2(KEYINPUT117), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(KEYINPUT117), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n840), .A2(new_n727), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  XOR2_X1   g657(.A(KEYINPUT118), .B(KEYINPUT50), .Z(new_n844));
  OR2_X1    g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n843), .B1(KEYINPUT118), .B2(KEYINPUT50), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI22_X1  g661(.A1(new_n813), .A2(new_n816), .B1(new_n324), .B2(new_n821), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(new_n837), .A3(new_n809), .A4(new_n833), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n836), .A2(KEYINPUT51), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n698), .A2(new_n829), .A3(new_n766), .A4(new_n833), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT48), .ZN(new_n852));
  OAI221_X1 g666(.A(new_n258), .B1(new_n830), .B2(new_n665), .C1(new_n838), .C2(new_n749), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AND4_X1   g668(.A1(new_n847), .A2(new_n849), .A3(new_n834), .A4(new_n831), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n850), .B(new_n854), .C1(new_n855), .C2(KEYINPUT51), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT113), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n673), .A2(new_n255), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n859), .A2(new_n321), .A3(new_n703), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n779), .A2(new_n781), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n862), .B1(new_n775), .B2(new_n776), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n688), .A2(new_n430), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n858), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n861), .B1(new_n616), .B2(new_n633), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n866), .A2(KEYINPUT113), .A3(new_n695), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n777), .A2(new_n705), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n865), .A2(new_n867), .B1(new_n868), .B2(new_n790), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n698), .B(new_n641), .C1(new_n742), .C2(new_n746), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n769), .A2(new_n751), .A3(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n756), .A2(new_n786), .A3(new_n688), .A4(new_n768), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n869), .A2(new_n871), .A3(new_n788), .A4(new_n872), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n493), .B(new_n491), .C1(new_n690), .C2(new_n634), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n666), .A2(new_n489), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n642), .A2(new_n651), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n489), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n804), .A2(new_n671), .A3(new_n321), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT112), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n642), .A2(new_n651), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n874), .A2(new_n876), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT114), .B1(new_n873), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n684), .A2(new_n703), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n723), .A2(new_n430), .A3(new_n764), .A4(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n772), .A2(new_n707), .A3(new_n736), .A4(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT52), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n735), .B(new_n698), .C1(new_n706), .C2(new_n732), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n889), .A2(new_n772), .A3(KEYINPUT52), .A4(new_n885), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n863), .A2(new_n858), .A3(new_n864), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT113), .B1(new_n866), .B2(new_n695), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n791), .B(new_n872), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  AOI211_X1 g709(.A(new_n774), .B(new_n544), .C1(new_n616), .C2(new_n633), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n786), .A2(new_n698), .A3(new_n641), .ZN(new_n897));
  AOI22_X1  g711(.A1(new_n786), .A2(new_n896), .B1(new_n897), .B2(new_n774), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n769), .A2(new_n751), .A3(new_n870), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n882), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT114), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n895), .A2(new_n900), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n883), .A2(new_n891), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n891), .A2(KEYINPUT53), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n895), .A2(new_n900), .A3(new_n901), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT116), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n870), .A2(new_n751), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n788), .A2(new_n908), .A3(new_n769), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n909), .A2(new_n894), .A3(new_n882), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT116), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n857), .B1(new_n888), .B2(new_n890), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI22_X1  g727(.A1(new_n857), .A2(new_n904), .B1(new_n907), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT54), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT53), .B1(new_n891), .B2(KEYINPUT115), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n904), .B(new_n917), .Z(new_n918));
  OAI21_X1  g732(.A(new_n916), .B1(new_n918), .B2(new_n915), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n856), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(G952), .A2(G953), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n827), .B1(new_n920), .B2(new_n921), .ZN(G75));
  NOR2_X1   g736(.A1(new_n914), .A2(new_n252), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(G210), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n462), .A2(new_n464), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(new_n469), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT55), .Z(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT121), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n929), .A2(KEYINPUT56), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n924), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n928), .B1(new_n924), .B2(new_n930), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n257), .A2(G952), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(G51));
  XNOR2_X1  g748(.A(new_n914), .B(KEYINPUT54), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n796), .B(KEYINPUT57), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n410), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OR3_X1    g751(.A1(new_n914), .A2(new_n252), .A3(new_n795), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n933), .B1(new_n937), .B2(new_n938), .ZN(G54));
  NAND3_X1  g753(.A1(new_n923), .A2(KEYINPUT58), .A3(G475), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n940), .A2(new_n244), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n940), .A2(new_n244), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n941), .A2(new_n942), .A3(new_n933), .ZN(G60));
  INV_X1    g757(.A(new_n663), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n656), .B(KEYINPUT59), .Z(new_n945));
  AOI21_X1  g759(.A(new_n944), .B1(new_n919), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n933), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n944), .A2(new_n945), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n947), .B1(new_n935), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n946), .A2(new_n949), .ZN(G63));
  INV_X1    g764(.A(new_n534), .ZN(new_n951));
  NAND2_X1  g765(.A1(G217), .A2(G902), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT60), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n914), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n953), .ZN(new_n955));
  AOI22_X1  g769(.A1(new_n906), .A2(KEYINPUT114), .B1(new_n888), .B2(new_n890), .ZN(new_n956));
  AOI21_X1  g770(.A(KEYINPUT53), .B1(new_n956), .B2(new_n903), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n911), .B1(new_n910), .B2(new_n912), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n682), .B(new_n955), .C1(new_n957), .C2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n954), .A2(new_n947), .A3(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT122), .ZN(new_n963));
  XNOR2_X1  g777(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n964), .B1(new_n962), .B2(new_n963), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(G66));
  INV_X1    g781(.A(G224), .ZN(new_n968));
  OAI21_X1  g782(.A(G953), .B1(new_n264), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n882), .A2(new_n899), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n969), .B1(new_n970), .B2(G953), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n925), .B1(G898), .B2(new_n257), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(G69));
  NAND4_X1  g787(.A1(new_n803), .A2(new_n698), .A3(new_n766), .A4(new_n764), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n974), .A2(new_n788), .A3(new_n791), .ZN(new_n975));
  INV_X1    g789(.A(new_n810), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n976), .A2(new_n818), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n889), .A2(new_n772), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n975), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT126), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n979), .A2(new_n980), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n981), .A2(new_n257), .A3(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n236), .A2(new_n237), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n594), .B(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n985), .B1(G900), .B2(G953), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n729), .A2(new_n978), .ZN(new_n988));
  OR2_X1    g802(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n804), .A2(new_n321), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n991), .A2(new_n665), .ZN(new_n992));
  NOR4_X1   g806(.A1(new_n711), .A2(new_n777), .A3(new_n782), .A4(new_n992), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n976), .A2(new_n818), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n989), .A2(new_n990), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n257), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n985), .B(KEYINPUT124), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n987), .A2(KEYINPUT125), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n257), .B1(G227), .B2(G900), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1000), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n987), .A2(new_n998), .A3(KEYINPUT125), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1001), .A2(new_n1003), .ZN(G72));
  NAND3_X1  g818(.A1(new_n981), .A2(new_n970), .A3(new_n982), .ZN(new_n1005));
  XNOR2_X1  g819(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n644), .A2(new_n252), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  AOI211_X1 g822(.A(new_n553), .B(new_n628), .C1(new_n1005), .C2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n970), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1008), .B1(new_n995), .B2(new_n1010), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n1011), .A2(new_n553), .A3(new_n628), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n599), .A2(new_n553), .ZN(new_n1013));
  INV_X1    g827(.A(new_n597), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1008), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n918), .A2(new_n1015), .ZN(new_n1016));
  NOR4_X1   g830(.A1(new_n1009), .A2(new_n933), .A3(new_n1012), .A4(new_n1016), .ZN(G57));
endmodule


