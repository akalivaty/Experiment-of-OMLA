

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U547 ( .A1(n714), .A2(n707), .ZN(n709) );
  NOR2_X1 U548 ( .A1(G2104), .A2(G2105), .ZN(n549) );
  NAND2_X1 U549 ( .A1(G29), .A2(n968), .ZN(n512) );
  OR2_X1 U550 ( .A1(n788), .A2(n787), .ZN(n513) );
  AND2_X1 U551 ( .A1(n791), .A2(n790), .ZN(n514) );
  INV_X1 U552 ( .A(n973), .ZN(n705) );
  INV_X1 U553 ( .A(KEYINPUT96), .ZN(n708) );
  INV_X1 U554 ( .A(n747), .ZN(n720) );
  BUF_X1 U555 ( .A(n720), .Z(n733) );
  NOR2_X1 U556 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U557 ( .A(n755), .B(KEYINPUT32), .ZN(n763) );
  NAND2_X1 U558 ( .A1(n763), .A2(n762), .ZN(n765) );
  AND2_X1 U559 ( .A1(n789), .A2(n513), .ZN(n790) );
  NOR2_X1 U560 ( .A1(G164), .A2(G1384), .ZN(n700) );
  AND2_X1 U561 ( .A1(n822), .A2(n833), .ZN(n824) );
  XNOR2_X1 U562 ( .A(n619), .B(n618), .ZN(n970) );
  INV_X1 U563 ( .A(KEYINPUT17), .ZN(n548) );
  AND2_X1 U564 ( .A1(n824), .A2(n823), .ZN(n825) );
  BUF_X1 U565 ( .A(n521), .Z(n646) );
  NAND2_X1 U566 ( .A1(n905), .A2(G138), .ZN(n588) );
  NOR2_X2 U567 ( .A1(G2104), .A2(n540), .ZN(n897) );
  NOR2_X1 U568 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U569 ( .A1(n610), .A2(n609), .ZN(n973) );
  NOR2_X1 U570 ( .A1(G651), .A2(G543), .ZN(n652) );
  NAND2_X1 U571 ( .A1(n652), .A2(G89), .ZN(n515) );
  XNOR2_X1 U572 ( .A(n515), .B(KEYINPUT4), .ZN(n517) );
  XOR2_X1 U573 ( .A(KEYINPUT0), .B(G543), .Z(n521) );
  INV_X1 U574 ( .A(G651), .ZN(n519) );
  NOR2_X1 U575 ( .A1(n521), .A2(n519), .ZN(n657) );
  NAND2_X1 U576 ( .A1(G76), .A2(n657), .ZN(n516) );
  NAND2_X1 U577 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U578 ( .A(KEYINPUT5), .B(n518), .ZN(n527) );
  NOR2_X1 U579 ( .A1(G543), .A2(n519), .ZN(n520) );
  XOR2_X2 U580 ( .A(KEYINPUT1), .B(n520), .Z(n653) );
  NAND2_X1 U581 ( .A1(G63), .A2(n653), .ZN(n523) );
  NOR2_X2 U582 ( .A1(G651), .A2(n646), .ZN(n662) );
  NAND2_X1 U583 ( .A1(G51), .A2(n662), .ZN(n522) );
  NAND2_X1 U584 ( .A1(n523), .A2(n522), .ZN(n525) );
  XOR2_X1 U585 ( .A(KEYINPUT76), .B(KEYINPUT6), .Z(n524) );
  XNOR2_X1 U586 ( .A(n525), .B(n524), .ZN(n526) );
  NAND2_X1 U587 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U588 ( .A(KEYINPUT7), .B(n528), .ZN(G168) );
  XOR2_X1 U589 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U590 ( .A1(G91), .A2(n652), .ZN(n529) );
  XOR2_X1 U591 ( .A(KEYINPUT68), .B(n529), .Z(n534) );
  NAND2_X1 U592 ( .A1(G65), .A2(n653), .ZN(n531) );
  NAND2_X1 U593 ( .A1(G53), .A2(n662), .ZN(n530) );
  NAND2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U595 ( .A(KEYINPUT69), .B(n532), .Z(n533) );
  NOR2_X1 U596 ( .A1(n534), .A2(n533), .ZN(n536) );
  NAND2_X1 U597 ( .A1(n657), .A2(G78), .ZN(n535) );
  NAND2_X1 U598 ( .A1(n536), .A2(n535), .ZN(G299) );
  INV_X1 U599 ( .A(KEYINPUT23), .ZN(n539) );
  INV_X1 U600 ( .A(G2105), .ZN(n537) );
  AND2_X1 U601 ( .A1(n537), .A2(G2104), .ZN(n902) );
  NAND2_X1 U602 ( .A1(n902), .A2(G101), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(n544) );
  INV_X1 U604 ( .A(G2105), .ZN(n540) );
  NAND2_X1 U605 ( .A1(n897), .A2(G125), .ZN(n543) );
  AND2_X1 U606 ( .A1(n544), .A2(n543), .ZN(n542) );
  INV_X1 U607 ( .A(KEYINPUT65), .ZN(n541) );
  NAND2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n547) );
  NAND2_X1 U609 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U610 ( .A1(n545), .A2(KEYINPUT65), .ZN(n546) );
  NAND2_X1 U611 ( .A1(n547), .A2(n546), .ZN(n696) );
  XNOR2_X2 U612 ( .A(n549), .B(n548), .ZN(n905) );
  NAND2_X1 U613 ( .A1(G137), .A2(n905), .ZN(n691) );
  AND2_X1 U614 ( .A1(n696), .A2(n691), .ZN(n551) );
  AND2_X1 U615 ( .A1(G2104), .A2(G2105), .ZN(n898) );
  NAND2_X1 U616 ( .A1(G113), .A2(n898), .ZN(n550) );
  XNOR2_X1 U617 ( .A(KEYINPUT66), .B(n550), .ZN(n690) );
  AND2_X1 U618 ( .A1(n551), .A2(n690), .ZN(G160) );
  NAND2_X1 U619 ( .A1(G85), .A2(n652), .ZN(n553) );
  NAND2_X1 U620 ( .A1(G72), .A2(n657), .ZN(n552) );
  NAND2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n557) );
  NAND2_X1 U622 ( .A1(G60), .A2(n653), .ZN(n555) );
  NAND2_X1 U623 ( .A1(G47), .A2(n662), .ZN(n554) );
  NAND2_X1 U624 ( .A1(n555), .A2(n554), .ZN(n556) );
  OR2_X1 U625 ( .A1(n557), .A2(n556), .ZN(G290) );
  XOR2_X1 U626 ( .A(KEYINPUT107), .B(KEYINPUT109), .Z(n559) );
  XNOR2_X1 U627 ( .A(G2446), .B(G2451), .ZN(n558) );
  XNOR2_X1 U628 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U629 ( .A(n560), .B(G2430), .Z(n562) );
  XNOR2_X1 U630 ( .A(G1348), .B(G1341), .ZN(n561) );
  XNOR2_X1 U631 ( .A(n562), .B(n561), .ZN(n566) );
  XOR2_X1 U632 ( .A(KEYINPUT108), .B(G2435), .Z(n564) );
  XNOR2_X1 U633 ( .A(G2438), .B(G2454), .ZN(n563) );
  XNOR2_X1 U634 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U635 ( .A(n566), .B(n565), .Z(n568) );
  XNOR2_X1 U636 ( .A(G2443), .B(G2427), .ZN(n567) );
  XNOR2_X1 U637 ( .A(n568), .B(n567), .ZN(n569) );
  AND2_X1 U638 ( .A1(n569), .A2(G14), .ZN(G401) );
  NAND2_X1 U639 ( .A1(G90), .A2(n652), .ZN(n571) );
  NAND2_X1 U640 ( .A1(G77), .A2(n657), .ZN(n570) );
  NAND2_X1 U641 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U642 ( .A(n572), .B(KEYINPUT9), .ZN(n574) );
  NAND2_X1 U643 ( .A1(G52), .A2(n662), .ZN(n573) );
  NAND2_X1 U644 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U645 ( .A1(G64), .A2(n653), .ZN(n575) );
  XNOR2_X1 U646 ( .A(KEYINPUT67), .B(n575), .ZN(n576) );
  NOR2_X1 U647 ( .A1(n577), .A2(n576), .ZN(G171) );
  AND2_X1 U648 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U649 ( .A1(G135), .A2(n905), .ZN(n584) );
  NAND2_X1 U650 ( .A1(G99), .A2(n902), .ZN(n579) );
  NAND2_X1 U651 ( .A1(G111), .A2(n898), .ZN(n578) );
  NAND2_X1 U652 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U653 ( .A1(n897), .A2(G123), .ZN(n580) );
  XOR2_X1 U654 ( .A(KEYINPUT18), .B(n580), .Z(n581) );
  NOR2_X1 U655 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U656 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U657 ( .A(n585), .B(KEYINPUT80), .ZN(n951) );
  XNOR2_X1 U658 ( .A(n951), .B(G2096), .ZN(n586) );
  OR2_X1 U659 ( .A1(G2100), .A2(n586), .ZN(G156) );
  NAND2_X1 U660 ( .A1(G102), .A2(n902), .ZN(n587) );
  NAND2_X1 U661 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U662 ( .A1(G126), .A2(n897), .ZN(n590) );
  NAND2_X1 U663 ( .A1(G114), .A2(n898), .ZN(n589) );
  NAND2_X1 U664 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U665 ( .A1(n592), .A2(n591), .ZN(G164) );
  INV_X1 U666 ( .A(G132), .ZN(G219) );
  INV_X1 U667 ( .A(G82), .ZN(G220) );
  INV_X1 U668 ( .A(G57), .ZN(G237) );
  INV_X1 U669 ( .A(G108), .ZN(G238) );
  INV_X1 U670 ( .A(G120), .ZN(G236) );
  NAND2_X1 U671 ( .A1(G88), .A2(n652), .ZN(n594) );
  NAND2_X1 U672 ( .A1(G75), .A2(n657), .ZN(n593) );
  NAND2_X1 U673 ( .A1(n594), .A2(n593), .ZN(n598) );
  NAND2_X1 U674 ( .A1(G62), .A2(n653), .ZN(n596) );
  NAND2_X1 U675 ( .A1(G50), .A2(n662), .ZN(n595) );
  NAND2_X1 U676 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U677 ( .A1(n598), .A2(n597), .ZN(G166) );
  NAND2_X1 U678 ( .A1(G7), .A2(G661), .ZN(n599) );
  XNOR2_X1 U679 ( .A(n599), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U680 ( .A(G223), .ZN(n844) );
  NAND2_X1 U681 ( .A1(n844), .A2(G567), .ZN(n600) );
  XOR2_X1 U682 ( .A(KEYINPUT11), .B(n600), .Z(G234) );
  NAND2_X1 U683 ( .A1(n652), .A2(G81), .ZN(n601) );
  XNOR2_X1 U684 ( .A(n601), .B(KEYINPUT12), .ZN(n603) );
  NAND2_X1 U685 ( .A1(G68), .A2(n657), .ZN(n602) );
  NAND2_X1 U686 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U687 ( .A(KEYINPUT13), .B(n604), .ZN(n610) );
  NAND2_X1 U688 ( .A1(G56), .A2(n653), .ZN(n605) );
  XOR2_X1 U689 ( .A(KEYINPUT14), .B(n605), .Z(n608) );
  NAND2_X1 U690 ( .A1(n662), .A2(G43), .ZN(n606) );
  XOR2_X1 U691 ( .A(KEYINPUT70), .B(n606), .Z(n607) );
  XNOR2_X1 U692 ( .A(G860), .B(KEYINPUT71), .ZN(n626) );
  OR2_X1 U693 ( .A1(n973), .A2(n626), .ZN(G153) );
  XOR2_X1 U694 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  NAND2_X1 U695 ( .A1(G868), .A2(G301), .ZN(n611) );
  XNOR2_X1 U696 ( .A(n611), .B(KEYINPUT73), .ZN(n621) );
  NAND2_X1 U697 ( .A1(G92), .A2(n652), .ZN(n613) );
  NAND2_X1 U698 ( .A1(n657), .A2(G79), .ZN(n612) );
  NAND2_X1 U699 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U700 ( .A1(G66), .A2(n653), .ZN(n615) );
  NAND2_X1 U701 ( .A1(G54), .A2(n662), .ZN(n614) );
  NAND2_X1 U702 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U703 ( .A1(n617), .A2(n616), .ZN(n619) );
  XNOR2_X1 U704 ( .A(KEYINPUT74), .B(KEYINPUT15), .ZN(n618) );
  INV_X1 U705 ( .A(n970), .ZN(n704) );
  NOR2_X1 U706 ( .A1(n704), .A2(G868), .ZN(n620) );
  NOR2_X1 U707 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U708 ( .A(KEYINPUT75), .B(n622), .ZN(G284) );
  INV_X1 U709 ( .A(G868), .ZN(n673) );
  NOR2_X1 U710 ( .A1(G286), .A2(n673), .ZN(n624) );
  NOR2_X1 U711 ( .A1(G868), .A2(G299), .ZN(n623) );
  NOR2_X1 U712 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U713 ( .A(KEYINPUT77), .B(n625), .Z(G297) );
  NAND2_X1 U714 ( .A1(n626), .A2(G559), .ZN(n627) );
  NAND2_X1 U715 ( .A1(n627), .A2(n704), .ZN(n628) );
  XNOR2_X1 U716 ( .A(n628), .B(KEYINPUT16), .ZN(n629) );
  XNOR2_X1 U717 ( .A(KEYINPUT78), .B(n629), .ZN(G148) );
  NOR2_X1 U718 ( .A1(G868), .A2(n973), .ZN(n632) );
  NAND2_X1 U719 ( .A1(n704), .A2(G868), .ZN(n630) );
  NOR2_X1 U720 ( .A1(G559), .A2(n630), .ZN(n631) );
  NOR2_X1 U721 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U722 ( .A(KEYINPUT79), .B(n633), .Z(G282) );
  NAND2_X1 U723 ( .A1(G80), .A2(n657), .ZN(n634) );
  XNOR2_X1 U724 ( .A(n634), .B(KEYINPUT82), .ZN(n641) );
  NAND2_X1 U725 ( .A1(G93), .A2(n652), .ZN(n636) );
  NAND2_X1 U726 ( .A1(G55), .A2(n662), .ZN(n635) );
  NAND2_X1 U727 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U728 ( .A1(G67), .A2(n653), .ZN(n637) );
  XNOR2_X1 U729 ( .A(KEYINPUT83), .B(n637), .ZN(n638) );
  NOR2_X1 U730 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U731 ( .A1(n641), .A2(n640), .ZN(n672) );
  XNOR2_X1 U732 ( .A(n973), .B(KEYINPUT81), .ZN(n643) );
  NAND2_X1 U733 ( .A1(n704), .A2(G559), .ZN(n642) );
  XOR2_X1 U734 ( .A(n643), .B(n642), .Z(n670) );
  NOR2_X1 U735 ( .A1(G860), .A2(n670), .ZN(n644) );
  XOR2_X1 U736 ( .A(n672), .B(n644), .Z(G145) );
  NAND2_X1 U737 ( .A1(G49), .A2(n662), .ZN(n645) );
  XNOR2_X1 U738 ( .A(n645), .B(KEYINPUT84), .ZN(n651) );
  NAND2_X1 U739 ( .A1(G87), .A2(n646), .ZN(n648) );
  NAND2_X1 U740 ( .A1(G74), .A2(G651), .ZN(n647) );
  NAND2_X1 U741 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U742 ( .A1(n653), .A2(n649), .ZN(n650) );
  NAND2_X1 U743 ( .A1(n651), .A2(n650), .ZN(G288) );
  NAND2_X1 U744 ( .A1(G86), .A2(n652), .ZN(n655) );
  NAND2_X1 U745 ( .A1(G61), .A2(n653), .ZN(n654) );
  NAND2_X1 U746 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U747 ( .A(KEYINPUT85), .B(n656), .Z(n660) );
  NAND2_X1 U748 ( .A1(n657), .A2(G73), .ZN(n658) );
  XOR2_X1 U749 ( .A(KEYINPUT2), .B(n658), .Z(n659) );
  NOR2_X1 U750 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U751 ( .A(n661), .B(KEYINPUT86), .ZN(n664) );
  NAND2_X1 U752 ( .A1(G48), .A2(n662), .ZN(n663) );
  NAND2_X1 U753 ( .A1(n664), .A2(n663), .ZN(G305) );
  XOR2_X1 U754 ( .A(G299), .B(G290), .Z(n665) );
  XNOR2_X1 U755 ( .A(n665), .B(G288), .ZN(n666) );
  XNOR2_X1 U756 ( .A(n672), .B(n666), .ZN(n668) );
  XNOR2_X1 U757 ( .A(G166), .B(KEYINPUT19), .ZN(n667) );
  XNOR2_X1 U758 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U759 ( .A(n669), .B(G305), .ZN(n913) );
  XOR2_X1 U760 ( .A(n670), .B(n913), .Z(n671) );
  NAND2_X1 U761 ( .A1(n671), .A2(G868), .ZN(n675) );
  NAND2_X1 U762 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U763 ( .A1(n675), .A2(n674), .ZN(G295) );
  NAND2_X1 U764 ( .A1(G2078), .A2(G2084), .ZN(n676) );
  XOR2_X1 U765 ( .A(KEYINPUT20), .B(n676), .Z(n677) );
  NAND2_X1 U766 ( .A1(G2090), .A2(n677), .ZN(n678) );
  XNOR2_X1 U767 ( .A(KEYINPUT21), .B(n678), .ZN(n679) );
  NAND2_X1 U768 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U769 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U770 ( .A1(G661), .A2(G483), .ZN(n688) );
  NOR2_X1 U771 ( .A1(G236), .A2(G238), .ZN(n680) );
  NAND2_X1 U772 ( .A1(G69), .A2(n680), .ZN(n681) );
  NOR2_X1 U773 ( .A1(n681), .A2(G237), .ZN(n682) );
  XNOR2_X1 U774 ( .A(n682), .B(KEYINPUT87), .ZN(n848) );
  NAND2_X1 U775 ( .A1(n848), .A2(G567), .ZN(n687) );
  NOR2_X1 U776 ( .A1(G220), .A2(G219), .ZN(n683) );
  XOR2_X1 U777 ( .A(KEYINPUT22), .B(n683), .Z(n684) );
  NOR2_X1 U778 ( .A1(G218), .A2(n684), .ZN(n685) );
  NAND2_X1 U779 ( .A1(G96), .A2(n685), .ZN(n849) );
  NAND2_X1 U780 ( .A1(n849), .A2(G2106), .ZN(n686) );
  NAND2_X1 U781 ( .A1(n687), .A2(n686), .ZN(n850) );
  NOR2_X1 U782 ( .A1(n688), .A2(n850), .ZN(n689) );
  XNOR2_X1 U783 ( .A(n689), .B(KEYINPUT88), .ZN(n847) );
  NAND2_X1 U784 ( .A1(G36), .A2(n847), .ZN(G176) );
  INV_X1 U785 ( .A(G166), .ZN(G303) );
  INV_X1 U786 ( .A(KEYINPUT26), .ZN(n703) );
  AND2_X1 U787 ( .A1(n690), .A2(G40), .ZN(n692) );
  AND2_X1 U788 ( .A1(n692), .A2(n691), .ZN(n694) );
  NAND2_X1 U789 ( .A1(n696), .A2(n694), .ZN(n810) );
  NAND2_X1 U790 ( .A1(n810), .A2(KEYINPUT93), .ZN(n698) );
  INV_X1 U791 ( .A(KEYINPUT93), .ZN(n693) );
  AND2_X1 U792 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U793 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U794 ( .A1(n698), .A2(n697), .ZN(n701) );
  XNOR2_X1 U795 ( .A(n700), .B(KEYINPUT64), .ZN(n809) );
  NAND2_X2 U796 ( .A1(n701), .A2(n809), .ZN(n747) );
  NAND2_X1 U797 ( .A1(G1996), .A2(n720), .ZN(n702) );
  XNOR2_X1 U798 ( .A(n703), .B(n702), .ZN(n714) );
  NAND2_X1 U799 ( .A1(G1341), .A2(n747), .ZN(n715) );
  AND2_X1 U800 ( .A1(n704), .A2(n715), .ZN(n706) );
  NAND2_X1 U801 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U802 ( .A(n709), .B(n708), .ZN(n713) );
  NOR2_X1 U803 ( .A1(n733), .A2(G1348), .ZN(n711) );
  NOR2_X1 U804 ( .A1(G2067), .A2(n747), .ZN(n710) );
  NOR2_X1 U805 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U806 ( .A1(n713), .A2(n712), .ZN(n719) );
  NOR2_X1 U807 ( .A1(n973), .A2(n714), .ZN(n716) );
  NAND2_X1 U808 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U809 ( .A1(n970), .A2(n717), .ZN(n718) );
  NAND2_X1 U810 ( .A1(n719), .A2(n718), .ZN(n725) );
  NAND2_X1 U811 ( .A1(n720), .A2(G2072), .ZN(n721) );
  XNOR2_X1 U812 ( .A(n721), .B(KEYINPUT27), .ZN(n723) );
  INV_X1 U813 ( .A(G1956), .ZN(n1006) );
  NOR2_X1 U814 ( .A1(n1006), .A2(n733), .ZN(n722) );
  OR2_X1 U815 ( .A1(n723), .A2(n722), .ZN(n727) );
  OR2_X1 U816 ( .A1(G299), .A2(n727), .ZN(n724) );
  NAND2_X1 U817 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U818 ( .A(n726), .B(KEYINPUT97), .ZN(n731) );
  XNOR2_X1 U819 ( .A(KEYINPUT28), .B(KEYINPUT95), .ZN(n729) );
  NAND2_X1 U820 ( .A1(n727), .A2(G299), .ZN(n728) );
  XNOR2_X1 U821 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U822 ( .A(n732), .B(KEYINPUT29), .ZN(n737) );
  OR2_X1 U823 ( .A1(n733), .A2(G1961), .ZN(n735) );
  XNOR2_X1 U824 ( .A(G2078), .B(KEYINPUT25), .ZN(n931) );
  NAND2_X1 U825 ( .A1(n733), .A2(n931), .ZN(n734) );
  NAND2_X1 U826 ( .A1(n735), .A2(n734), .ZN(n741) );
  NAND2_X1 U827 ( .A1(G171), .A2(n741), .ZN(n736) );
  NAND2_X1 U828 ( .A1(n737), .A2(n736), .ZN(n746) );
  NAND2_X1 U829 ( .A1(G8), .A2(n747), .ZN(n788) );
  NOR2_X1 U830 ( .A1(G1966), .A2(n788), .ZN(n761) );
  NOR2_X1 U831 ( .A1(G2084), .A2(n747), .ZN(n756) );
  NOR2_X1 U832 ( .A1(n761), .A2(n756), .ZN(n738) );
  NAND2_X1 U833 ( .A1(G8), .A2(n738), .ZN(n739) );
  XNOR2_X1 U834 ( .A(KEYINPUT30), .B(n739), .ZN(n740) );
  NOR2_X1 U835 ( .A1(G168), .A2(n740), .ZN(n743) );
  NOR2_X1 U836 ( .A1(G171), .A2(n741), .ZN(n742) );
  NOR2_X1 U837 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U838 ( .A(KEYINPUT31), .B(n744), .Z(n745) );
  NAND2_X1 U839 ( .A1(n746), .A2(n745), .ZN(n758) );
  NAND2_X1 U840 ( .A1(n758), .A2(G286), .ZN(n753) );
  NOR2_X1 U841 ( .A1(G1971), .A2(n788), .ZN(n749) );
  NOR2_X1 U842 ( .A1(G2090), .A2(n747), .ZN(n748) );
  NOR2_X1 U843 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U844 ( .A1(n750), .A2(G303), .ZN(n751) );
  XNOR2_X1 U845 ( .A(n751), .B(KEYINPUT98), .ZN(n752) );
  NAND2_X1 U846 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U847 ( .A1(n754), .A2(G8), .ZN(n755) );
  NAND2_X1 U848 ( .A1(G8), .A2(n756), .ZN(n757) );
  XNOR2_X1 U849 ( .A(n757), .B(KEYINPUT94), .ZN(n759) );
  NAND2_X1 U850 ( .A1(n759), .A2(n758), .ZN(n760) );
  OR2_X1 U851 ( .A1(n761), .A2(n760), .ZN(n762) );
  INV_X1 U852 ( .A(KEYINPUT99), .ZN(n764) );
  XNOR2_X1 U853 ( .A(n765), .B(n764), .ZN(n783) );
  NOR2_X1 U854 ( .A1(G1971), .A2(G303), .ZN(n766) );
  NOR2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n974) );
  NOR2_X1 U856 ( .A1(n766), .A2(n974), .ZN(n768) );
  INV_X1 U857 ( .A(n788), .ZN(n772) );
  NAND2_X1 U858 ( .A1(n974), .A2(n772), .ZN(n767) );
  NAND2_X1 U859 ( .A1(n767), .A2(KEYINPUT33), .ZN(n770) );
  AND2_X1 U860 ( .A1(n768), .A2(n770), .ZN(n769) );
  AND2_X1 U861 ( .A1(n783), .A2(n769), .ZN(n777) );
  INV_X1 U862 ( .A(n770), .ZN(n775) );
  INV_X1 U863 ( .A(KEYINPUT33), .ZN(n771) );
  NAND2_X1 U864 ( .A1(G1976), .A2(G288), .ZN(n976) );
  AND2_X1 U865 ( .A1(n771), .A2(n976), .ZN(n773) );
  AND2_X1 U866 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U867 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U868 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U869 ( .A(n778), .B(KEYINPUT100), .ZN(n780) );
  XNOR2_X1 U870 ( .A(KEYINPUT101), .B(G1981), .ZN(n779) );
  XNOR2_X1 U871 ( .A(n779), .B(G305), .ZN(n989) );
  NAND2_X1 U872 ( .A1(n780), .A2(n989), .ZN(n791) );
  NOR2_X1 U873 ( .A1(G2090), .A2(G303), .ZN(n781) );
  NAND2_X1 U874 ( .A1(G8), .A2(n781), .ZN(n782) );
  NAND2_X1 U875 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U876 ( .A1(n784), .A2(n788), .ZN(n785) );
  XNOR2_X1 U877 ( .A(n785), .B(KEYINPUT102), .ZN(n789) );
  NOR2_X1 U878 ( .A1(G1981), .A2(G305), .ZN(n786) );
  XOR2_X1 U879 ( .A(n786), .B(KEYINPUT24), .Z(n787) );
  XNOR2_X1 U880 ( .A(n514), .B(KEYINPUT103), .ZN(n826) );
  NAND2_X1 U881 ( .A1(G105), .A2(n902), .ZN(n792) );
  XNOR2_X1 U882 ( .A(n792), .B(KEYINPUT38), .ZN(n799) );
  NAND2_X1 U883 ( .A1(G117), .A2(n898), .ZN(n794) );
  NAND2_X1 U884 ( .A1(G141), .A2(n905), .ZN(n793) );
  NAND2_X1 U885 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U886 ( .A1(n897), .A2(G129), .ZN(n795) );
  XOR2_X1 U887 ( .A(KEYINPUT90), .B(n795), .Z(n796) );
  NOR2_X1 U888 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U889 ( .A1(n799), .A2(n798), .ZN(n893) );
  NAND2_X1 U890 ( .A1(G1996), .A2(n893), .ZN(n808) );
  NAND2_X1 U891 ( .A1(G95), .A2(n902), .ZN(n801) );
  NAND2_X1 U892 ( .A1(G131), .A2(n905), .ZN(n800) );
  NAND2_X1 U893 ( .A1(n801), .A2(n800), .ZN(n804) );
  NAND2_X1 U894 ( .A1(G119), .A2(n897), .ZN(n802) );
  XNOR2_X1 U895 ( .A(KEYINPUT89), .B(n802), .ZN(n803) );
  NOR2_X1 U896 ( .A1(n804), .A2(n803), .ZN(n806) );
  NAND2_X1 U897 ( .A1(n898), .A2(G107), .ZN(n805) );
  NAND2_X1 U898 ( .A1(n806), .A2(n805), .ZN(n887) );
  NAND2_X1 U899 ( .A1(G1991), .A2(n887), .ZN(n807) );
  NAND2_X1 U900 ( .A1(n808), .A2(n807), .ZN(n949) );
  NOR2_X1 U901 ( .A1(n810), .A2(n809), .ZN(n838) );
  XOR2_X1 U902 ( .A(n838), .B(KEYINPUT91), .Z(n811) );
  NAND2_X1 U903 ( .A1(n949), .A2(n811), .ZN(n812) );
  XOR2_X1 U904 ( .A(KEYINPUT92), .B(n812), .Z(n830) );
  INV_X1 U905 ( .A(n830), .ZN(n822) );
  NAND2_X1 U906 ( .A1(G104), .A2(n902), .ZN(n814) );
  NAND2_X1 U907 ( .A1(G140), .A2(n905), .ZN(n813) );
  NAND2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U909 ( .A(KEYINPUT34), .B(n815), .ZN(n820) );
  NAND2_X1 U910 ( .A1(G128), .A2(n897), .ZN(n817) );
  NAND2_X1 U911 ( .A1(G116), .A2(n898), .ZN(n816) );
  NAND2_X1 U912 ( .A1(n817), .A2(n816), .ZN(n818) );
  XOR2_X1 U913 ( .A(KEYINPUT35), .B(n818), .Z(n819) );
  NOR2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U915 ( .A(KEYINPUT36), .B(n821), .ZN(n909) );
  XNOR2_X1 U916 ( .A(KEYINPUT37), .B(G2067), .ZN(n836) );
  NOR2_X1 U917 ( .A1(n909), .A2(n836), .ZN(n946) );
  NAND2_X1 U918 ( .A1(n838), .A2(n946), .ZN(n833) );
  XNOR2_X1 U919 ( .A(G1986), .B(G290), .ZN(n979) );
  NAND2_X1 U920 ( .A1(n979), .A2(n838), .ZN(n823) );
  NAND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n841) );
  NOR2_X1 U922 ( .A1(G1996), .A2(n893), .ZN(n961) );
  NOR2_X1 U923 ( .A1(G1986), .A2(G290), .ZN(n828) );
  NOR2_X1 U924 ( .A1(n887), .A2(G1991), .ZN(n827) );
  XNOR2_X1 U925 ( .A(n827), .B(KEYINPUT104), .ZN(n953) );
  NOR2_X1 U926 ( .A1(n828), .A2(n953), .ZN(n829) );
  NOR2_X1 U927 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U928 ( .A1(n961), .A2(n831), .ZN(n832) );
  XNOR2_X1 U929 ( .A(n832), .B(KEYINPUT39), .ZN(n834) );
  NAND2_X1 U930 ( .A1(n834), .A2(n833), .ZN(n835) );
  XOR2_X1 U931 ( .A(KEYINPUT105), .B(n835), .Z(n837) );
  NAND2_X1 U932 ( .A1(n909), .A2(n836), .ZN(n945) );
  NAND2_X1 U933 ( .A1(n837), .A2(n945), .ZN(n839) );
  NAND2_X1 U934 ( .A1(n839), .A2(n838), .ZN(n840) );
  NAND2_X1 U935 ( .A1(n841), .A2(n840), .ZN(n843) );
  XNOR2_X1 U936 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n842) );
  XNOR2_X1 U937 ( .A(n843), .B(n842), .ZN(G329) );
  NAND2_X1 U938 ( .A1(G2106), .A2(n844), .ZN(G217) );
  AND2_X1 U939 ( .A1(G15), .A2(G2), .ZN(n845) );
  NAND2_X1 U940 ( .A1(G661), .A2(n845), .ZN(G259) );
  NAND2_X1 U941 ( .A1(G3), .A2(G1), .ZN(n846) );
  NAND2_X1 U942 ( .A1(n847), .A2(n846), .ZN(G188) );
  INV_X1 U944 ( .A(G96), .ZN(G221) );
  NOR2_X1 U945 ( .A1(n849), .A2(n848), .ZN(G325) );
  INV_X1 U946 ( .A(G325), .ZN(G261) );
  INV_X1 U947 ( .A(n850), .ZN(G319) );
  XOR2_X1 U948 ( .A(KEYINPUT112), .B(G1991), .Z(n852) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1986), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U951 ( .A(n853), .B(KEYINPUT41), .Z(n855) );
  XNOR2_X1 U952 ( .A(G1981), .B(G1966), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U954 ( .A(G1956), .B(G1961), .Z(n857) );
  XNOR2_X1 U955 ( .A(G1976), .B(G1971), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U957 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U958 ( .A(KEYINPUT111), .B(G2474), .ZN(n860) );
  XNOR2_X1 U959 ( .A(n861), .B(n860), .ZN(G229) );
  XOR2_X1 U960 ( .A(G2096), .B(KEYINPUT43), .Z(n863) );
  XNOR2_X1 U961 ( .A(G2072), .B(G2678), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U963 ( .A(n864), .B(KEYINPUT110), .Z(n866) );
  XNOR2_X1 U964 ( .A(G2067), .B(G2090), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U966 ( .A(KEYINPUT42), .B(G2100), .Z(n868) );
  XNOR2_X1 U967 ( .A(G2078), .B(G2084), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U969 ( .A(n870), .B(n869), .ZN(G227) );
  NAND2_X1 U970 ( .A1(G100), .A2(n902), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G112), .A2(n898), .ZN(n871) );
  NAND2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U973 ( .A(n873), .B(KEYINPUT113), .ZN(n875) );
  NAND2_X1 U974 ( .A1(G136), .A2(n905), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n878) );
  NAND2_X1 U976 ( .A1(n897), .A2(G124), .ZN(n876) );
  XOR2_X1 U977 ( .A(KEYINPUT44), .B(n876), .Z(n877) );
  NOR2_X1 U978 ( .A1(n878), .A2(n877), .ZN(G162) );
  NAND2_X1 U979 ( .A1(G130), .A2(n897), .ZN(n880) );
  NAND2_X1 U980 ( .A1(G118), .A2(n898), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U982 ( .A(KEYINPUT114), .B(n881), .ZN(n886) );
  NAND2_X1 U983 ( .A1(G106), .A2(n902), .ZN(n883) );
  NAND2_X1 U984 ( .A1(G142), .A2(n905), .ZN(n882) );
  NAND2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U986 ( .A(n884), .B(KEYINPUT45), .Z(n885) );
  NOR2_X1 U987 ( .A1(n886), .A2(n885), .ZN(n888) );
  XNOR2_X1 U988 ( .A(n888), .B(n887), .ZN(n892) );
  XOR2_X1 U989 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n890) );
  XNOR2_X1 U990 ( .A(G160), .B(G164), .ZN(n889) );
  XNOR2_X1 U991 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U992 ( .A(n892), .B(n891), .ZN(n895) );
  XNOR2_X1 U993 ( .A(n893), .B(G162), .ZN(n894) );
  XNOR2_X1 U994 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n951), .B(n896), .ZN(n911) );
  NAND2_X1 U996 ( .A1(G127), .A2(n897), .ZN(n900) );
  NAND2_X1 U997 ( .A1(G115), .A2(n898), .ZN(n899) );
  NAND2_X1 U998 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n901), .B(KEYINPUT47), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(G103), .A2(n902), .ZN(n903) );
  NAND2_X1 U1001 ( .A1(n904), .A2(n903), .ZN(n908) );
  NAND2_X1 U1002 ( .A1(G139), .A2(n905), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(KEYINPUT115), .B(n906), .ZN(n907) );
  NOR2_X1 U1004 ( .A1(n908), .A2(n907), .ZN(n956) );
  XNOR2_X1 U1005 ( .A(n909), .B(n956), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n912), .ZN(G395) );
  XOR2_X1 U1008 ( .A(n913), .B(G286), .Z(n915) );
  XNOR2_X1 U1009 ( .A(G171), .B(n970), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(n915), .B(n914), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(n916), .B(n973), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n917), .ZN(G397) );
  NOR2_X1 U1013 ( .A1(G229), .A2(G227), .ZN(n918) );
  XOR2_X1 U1014 ( .A(KEYINPUT49), .B(n918), .Z(n919) );
  NAND2_X1 U1015 ( .A1(G319), .A2(n919), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(G401), .A2(n920), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(KEYINPUT116), .B(n921), .ZN(n923) );
  NOR2_X1 U1018 ( .A1(G395), .A2(G397), .ZN(n922) );
  NAND2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  INV_X1 U1021 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1022 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n944) );
  XNOR2_X1 U1023 ( .A(G2090), .B(G35), .ZN(n936) );
  XNOR2_X1 U1024 ( .A(G2067), .B(G26), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(G33), .B(G2072), .ZN(n924) );
  NOR2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n930) );
  XOR2_X1 U1027 ( .A(G1991), .B(G25), .Z(n926) );
  NAND2_X1 U1028 ( .A1(n926), .A2(G28), .ZN(n928) );
  XNOR2_X1 U1029 ( .A(G32), .B(G1996), .ZN(n927) );
  NOR2_X1 U1030 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n933) );
  XOR2_X1 U1032 ( .A(G27), .B(n931), .Z(n932) );
  NOR2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1034 ( .A(KEYINPUT53), .B(n934), .ZN(n935) );
  NOR2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1036 ( .A(n937), .B(KEYINPUT118), .ZN(n940) );
  XOR2_X1 U1037 ( .A(G2084), .B(G34), .Z(n938) );
  XNOR2_X1 U1038 ( .A(KEYINPUT54), .B(n938), .ZN(n939) );
  NAND2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n942) );
  INV_X1 U1040 ( .A(G29), .ZN(n941) );
  NAND2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1042 ( .A(n944), .B(n943), .ZN(n969) );
  INV_X1 U1043 ( .A(n945), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n955) );
  XOR2_X1 U1045 ( .A(G160), .B(G2084), .Z(n948) );
  NOR2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n966) );
  XOR2_X1 U1050 ( .A(G2072), .B(n956), .Z(n958) );
  XOR2_X1 U1051 ( .A(G164), .B(G2078), .Z(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(KEYINPUT50), .B(n959), .ZN(n964) );
  XOR2_X1 U1054 ( .A(G2090), .B(G162), .Z(n960) );
  NOR2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1056 ( .A(KEYINPUT51), .B(n962), .Z(n963) );
  NAND2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1059 ( .A(n967), .B(KEYINPUT52), .Z(n968) );
  NAND2_X1 U1060 ( .A1(n969), .A2(n512), .ZN(n1026) );
  XNOR2_X1 U1061 ( .A(G16), .B(KEYINPUT56), .ZN(n995) );
  XOR2_X1 U1062 ( .A(G1348), .B(n970), .Z(n972) );
  XNOR2_X1 U1063 ( .A(G171), .B(G1961), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n988) );
  XOR2_X1 U1065 ( .A(n973), .B(G1341), .Z(n986) );
  XNOR2_X1 U1066 ( .A(G1971), .B(G166), .ZN(n981) );
  INV_X1 U1067 ( .A(n974), .ZN(n975) );
  NAND2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1069 ( .A(KEYINPUT119), .B(n977), .Z(n978) );
  NOR2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(G1956), .B(G299), .ZN(n982) );
  NOR2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1074 ( .A(KEYINPUT120), .B(n984), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1076 ( .A1(n988), .A2(n987), .ZN(n993) );
  XNOR2_X1 U1077 ( .A(G1966), .B(G168), .ZN(n990) );
  NAND2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1079 ( .A(n991), .B(KEYINPUT57), .ZN(n992) );
  NAND2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1081 ( .A1(n995), .A2(n994), .ZN(n1023) );
  XNOR2_X1 U1082 ( .A(G1986), .B(G24), .ZN(n1000) );
  XNOR2_X1 U1083 ( .A(G1976), .B(G23), .ZN(n997) );
  XNOR2_X1 U1084 ( .A(G22), .B(G1971), .ZN(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(KEYINPUT123), .B(n998), .ZN(n999) );
  NOR2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(KEYINPUT124), .B(n1001), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(n1002), .B(KEYINPUT58), .ZN(n1016) );
  XNOR2_X1 U1090 ( .A(G1981), .B(G6), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G1341), .B(G19), .ZN(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(KEYINPUT122), .B(n1005), .ZN(n1008) );
  XNOR2_X1 U1094 ( .A(n1006), .B(G20), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XOR2_X1 U1096 ( .A(KEYINPUT59), .B(G1348), .Z(n1009) );
  XNOR2_X1 U1097 ( .A(G4), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1099 ( .A(KEYINPUT60), .B(n1012), .Z(n1014) );
  XNOR2_X1 U1100 ( .A(G1961), .B(G5), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XNOR2_X1 U1103 ( .A(G21), .B(G1966), .ZN(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(n1019), .B(KEYINPUT61), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(G16), .B(KEYINPUT121), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1109 ( .A(KEYINPUT125), .B(n1024), .Z(n1025) );
  NOR2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1111 ( .A1(n1027), .A2(G11), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(n1028), .B(KEYINPUT126), .ZN(n1029) );
  XNOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1029), .ZN(G150) );
  INV_X1 U1114 ( .A(G150), .ZN(G311) );
endmodule

