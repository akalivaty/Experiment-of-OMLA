

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732;

  AND2_X1 U360 ( .A1(n411), .A2(n410), .ZN(n409) );
  NOR2_X1 U361 ( .A1(n545), .A2(n544), .ZN(n620) );
  XNOR2_X2 U362 ( .A(G101), .B(KEYINPUT75), .ZN(n424) );
  XNOR2_X2 U363 ( .A(n406), .B(KEYINPUT69), .ZN(n388) );
  XNOR2_X2 U364 ( .A(n380), .B(n369), .ZN(n712) );
  XNOR2_X2 U365 ( .A(n379), .B(n342), .ZN(n369) );
  XNOR2_X1 U366 ( .A(n551), .B(n462), .ZN(n586) );
  INV_X1 U367 ( .A(n551), .ZN(n687) );
  XNOR2_X2 U368 ( .A(n499), .B(G478), .ZN(n536) );
  XNOR2_X2 U369 ( .A(n719), .B(G146), .ZN(n449) );
  NOR2_X1 U370 ( .A1(n732), .A2(n731), .ZN(n405) );
  NOR2_X1 U371 ( .A1(n527), .A2(n356), .ZN(n397) );
  NOR2_X1 U372 ( .A1(n672), .A2(n671), .ZN(n569) );
  XNOR2_X1 U373 ( .A(n448), .B(KEYINPUT74), .ZN(n527) );
  NAND2_X1 U374 ( .A1(n706), .A2(n720), .ZN(n367) );
  AND2_X1 U375 ( .A1(n340), .A2(n348), .ZN(n347) );
  XNOR2_X1 U376 ( .A(n405), .B(KEYINPUT46), .ZN(n404) );
  XNOR2_X1 U377 ( .A(n563), .B(n562), .ZN(n732) );
  XNOR2_X1 U378 ( .A(n418), .B(n344), .ZN(n663) );
  AND2_X1 U379 ( .A1(n396), .A2(n392), .ZN(n391) );
  XNOR2_X1 U380 ( .A(n397), .B(KEYINPUT33), .ZN(n699) );
  INV_X1 U381 ( .A(n586), .ZN(n356) );
  XNOR2_X1 U382 ( .A(n362), .B(n337), .ZN(n534) );
  XNOR2_X1 U383 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U384 ( .A(n401), .B(G146), .ZN(n467) );
  XNOR2_X1 U385 ( .A(n423), .B(G137), .ZN(n421) );
  XNOR2_X1 U386 ( .A(KEYINPUT4), .B(G131), .ZN(n423) );
  XNOR2_X1 U387 ( .A(G107), .B(G104), .ZN(n425) );
  XNOR2_X2 U388 ( .A(n561), .B(KEYINPUT39), .ZN(n599) );
  NOR2_X1 U389 ( .A1(G237), .A2(G953), .ZN(n454) );
  XNOR2_X1 U390 ( .A(n467), .B(n430), .ZN(n501) );
  INV_X1 U391 ( .A(KEYINPUT10), .ZN(n430) );
  XNOR2_X1 U392 ( .A(n425), .B(n424), .ZN(n379) );
  NOR2_X1 U393 ( .A1(n620), .A2(n547), .ZN(n414) );
  XOR2_X1 U394 ( .A(KEYINPUT68), .B(G140), .Z(n431) );
  NAND2_X1 U395 ( .A1(n360), .A2(n403), .ZN(n359) );
  INV_X1 U396 ( .A(G237), .ZN(n472) );
  NOR2_X1 U397 ( .A1(n557), .A2(n564), .ZN(n558) );
  NAND2_X1 U398 ( .A1(n638), .A2(n473), .ZN(n428) );
  OR2_X1 U399 ( .A1(n631), .A2(G902), .ZN(n362) );
  XNOR2_X1 U400 ( .A(n402), .B(n444), .ZN(n679) );
  XNOR2_X1 U401 ( .A(n383), .B(n459), .ZN(n608) );
  XNOR2_X1 U402 ( .A(G110), .B(G119), .ZN(n435) );
  XNOR2_X1 U403 ( .A(n501), .B(n431), .ZN(n718) );
  XNOR2_X1 U404 ( .A(n489), .B(n488), .ZN(n490) );
  INV_X1 U405 ( .A(KEYINPUT9), .ZN(n488) );
  XNOR2_X1 U406 ( .A(G107), .B(G122), .ZN(n489) );
  XNOR2_X1 U407 ( .A(n365), .B(n363), .ZN(n506) );
  XNOR2_X1 U408 ( .A(n502), .B(n366), .ZN(n365) );
  XNOR2_X1 U409 ( .A(n503), .B(n364), .ZN(n363) );
  XNOR2_X1 U410 ( .A(KEYINPUT11), .B(KEYINPUT95), .ZN(n366) );
  INV_X1 U411 ( .A(KEYINPUT89), .ZN(n420) );
  INV_X1 U412 ( .A(n431), .ZN(n407) );
  XNOR2_X1 U413 ( .A(n465), .B(n466), .ZN(n378) );
  XNOR2_X1 U414 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n466) );
  INV_X1 U415 ( .A(G125), .ZN(n401) );
  XNOR2_X1 U416 ( .A(KEYINPUT79), .B(KEYINPUT4), .ZN(n469) );
  XNOR2_X1 U417 ( .A(n464), .B(n463), .ZN(n380) );
  XNOR2_X1 U418 ( .A(KEYINPUT16), .B(G122), .ZN(n463) );
  INV_X1 U419 ( .A(G953), .ZN(n721) );
  AND2_X1 U420 ( .A1(n393), .A2(n682), .ZN(n392) );
  NAND2_X1 U421 ( .A1(n395), .A2(n394), .ZN(n393) );
  INV_X1 U422 ( .A(n588), .ZN(n394) );
  NAND2_X1 U423 ( .A1(n477), .A2(KEYINPUT85), .ZN(n410) );
  XNOR2_X1 U424 ( .A(G131), .B(G113), .ZN(n364) );
  XNOR2_X1 U425 ( .A(G140), .B(G143), .ZN(n503) );
  XNOR2_X1 U426 ( .A(G104), .B(G122), .ZN(n502) );
  INV_X1 U427 ( .A(KEYINPUT104), .ZN(n415) );
  NAND2_X1 U428 ( .A1(n351), .A2(n412), .ZN(n350) );
  AND2_X2 U429 ( .A1(n361), .A2(n384), .ZN(n720) );
  AND2_X1 U430 ( .A1(n385), .A2(n601), .ZN(n384) );
  NAND2_X1 U431 ( .A1(n359), .A2(n358), .ZN(n361) );
  INV_X1 U432 ( .A(n590), .ZN(n597) );
  NOR2_X1 U433 ( .A1(n699), .A2(n528), .ZN(n485) );
  OR2_X1 U434 ( .A1(n586), .A2(n355), .ZN(n521) );
  INV_X1 U435 ( .A(n372), .ZN(n355) );
  INV_X1 U436 ( .A(n688), .ZN(n419) );
  NOR2_X1 U437 ( .A1(n560), .A2(n559), .ZN(n593) );
  XNOR2_X1 U438 ( .A(n534), .B(n535), .ZN(n537) );
  XOR2_X1 U439 ( .A(KEYINPUT72), .B(KEYINPUT22), .Z(n515) );
  XOR2_X1 U440 ( .A(n609), .B(KEYINPUT62), .Z(n610) );
  XNOR2_X1 U441 ( .A(n718), .B(n434), .ZN(n371) );
  XNOR2_X1 U442 ( .A(n491), .B(n490), .ZN(n498) );
  XNOR2_X1 U443 ( .A(n507), .B(n508), .ZN(n631) );
  XNOR2_X1 U444 ( .A(KEYINPUT12), .B(KEYINPUT96), .ZN(n500) );
  XNOR2_X1 U445 ( .A(n449), .B(n398), .ZN(n638) );
  XNOR2_X1 U446 ( .A(n407), .B(n400), .ZN(n399) );
  XNOR2_X1 U447 ( .A(n426), .B(n420), .ZN(n400) );
  XNOR2_X1 U448 ( .A(n470), .B(n377), .ZN(n376) );
  XNOR2_X1 U449 ( .A(n467), .B(n378), .ZN(n377) );
  NOR2_X1 U450 ( .A1(n373), .A2(G952), .ZN(n647) );
  BUF_X1 U451 ( .A(n721), .Z(n373) );
  XNOR2_X1 U452 ( .A(n589), .B(KEYINPUT110), .ZN(n357) );
  NAND2_X1 U453 ( .A1(n391), .A2(n389), .ZN(n589) );
  NAND2_X1 U454 ( .A1(n390), .A2(n394), .ZN(n389) );
  AND2_X1 U455 ( .A1(n583), .A2(n582), .ZN(n336) );
  XOR2_X1 U456 ( .A(n509), .B(G475), .Z(n337) );
  XOR2_X1 U457 ( .A(n475), .B(n474), .Z(n338) );
  OR2_X1 U458 ( .A1(n477), .A2(KEYINPUT85), .ZN(n339) );
  XOR2_X1 U459 ( .A(n540), .B(n415), .Z(n340) );
  AND2_X1 U460 ( .A1(n357), .A2(n657), .ZN(n341) );
  XOR2_X1 U461 ( .A(KEYINPUT86), .B(G110), .Z(n342) );
  AND2_X1 U462 ( .A1(n381), .A2(n588), .ZN(n343) );
  XOR2_X1 U463 ( .A(n529), .B(KEYINPUT93), .Z(n344) );
  XNOR2_X1 U464 ( .A(KEYINPUT66), .B(KEYINPUT0), .ZN(n345) );
  XNOR2_X1 U465 ( .A(n371), .B(n441), .ZN(n605) );
  XNOR2_X1 U466 ( .A(G119), .B(KEYINPUT126), .ZN(n346) );
  NAND2_X2 U467 ( .A1(n349), .A2(n347), .ZN(n368) );
  NAND2_X1 U468 ( .A1(n625), .A2(n549), .ZN(n348) );
  AND2_X2 U469 ( .A1(n352), .A2(n350), .ZN(n349) );
  NAND2_X1 U470 ( .A1(n414), .A2(n375), .ZN(n351) );
  NAND2_X1 U471 ( .A1(n354), .A2(n353), .ZN(n352) );
  NAND2_X1 U472 ( .A1(n526), .A2(KEYINPUT84), .ZN(n353) );
  INV_X1 U473 ( .A(n625), .ZN(n354) );
  XNOR2_X1 U474 ( .A(n357), .B(G125), .ZN(n729) );
  NAND2_X1 U475 ( .A1(n388), .A2(n387), .ZN(n358) );
  INV_X1 U476 ( .A(n388), .ZN(n360) );
  XNOR2_X2 U477 ( .A(n367), .B(KEYINPUT2), .ZN(n667) );
  XNOR2_X2 U478 ( .A(n368), .B(n550), .ZN(n706) );
  XNOR2_X1 U479 ( .A(n399), .B(n369), .ZN(n398) );
  XNOR2_X2 U480 ( .A(n370), .B(n345), .ZN(n531) );
  NOR2_X2 U481 ( .A1(n573), .A2(n484), .ZN(n370) );
  XNOR2_X2 U482 ( .A(n381), .B(KEYINPUT19), .ZN(n573) );
  NAND2_X2 U483 ( .A1(n409), .A2(n408), .ZN(n381) );
  XNOR2_X1 U484 ( .A(n712), .B(n376), .ZN(n644) );
  NAND2_X1 U485 ( .A1(n681), .A2(n530), .ZN(n557) );
  OR2_X2 U486 ( .A1(n644), .A2(n471), .ZN(n417) );
  NAND2_X1 U487 ( .A1(n541), .A2(n523), .ZN(n524) );
  XNOR2_X2 U488 ( .A(n516), .B(n515), .ZN(n541) );
  BUF_X2 U489 ( .A(n679), .Z(n372) );
  NOR2_X2 U490 ( .A1(n679), .A2(n678), .ZN(n681) );
  XNOR2_X1 U491 ( .A(n374), .B(n605), .ZN(n422) );
  NAND2_X1 U492 ( .A1(n642), .A2(G217), .ZN(n374) );
  NAND2_X1 U493 ( .A1(n525), .A2(n375), .ZN(n526) );
  XNOR2_X1 U494 ( .A(n375), .B(n346), .ZN(G21) );
  XNOR2_X2 U495 ( .A(n524), .B(KEYINPUT32), .ZN(n375) );
  XNOR2_X2 U496 ( .A(n457), .B(n456), .ZN(n464) );
  INV_X1 U497 ( .A(n381), .ZN(n395) );
  XNOR2_X2 U498 ( .A(n382), .B(n461), .ZN(n551) );
  NAND2_X1 U499 ( .A1(n608), .A2(n473), .ZN(n382) );
  NAND2_X1 U500 ( .A1(n452), .A2(n453), .ZN(n383) );
  NAND2_X1 U501 ( .A1(n386), .A2(KEYINPUT48), .ZN(n385) );
  INV_X1 U502 ( .A(n404), .ZN(n386) );
  NAND2_X1 U503 ( .A1(n404), .A2(n403), .ZN(n387) );
  INV_X1 U504 ( .A(n594), .ZN(n390) );
  NAND2_X1 U505 ( .A1(n594), .A2(n343), .ZN(n396) );
  XNOR2_X2 U506 ( .A(n587), .B(KEYINPUT107), .ZN(n594) );
  NAND2_X1 U507 ( .A1(n605), .A2(n473), .ZN(n402) );
  INV_X1 U508 ( .A(KEYINPUT48), .ZN(n403) );
  NAND2_X1 U509 ( .A1(n341), .A2(n336), .ZN(n406) );
  NOR2_X2 U510 ( .A1(n634), .A2(n647), .ZN(n635) );
  NOR2_X2 U511 ( .A1(n648), .A2(n647), .ZN(n649) );
  OR2_X1 U512 ( .A1(n590), .A2(n339), .ZN(n408) );
  XNOR2_X2 U513 ( .A(n417), .B(n338), .ZN(n590) );
  NAND2_X1 U514 ( .A1(n590), .A2(KEYINPUT85), .ZN(n411) );
  XNOR2_X2 U515 ( .A(G116), .B(G113), .ZN(n457) );
  NAND2_X1 U516 ( .A1(n416), .A2(n413), .ZN(n412) );
  INV_X1 U517 ( .A(n548), .ZN(n413) );
  INV_X1 U518 ( .A(n620), .ZN(n416) );
  INV_X1 U519 ( .A(n531), .ZN(n528) );
  NAND2_X1 U520 ( .A1(n531), .A2(n419), .ZN(n418) );
  XNOR2_X2 U521 ( .A(n486), .B(n421), .ZN(n719) );
  NOR2_X2 U522 ( .A1(n612), .A2(n647), .ZN(n614) );
  XNOR2_X2 U523 ( .A(KEYINPUT3), .B(G119), .ZN(n456) );
  XNOR2_X1 U524 ( .A(n501), .B(n500), .ZN(n508) );
  XNOR2_X1 U525 ( .A(KEYINPUT109), .B(KEYINPUT36), .ZN(n588) );
  NAND2_X1 U526 ( .A1(n593), .A2(n669), .ZN(n561) );
  INV_X1 U527 ( .A(n647), .ZN(n606) );
  INV_X1 U528 ( .A(KEYINPUT63), .ZN(n613) );
  NAND2_X1 U529 ( .A1(n422), .A2(n606), .ZN(n607) );
  XNOR2_X1 U530 ( .A(n607), .B(KEYINPUT121), .ZN(G66) );
  XNOR2_X2 U531 ( .A(G143), .B(G128), .ZN(n468) );
  XNOR2_X2 U532 ( .A(n468), .B(G134), .ZN(n486) );
  NAND2_X1 U533 ( .A1(G227), .A2(n721), .ZN(n426) );
  INV_X1 U534 ( .A(G902), .ZN(n473) );
  XOR2_X1 U535 ( .A(KEYINPUT70), .B(G469), .Z(n427) );
  XNOR2_X2 U536 ( .A(n428), .B(n427), .ZN(n567) );
  XNOR2_X1 U537 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n429) );
  XNOR2_X1 U538 ( .A(n567), .B(n429), .ZN(n517) );
  XOR2_X1 U539 ( .A(KEYINPUT90), .B(KEYINPUT24), .Z(n433) );
  XNOR2_X1 U540 ( .A(KEYINPUT78), .B(KEYINPUT23), .ZN(n432) );
  XNOR2_X1 U541 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U542 ( .A(G137), .B(G128), .Z(n436) );
  XNOR2_X1 U543 ( .A(n436), .B(n435), .ZN(n440) );
  NAND2_X1 U544 ( .A1(n721), .A2(G234), .ZN(n438) );
  XNOR2_X1 U545 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n437) );
  XNOR2_X1 U546 ( .A(n438), .B(n437), .ZN(n492) );
  NAND2_X1 U547 ( .A1(n492), .A2(G221), .ZN(n439) );
  XNOR2_X1 U548 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U549 ( .A(KEYINPUT15), .B(G902), .ZN(n602) );
  NAND2_X1 U550 ( .A1(G234), .A2(n602), .ZN(n442) );
  XNOR2_X1 U551 ( .A(KEYINPUT20), .B(n442), .ZN(n445) );
  NAND2_X1 U552 ( .A1(n445), .A2(G217), .ZN(n443) );
  XNOR2_X1 U553 ( .A(n443), .B(KEYINPUT25), .ZN(n444) );
  NAND2_X1 U554 ( .A1(n445), .A2(G221), .ZN(n447) );
  XOR2_X1 U555 ( .A(KEYINPUT21), .B(KEYINPUT91), .Z(n446) );
  XNOR2_X1 U556 ( .A(n447), .B(n446), .ZN(n678) );
  NAND2_X1 U557 ( .A1(n517), .A2(n681), .ZN(n448) );
  NAND2_X1 U558 ( .A1(KEYINPUT5), .A2(n449), .ZN(n453) );
  INV_X1 U559 ( .A(KEYINPUT5), .ZN(n451) );
  INV_X1 U560 ( .A(n449), .ZN(n450) );
  NAND2_X1 U561 ( .A1(n451), .A2(n450), .ZN(n452) );
  XNOR2_X1 U562 ( .A(n454), .B(KEYINPUT76), .ZN(n504) );
  NAND2_X1 U563 ( .A1(n504), .A2(G210), .ZN(n455) );
  XNOR2_X1 U564 ( .A(n455), .B(G101), .ZN(n458) );
  XOR2_X1 U565 ( .A(n464), .B(n458), .Z(n459) );
  INV_X1 U566 ( .A(KEYINPUT71), .ZN(n460) );
  XNOR2_X1 U567 ( .A(n460), .B(G472), .ZN(n461) );
  INV_X1 U568 ( .A(KEYINPUT6), .ZN(n462) );
  NAND2_X1 U569 ( .A1(n721), .A2(G224), .ZN(n465) );
  XNOR2_X1 U570 ( .A(n468), .B(n469), .ZN(n470) );
  INV_X1 U571 ( .A(n602), .ZN(n471) );
  NAND2_X1 U572 ( .A1(n473), .A2(n472), .ZN(n476) );
  NAND2_X1 U573 ( .A1(n476), .A2(G210), .ZN(n475) );
  INV_X1 U574 ( .A(KEYINPUT82), .ZN(n474) );
  NAND2_X1 U575 ( .A1(n476), .A2(G214), .ZN(n668) );
  INV_X1 U576 ( .A(n668), .ZN(n477) );
  XOR2_X1 U577 ( .A(KEYINPUT14), .B(KEYINPUT87), .Z(n479) );
  NAND2_X1 U578 ( .A1(G237), .A2(G234), .ZN(n478) );
  XNOR2_X1 U579 ( .A(n479), .B(n478), .ZN(n482) );
  AND2_X1 U580 ( .A1(G953), .A2(G902), .ZN(n480) );
  NAND2_X1 U581 ( .A1(n482), .A2(n480), .ZN(n553) );
  NOR2_X1 U582 ( .A1(G898), .A2(n553), .ZN(n481) );
  XNOR2_X1 U583 ( .A(n481), .B(KEYINPUT88), .ZN(n483) );
  NAND2_X1 U584 ( .A1(G952), .A2(n482), .ZN(n697) );
  NOR2_X1 U585 ( .A1(n697), .A2(G953), .ZN(n556) );
  NOR2_X1 U586 ( .A1(n483), .A2(n556), .ZN(n484) );
  XNOR2_X1 U587 ( .A(n485), .B(KEYINPUT34), .ZN(n512) );
  XNOR2_X1 U588 ( .A(n486), .B(KEYINPUT101), .ZN(n487) );
  XNOR2_X1 U589 ( .A(n487), .B(KEYINPUT7), .ZN(n491) );
  NAND2_X1 U590 ( .A1(n492), .A2(G217), .ZN(n496) );
  XOR2_X1 U591 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n494) );
  XNOR2_X1 U592 ( .A(G116), .B(KEYINPUT102), .ZN(n493) );
  XNOR2_X1 U593 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U594 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U595 ( .A(n498), .B(n497), .ZN(n627) );
  NOR2_X1 U596 ( .A1(n627), .A2(G902), .ZN(n499) );
  NAND2_X1 U597 ( .A1(n504), .A2(G214), .ZN(n505) );
  XNOR2_X1 U598 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U599 ( .A(KEYINPUT97), .B(KEYINPUT13), .ZN(n509) );
  NOR2_X1 U600 ( .A1(n536), .A2(n534), .ZN(n510) );
  XNOR2_X1 U601 ( .A(n510), .B(KEYINPUT105), .ZN(n591) );
  INV_X1 U602 ( .A(n591), .ZN(n511) );
  NAND2_X1 U603 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X2 U604 ( .A(n513), .B(KEYINPUT35), .ZN(n625) );
  NAND2_X1 U605 ( .A1(n536), .A2(n534), .ZN(n671) );
  NOR2_X1 U606 ( .A1(n671), .A2(n678), .ZN(n514) );
  NAND2_X1 U607 ( .A1(n531), .A2(n514), .ZN(n516) );
  INV_X1 U608 ( .A(n517), .ZN(n543) );
  INV_X1 U609 ( .A(n543), .ZN(n682) );
  NAND2_X1 U610 ( .A1(n687), .A2(n372), .ZN(n518) );
  NOR2_X1 U611 ( .A1(n682), .A2(n518), .ZN(n519) );
  NAND2_X1 U612 ( .A1(n541), .A2(n519), .ZN(n615) );
  INV_X1 U613 ( .A(n615), .ZN(n520) );
  NOR2_X1 U614 ( .A1(n520), .A2(KEYINPUT44), .ZN(n525) );
  NOR2_X1 U615 ( .A1(n543), .A2(n521), .ZN(n522) );
  XNOR2_X1 U616 ( .A(n522), .B(KEYINPUT80), .ZN(n523) );
  OR2_X1 U617 ( .A1(n527), .A2(n687), .ZN(n688) );
  XOR2_X1 U618 ( .A(KEYINPUT94), .B(KEYINPUT31), .Z(n529) );
  INV_X1 U619 ( .A(n567), .ZN(n530) );
  NOR2_X1 U620 ( .A1(n557), .A2(n551), .ZN(n532) );
  NAND2_X1 U621 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U622 ( .A(n533), .B(KEYINPUT92), .ZN(n616) );
  NAND2_X1 U623 ( .A1(n663), .A2(n616), .ZN(n539) );
  INV_X1 U624 ( .A(KEYINPUT98), .ZN(n535) );
  NOR2_X1 U625 ( .A1(n537), .A2(n536), .ZN(n654) );
  NAND2_X1 U626 ( .A1(n537), .A2(n536), .ZN(n662) );
  INV_X1 U627 ( .A(n662), .ZN(n617) );
  NOR2_X1 U628 ( .A1(n654), .A2(n617), .ZN(n538) );
  XNOR2_X1 U629 ( .A(n538), .B(KEYINPUT103), .ZN(n579) );
  NAND2_X1 U630 ( .A1(n539), .A2(n579), .ZN(n540) );
  INV_X1 U631 ( .A(n541), .ZN(n545) );
  NOR2_X1 U632 ( .A1(n586), .A2(n372), .ZN(n542) );
  NAND2_X1 U633 ( .A1(n543), .A2(n542), .ZN(n544) );
  INV_X1 U634 ( .A(KEYINPUT44), .ZN(n546) );
  NAND2_X1 U635 ( .A1(n546), .A2(KEYINPUT84), .ZN(n548) );
  NAND2_X1 U636 ( .A1(n615), .A2(KEYINPUT44), .ZN(n547) );
  AND2_X1 U637 ( .A1(KEYINPUT84), .A2(n548), .ZN(n549) );
  XOR2_X1 U638 ( .A(KEYINPUT83), .B(KEYINPUT45), .Z(n550) );
  NAND2_X1 U639 ( .A1(n551), .A2(n668), .ZN(n552) );
  XNOR2_X1 U640 ( .A(KEYINPUT30), .B(n552), .ZN(n560) );
  XNOR2_X1 U641 ( .A(KEYINPUT106), .B(n553), .ZN(n554) );
  NOR2_X1 U642 ( .A1(G900), .A2(n554), .ZN(n555) );
  NOR2_X1 U643 ( .A1(n556), .A2(n555), .ZN(n564) );
  XNOR2_X1 U644 ( .A(n558), .B(KEYINPUT77), .ZN(n559) );
  XOR2_X1 U645 ( .A(KEYINPUT38), .B(n597), .Z(n669) );
  NAND2_X1 U646 ( .A1(n599), .A2(n617), .ZN(n563) );
  INV_X1 U647 ( .A(KEYINPUT40), .ZN(n562) );
  XOR2_X1 U648 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n572) );
  NOR2_X1 U649 ( .A1(n564), .A2(n678), .ZN(n565) );
  NAND2_X1 U650 ( .A1(n372), .A2(n565), .ZN(n584) );
  NOR2_X1 U651 ( .A1(n584), .A2(n687), .ZN(n566) );
  XOR2_X1 U652 ( .A(KEYINPUT28), .B(n566), .Z(n568) );
  NOR2_X1 U653 ( .A1(n568), .A2(n567), .ZN(n575) );
  NAND2_X1 U654 ( .A1(n669), .A2(n668), .ZN(n672) );
  XNOR2_X1 U655 ( .A(KEYINPUT41), .B(n569), .ZN(n698) );
  INV_X1 U656 ( .A(n698), .ZN(n570) );
  NAND2_X1 U657 ( .A1(n575), .A2(n570), .ZN(n571) );
  XNOR2_X1 U658 ( .A(n572), .B(n571), .ZN(n731) );
  INV_X1 U659 ( .A(n579), .ZN(n673) );
  NOR2_X1 U660 ( .A1(n673), .A2(KEYINPUT73), .ZN(n577) );
  INV_X1 U661 ( .A(n573), .ZN(n574) );
  NAND2_X1 U662 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X2 U663 ( .A(n576), .B(KEYINPUT81), .ZN(n659) );
  NAND2_X1 U664 ( .A1(n577), .A2(n659), .ZN(n578) );
  NAND2_X1 U665 ( .A1(n578), .A2(KEYINPUT47), .ZN(n583) );
  XNOR2_X1 U666 ( .A(KEYINPUT73), .B(n579), .ZN(n580) );
  NOR2_X1 U667 ( .A1(KEYINPUT47), .A2(n580), .ZN(n581) );
  NAND2_X1 U668 ( .A1(n581), .A2(n659), .ZN(n582) );
  NOR2_X1 U669 ( .A1(n584), .A2(n662), .ZN(n585) );
  NAND2_X1 U670 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U671 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U672 ( .A1(n593), .A2(n592), .ZN(n657) );
  NAND2_X1 U673 ( .A1(n594), .A2(n668), .ZN(n595) );
  NOR2_X1 U674 ( .A1(n682), .A2(n595), .ZN(n596) );
  XNOR2_X1 U675 ( .A(n596), .B(KEYINPUT43), .ZN(n598) );
  NOR2_X1 U676 ( .A1(n598), .A2(n597), .ZN(n621) );
  NAND2_X1 U677 ( .A1(n654), .A2(n599), .ZN(n666) );
  INV_X1 U678 ( .A(n666), .ZN(n600) );
  NOR2_X1 U679 ( .A1(n621), .A2(n600), .ZN(n601) );
  NAND2_X1 U680 ( .A1(n667), .A2(n471), .ZN(n604) );
  INV_X1 U681 ( .A(KEYINPUT64), .ZN(n603) );
  XNOR2_X2 U682 ( .A(n604), .B(n603), .ZN(n642) );
  NAND2_X1 U683 ( .A1(n642), .A2(G472), .ZN(n611) );
  BUF_X1 U684 ( .A(n608), .Z(n609) );
  XNOR2_X1 U685 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U686 ( .A(n614), .B(n613), .ZN(G57) );
  XNOR2_X1 U687 ( .A(n615), .B(G110), .ZN(G12) );
  INV_X1 U688 ( .A(n616), .ZN(n650) );
  NAND2_X1 U689 ( .A1(n650), .A2(n617), .ZN(n618) );
  XNOR2_X1 U690 ( .A(n618), .B(G104), .ZN(G6) );
  XNOR2_X1 U691 ( .A(G101), .B(KEYINPUT111), .ZN(n619) );
  XNOR2_X1 U692 ( .A(n620), .B(n619), .ZN(G3) );
  XOR2_X1 U693 ( .A(G140), .B(n621), .Z(G42) );
  XNOR2_X1 U694 ( .A(G116), .B(KEYINPUT115), .ZN(n624) );
  INV_X1 U695 ( .A(n663), .ZN(n622) );
  NAND2_X1 U696 ( .A1(n622), .A2(n654), .ZN(n623) );
  XOR2_X1 U697 ( .A(n624), .B(n623), .Z(G18) );
  XOR2_X1 U698 ( .A(n625), .B(G122), .Z(G24) );
  BUF_X1 U699 ( .A(n642), .Z(n626) );
  NAND2_X1 U700 ( .A1(n626), .A2(G478), .ZN(n628) );
  XNOR2_X1 U701 ( .A(n628), .B(n627), .ZN(n629) );
  NOR2_X1 U702 ( .A1(n629), .A2(n647), .ZN(G63) );
  NAND2_X1 U703 ( .A1(n642), .A2(G475), .ZN(n633) );
  XOR2_X1 U704 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n630) );
  XNOR2_X1 U705 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U706 ( .A(n635), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U707 ( .A1(n626), .A2(G469), .ZN(n640) );
  XOR2_X1 U708 ( .A(KEYINPUT119), .B(KEYINPUT57), .Z(n636) );
  XNOR2_X1 U709 ( .A(n636), .B(KEYINPUT58), .ZN(n637) );
  XNOR2_X1 U710 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U711 ( .A(n640), .B(n639), .ZN(n641) );
  NOR2_X1 U712 ( .A1(n641), .A2(n647), .ZN(G54) );
  NAND2_X1 U713 ( .A1(n642), .A2(G210), .ZN(n646) );
  XOR2_X1 U714 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n643) );
  XNOR2_X1 U715 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n646), .B(n645), .ZN(n648) );
  XNOR2_X1 U717 ( .A(n649), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U718 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n652) );
  NAND2_X1 U719 ( .A1(n650), .A2(n654), .ZN(n651) );
  XOR2_X1 U720 ( .A(n652), .B(n651), .Z(n653) );
  XNOR2_X1 U721 ( .A(G107), .B(n653), .ZN(G9) );
  XOR2_X1 U722 ( .A(G128), .B(KEYINPUT29), .Z(n656) );
  NAND2_X1 U723 ( .A1(n659), .A2(n654), .ZN(n655) );
  XNOR2_X1 U724 ( .A(n656), .B(n655), .ZN(G30) );
  XNOR2_X1 U725 ( .A(G143), .B(KEYINPUT112), .ZN(n658) );
  XNOR2_X1 U726 ( .A(n658), .B(n657), .ZN(G45) );
  XOR2_X1 U727 ( .A(G146), .B(KEYINPUT113), .Z(n661) );
  NAND2_X1 U728 ( .A1(n659), .A2(n617), .ZN(n660) );
  XNOR2_X1 U729 ( .A(n661), .B(n660), .ZN(G48) );
  NOR2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U731 ( .A(KEYINPUT114), .B(n664), .Z(n665) );
  XNOR2_X1 U732 ( .A(G113), .B(n665), .ZN(G15) );
  XNOR2_X1 U733 ( .A(G134), .B(n666), .ZN(G36) );
  BUF_X1 U734 ( .A(n667), .Z(n704) );
  NOR2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U736 ( .A1(n671), .A2(n670), .ZN(n675) );
  NOR2_X1 U737 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U738 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U739 ( .A(n676), .B(KEYINPUT118), .ZN(n677) );
  NOR2_X1 U740 ( .A1(n699), .A2(n677), .ZN(n694) );
  NAND2_X1 U741 ( .A1(n372), .A2(n678), .ZN(n680) );
  XNOR2_X1 U742 ( .A(n680), .B(KEYINPUT49), .ZN(n685) );
  NOR2_X1 U743 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U744 ( .A(n683), .B(KEYINPUT50), .ZN(n684) );
  NOR2_X1 U745 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U746 ( .A1(n687), .A2(n686), .ZN(n689) );
  NAND2_X1 U747 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U748 ( .A(n690), .B(KEYINPUT51), .ZN(n691) );
  XOR2_X1 U749 ( .A(KEYINPUT117), .B(n691), .Z(n692) );
  NOR2_X1 U750 ( .A1(n698), .A2(n692), .ZN(n693) );
  NOR2_X1 U751 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U752 ( .A(n695), .B(KEYINPUT52), .ZN(n696) );
  NOR2_X1 U753 ( .A1(n697), .A2(n696), .ZN(n701) );
  NOR2_X1 U754 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U755 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U756 ( .A1(n702), .A2(n373), .ZN(n703) );
  NOR2_X1 U757 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U758 ( .A(n705), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U759 ( .A1(n706), .A2(n373), .ZN(n707) );
  XNOR2_X1 U760 ( .A(n707), .B(KEYINPUT122), .ZN(n711) );
  NAND2_X1 U761 ( .A1(G953), .A2(G224), .ZN(n708) );
  XNOR2_X1 U762 ( .A(KEYINPUT61), .B(n708), .ZN(n709) );
  NAND2_X1 U763 ( .A1(n709), .A2(G898), .ZN(n710) );
  NAND2_X1 U764 ( .A1(n711), .A2(n710), .ZN(n717) );
  NOR2_X1 U765 ( .A1(G898), .A2(n373), .ZN(n713) );
  NOR2_X1 U766 ( .A1(n712), .A2(n713), .ZN(n715) );
  XOR2_X1 U767 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n714) );
  XNOR2_X1 U768 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U769 ( .A(n717), .B(n716), .ZN(G69) );
  XNOR2_X1 U770 ( .A(n719), .B(n718), .ZN(n723) );
  XOR2_X1 U771 ( .A(n723), .B(n720), .Z(n722) );
  NAND2_X1 U772 ( .A1(n722), .A2(n373), .ZN(n728) );
  XNOR2_X1 U773 ( .A(G227), .B(n723), .ZN(n724) );
  NAND2_X1 U774 ( .A1(n724), .A2(G900), .ZN(n725) );
  XOR2_X1 U775 ( .A(KEYINPUT125), .B(n725), .Z(n726) );
  NAND2_X1 U776 ( .A1(G953), .A2(n726), .ZN(n727) );
  NAND2_X1 U777 ( .A1(n728), .A2(n727), .ZN(G72) );
  XOR2_X1 U778 ( .A(KEYINPUT37), .B(KEYINPUT116), .Z(n730) );
  XNOR2_X1 U779 ( .A(n730), .B(n729), .ZN(G27) );
  XOR2_X1 U780 ( .A(G137), .B(n731), .Z(G39) );
  XOR2_X1 U781 ( .A(n732), .B(G131), .Z(G33) );
endmodule

