//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958;
  INV_X1    g000(.A(KEYINPUT2), .ZN(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  INV_X1    g002(.A(G162gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  INV_X1    g005(.A(G148gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(G141gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT74), .ZN(new_n209));
  AOI22_X1  g008(.A1(new_n205), .A2(new_n206), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G141gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G148gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n207), .A2(G141gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT74), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n211), .A2(G148gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n202), .B1(new_n208), .B2(new_n215), .ZN(new_n216));
  AND2_X1   g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n210), .A2(new_n214), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  OR2_X1    g020(.A1(G211gat), .A2(G218gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(G211gat), .A2(G218gat), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT69), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT22), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT22), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT69), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(new_n228), .A3(new_n223), .ZN(new_n229));
  XNOR2_X1  g028(.A(G197gat), .B(G204gat), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n224), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n224), .B1(new_n229), .B2(new_n230), .ZN(new_n232));
  NOR3_X1   g031(.A1(new_n231), .A2(new_n232), .A3(KEYINPUT29), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n221), .B1(new_n233), .B2(KEYINPUT3), .ZN(new_n234));
  NAND2_X1  g033(.A1(G228gat), .A2(G233gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n205), .A2(new_n206), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n208), .A2(new_n209), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(new_n214), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n239));
  XNOR2_X1  g038(.A(G141gat), .B(G148gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n219), .B1(new_n240), .B2(KEYINPUT2), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n238), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT75), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT75), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n238), .A2(new_n241), .A3(new_n244), .A4(new_n239), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT29), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n222), .A2(KEYINPUT70), .A3(new_n223), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n229), .A2(new_n247), .A3(new_n230), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n247), .B1(new_n229), .B2(new_n230), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n234), .B(new_n235), .C1(new_n246), .C2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT29), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n253), .B1(new_n248), .B2(new_n249), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n220), .B1(new_n254), .B2(new_n239), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n244), .B1(new_n220), .B2(new_n239), .ZN(new_n256));
  INV_X1    g055(.A(new_n245), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n253), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n255), .B1(new_n258), .B2(new_n250), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n252), .B1(new_n259), .B2(new_n235), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G22gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n235), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n243), .A2(new_n245), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n251), .B1(new_n263), .B2(new_n253), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n262), .B1(new_n264), .B2(new_n255), .ZN(new_n265));
  INV_X1    g064(.A(G22gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(new_n266), .A3(new_n252), .ZN(new_n267));
  XNOR2_X1  g066(.A(G78gat), .B(G106gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT31), .B(G50gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n270), .B(KEYINPUT77), .Z(new_n271));
  AND4_X1   g070(.A1(KEYINPUT78), .A2(new_n261), .A3(new_n267), .A4(new_n271), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n265), .A2(new_n266), .A3(new_n252), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n266), .B1(new_n265), .B2(new_n252), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT78), .B1(new_n275), .B2(new_n271), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n272), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G226gat), .A2(G233gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G183gat), .ZN(new_n281));
  INV_X1    g080(.A(G190gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT27), .B(G183gat), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT28), .B1(new_n285), .B2(new_n282), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(KEYINPUT27), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT27), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G183gat), .ZN(new_n289));
  AND4_X1   g088(.A1(KEYINPUT28), .A2(new_n287), .A3(new_n289), .A4(new_n282), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n284), .B1(new_n286), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G169gat), .ZN(new_n292));
  INV_X1    g091(.A(G176gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT64), .ZN(new_n295));
  NAND2_X1  g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n294), .B(new_n295), .C1(new_n297), .C2(KEYINPUT26), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n294), .A2(KEYINPUT26), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT64), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n298), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(G190gat), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT23), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n309), .A2(new_n292), .A3(new_n293), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(new_n297), .B2(new_n311), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n308), .A2(new_n312), .A3(KEYINPUT25), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT25), .B1(new_n308), .B2(new_n312), .ZN(new_n314));
  OAI22_X1  g113(.A1(new_n291), .A2(new_n303), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n280), .B1(new_n315), .B2(new_n253), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT25), .ZN(new_n317));
  NOR3_X1   g116(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n311), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n318), .B1(new_n319), .B2(new_n296), .ZN(new_n320));
  AND3_X1   g119(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n321), .B1(new_n305), .B2(new_n304), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n317), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n308), .A2(new_n312), .A3(KEYINPUT25), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n287), .A2(new_n289), .A3(new_n282), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT28), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n285), .A2(KEYINPUT28), .A3(new_n282), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n298), .A2(new_n299), .A3(new_n302), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(new_n331), .A3(new_n284), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n279), .B1(new_n325), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n250), .B1(new_n316), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n283), .B1(new_n328), .B2(new_n329), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n331), .A2(new_n335), .B1(new_n323), .B2(new_n324), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n279), .B1(new_n336), .B2(KEYINPUT29), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n315), .A2(new_n280), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n251), .A3(new_n338), .ZN(new_n339));
  XOR2_X1   g138(.A(G8gat), .B(G36gat), .Z(new_n340));
  XNOR2_X1  g139(.A(G64gat), .B(G92gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n334), .A2(new_n339), .A3(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT80), .B(KEYINPUT37), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n334), .A2(new_n339), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT81), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT81), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n334), .A2(new_n339), .A3(new_n350), .A4(new_n347), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n316), .A2(new_n250), .A3(new_n333), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n251), .B1(new_n337), .B2(new_n338), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT37), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT79), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT38), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n344), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT37), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n359), .B1(new_n334), .B2(new_n339), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n358), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n352), .A2(new_n356), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n355), .A2(new_n344), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n364), .B1(new_n349), .B2(new_n351), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n346), .B(new_n363), .C1(new_n365), .C2(new_n357), .ZN(new_n366));
  XNOR2_X1  g165(.A(G1gat), .B(G29gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(KEYINPUT0), .ZN(new_n368));
  XNOR2_X1  g167(.A(G57gat), .B(G85gat), .ZN(new_n369));
  XOR2_X1   g168(.A(new_n368), .B(new_n369), .Z(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G134gat), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT65), .B1(new_n372), .B2(G127gat), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT66), .ZN(new_n375));
  XNOR2_X1  g174(.A(G113gat), .B(G120gat), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n374), .B(new_n375), .C1(new_n376), .C2(KEYINPUT1), .ZN(new_n377));
  OAI211_X1 g176(.A(KEYINPUT66), .B(new_n373), .C1(new_n376), .C2(KEYINPUT1), .ZN(new_n378));
  XNOR2_X1  g177(.A(G127gat), .B(G134gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n377), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n380), .B1(new_n377), .B2(new_n378), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n221), .A2(KEYINPUT3), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n263), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n220), .B1(new_n381), .B2(new_n382), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g187(.A(KEYINPUT4), .B(new_n220), .C1(new_n381), .C2(new_n382), .ZN(new_n389));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n385), .A2(new_n388), .A3(new_n389), .A4(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT5), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n378), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n379), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n378), .A3(new_n380), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(new_n221), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n386), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n390), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n392), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n391), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n392), .A3(new_n390), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n394), .A2(new_n395), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT4), .B1(new_n403), .B2(new_n220), .ZN(new_n404));
  INV_X1    g203(.A(new_n389), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT76), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT76), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n388), .A2(new_n407), .A3(new_n389), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n402), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n371), .B1(new_n401), .B2(new_n409), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n388), .A2(new_n407), .A3(new_n389), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n407), .B1(new_n388), .B2(new_n389), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n400), .B(new_n370), .C1(new_n413), .C2(new_n402), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n410), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  OAI211_X1 g215(.A(KEYINPUT6), .B(new_n371), .C1(new_n401), .C2(new_n409), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n278), .B1(new_n366), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT30), .ZN(new_n420));
  OR2_X1    g219(.A1(new_n346), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n344), .B1(new_n353), .B2(new_n354), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n346), .A2(KEYINPUT73), .A3(new_n420), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT73), .B1(new_n346), .B2(new_n420), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n421), .B(new_n422), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n397), .A2(new_n398), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT39), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n263), .A2(new_n383), .A3(new_n384), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n429), .B1(new_n406), .B2(new_n408), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n428), .B1(new_n430), .B2(new_n390), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n385), .B1(new_n411), .B2(new_n412), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n432), .A2(new_n427), .A3(new_n398), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n431), .A2(new_n433), .A3(KEYINPUT40), .A4(new_n370), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n425), .A2(new_n434), .A3(new_n410), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n431), .A2(new_n433), .A3(new_n370), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT40), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n419), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n291), .A2(new_n303), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n313), .A2(new_n314), .ZN(new_n442));
  OAI22_X1  g241(.A1(new_n441), .A2(new_n442), .B1(new_n381), .B2(new_n382), .ZN(new_n443));
  INV_X1    g242(.A(G227gat), .ZN(new_n444));
  INV_X1    g243(.A(G233gat), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n394), .A2(new_n325), .A3(new_n332), .A4(new_n395), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n443), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT32), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT33), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  XOR2_X1   g250(.A(G15gat), .B(G43gat), .Z(new_n452));
  XNOR2_X1  g251(.A(new_n452), .B(KEYINPUT67), .ZN(new_n453));
  XOR2_X1   g252(.A(G71gat), .B(G99gat), .Z(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n449), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n455), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n448), .B(KEYINPUT32), .C1(new_n450), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT34), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n447), .ZN(new_n461));
  INV_X1    g260(.A(new_n446), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AOI211_X1 g262(.A(KEYINPUT34), .B(new_n446), .C1(new_n443), .C2(new_n447), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n459), .A2(KEYINPUT68), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n447), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n394), .A2(new_n395), .B1(new_n325), .B2(new_n332), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT34), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n461), .A2(new_n460), .A3(new_n462), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT68), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT68), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n473), .B1(new_n463), .B2(new_n464), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n472), .A2(new_n474), .A3(new_n458), .A4(new_n456), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n466), .A2(new_n475), .A3(KEYINPUT36), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n466), .A2(new_n475), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT36), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n425), .B1(new_n416), .B2(new_n417), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n476), .B(new_n479), .C1(new_n480), .C2(new_n278), .ZN(new_n481));
  INV_X1    g280(.A(new_n425), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n418), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n261), .A2(new_n267), .A3(new_n271), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT78), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n277), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n275), .A2(KEYINPUT78), .A3(new_n271), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n477), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n483), .A2(new_n488), .A3(KEYINPUT35), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT35), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n477), .A2(new_n486), .A3(new_n487), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n490), .B1(new_n491), .B2(new_n480), .ZN(new_n492));
  OAI22_X1  g291(.A1(new_n440), .A2(new_n481), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(G232gat), .A2(G233gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n494), .A2(KEYINPUT41), .ZN(new_n495));
  XNOR2_X1  g294(.A(G134gat), .B(G162gat), .ZN(new_n496));
  XOR2_X1   g295(.A(new_n495), .B(new_n496), .Z(new_n497));
  INV_X1    g296(.A(KEYINPUT93), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT84), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT82), .B1(G29gat), .B2(G36gat), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT14), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n502), .A2(new_n503), .B1(G29gat), .B2(G36gat), .ZN(new_n504));
  OR3_X1    g303(.A1(KEYINPUT82), .A2(G29gat), .A3(G36gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n505), .A2(KEYINPUT14), .A3(new_n501), .ZN(new_n506));
  INV_X1    g305(.A(G43gat), .ZN(new_n507));
  INV_X1    g306(.A(G50gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G43gat), .A2(G50gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT15), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT15), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n509), .A2(new_n513), .A3(new_n510), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n504), .A2(new_n506), .A3(new_n512), .A4(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n512), .B1(new_n504), .B2(new_n506), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n515), .B1(new_n516), .B2(KEYINPUT83), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n512), .A2(new_n514), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT83), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n518), .A2(new_n519), .A3(new_n506), .A4(new_n504), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n500), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n517), .A2(new_n520), .A3(new_n500), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(G99gat), .ZN(new_n525));
  INV_X1    g324(.A(G106gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G99gat), .A2(G106gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT90), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n527), .A2(KEYINPUT90), .A3(new_n528), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(G85gat), .ZN(new_n534));
  INV_X1    g333(.A(G92gat), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT88), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT88), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(G85gat), .A3(G92gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n538), .A3(KEYINPUT7), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n528), .A2(KEYINPUT8), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT89), .B(G85gat), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n539), .B(new_n540), .C1(G92gat), .C2(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT7), .B1(new_n536), .B2(new_n538), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n533), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n541), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n545), .A2(new_n535), .B1(KEYINPUT8), .B2(new_n528), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n532), .ZN(new_n547));
  INV_X1    g346(.A(new_n543), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n546), .A2(new_n547), .A3(new_n548), .A4(new_n539), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n544), .A2(KEYINPUT91), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT91), .B1(new_n544), .B2(new_n549), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n524), .A2(new_n553), .B1(KEYINPUT41), .B2(new_n494), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT17), .ZN(new_n555));
  INV_X1    g354(.A(new_n523), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n555), .B1(new_n556), .B2(new_n521), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n517), .A2(new_n520), .A3(KEYINPUT17), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n544), .A2(new_n549), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT91), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n550), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n557), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT92), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n554), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G190gat), .B(G218gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n564), .B1(new_n554), .B2(new_n563), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI211_X1 g368(.A(new_n564), .B(new_n566), .C1(new_n554), .C2(new_n563), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n499), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n568), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n572), .A2(new_n565), .A3(new_n566), .ZN(new_n573));
  INV_X1    g372(.A(new_n570), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n497), .B(new_n498), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT9), .ZN(new_n578));
  INV_X1    g377(.A(G71gat), .ZN(new_n579));
  INV_X1    g378(.A(G78gat), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G57gat), .A2(G64gat), .ZN(new_n582));
  OR2_X1    g381(.A1(G57gat), .A2(G64gat), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n579), .A2(new_n580), .ZN(new_n585));
  AOI22_X1  g384(.A1(KEYINPUT86), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n585), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n588), .A2(new_n581), .A3(new_n582), .A4(new_n583), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT21), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(G127gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n590), .B(KEYINPUT87), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT21), .ZN(new_n597));
  XNOR2_X1  g396(.A(G15gat), .B(G22gat), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT16), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n598), .B1(new_n599), .B2(G1gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n600), .B1(G1gat), .B2(new_n598), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n601), .B(G8gat), .Z(new_n602));
  NAND2_X1  g401(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n595), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(G155gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(G183gat), .B(G211gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n604), .B(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n577), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n602), .B1(new_n522), .B2(new_n523), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n602), .A2(new_n558), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n611), .B1(new_n557), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G229gat), .A2(G233gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n615), .B(KEYINPUT85), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n614), .A2(KEYINPUT18), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n602), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n619), .B1(new_n556), .B2(new_n521), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT17), .B1(new_n522), .B2(new_n523), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n617), .B(new_n620), .C1(new_n621), .C2(new_n612), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT18), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n616), .B(KEYINPUT13), .Z(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n524), .A2(new_n619), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(new_n627), .B2(new_n611), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n618), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G113gat), .B(G141gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G197gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT11), .B(G169gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n629), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n618), .A2(new_n624), .A3(new_n634), .A4(new_n628), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(G230gat), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n639), .A2(new_n445), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n561), .A2(KEYINPUT10), .A3(new_n596), .A4(new_n550), .ZN(new_n641));
  INV_X1    g440(.A(new_n590), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n533), .A2(KEYINPUT94), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n559), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n544), .A2(new_n642), .A3(new_n549), .A4(new_n643), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n640), .B1(new_n641), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n645), .A2(new_n647), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n640), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(G120gat), .B(G148gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT95), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n650), .A2(new_n652), .A3(new_n657), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  AND4_X1   g461(.A1(new_n493), .A2(new_n610), .A3(new_n638), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT96), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(new_n418), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g465(.A1(new_n664), .A2(new_n482), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n667), .A2(KEYINPUT97), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(KEYINPUT97), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n668), .A2(G8gat), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT16), .B(G8gat), .Z(new_n671));
  NAND3_X1  g470(.A1(new_n667), .A2(KEYINPUT42), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n671), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n673), .B1(new_n668), .B2(new_n669), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n670), .B(new_n672), .C1(new_n674), .C2(KEYINPUT42), .ZN(G1325gat));
  NAND2_X1  g474(.A1(new_n479), .A2(new_n476), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(G15gat), .B1(new_n664), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n477), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n679), .A2(G15gat), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n678), .B1(new_n664), .B2(new_n680), .ZN(G1326gat));
  NOR2_X1   g480(.A1(new_n664), .A2(new_n278), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT43), .B(G22gat), .Z(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1327gat));
  INV_X1    g483(.A(new_n609), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n636), .A2(new_n637), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n685), .A2(new_n686), .A3(new_n661), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n493), .A2(new_n577), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(G29gat), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n688), .A2(new_n689), .A3(new_n416), .A4(new_n417), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT98), .B(KEYINPUT45), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n493), .A2(KEYINPUT44), .A3(new_n577), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n687), .B(KEYINPUT99), .Z(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n577), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n440), .A2(KEYINPUT100), .A3(new_n481), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT100), .ZN(new_n699));
  INV_X1    g498(.A(new_n278), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n676), .B1(new_n483), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n436), .A2(new_n437), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n702), .A2(new_n410), .A3(new_n425), .A4(new_n434), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n703), .B(new_n278), .C1(new_n418), .C2(new_n366), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n699), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n698), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT101), .B1(new_n489), .B2(new_n492), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT35), .B1(new_n483), .B2(new_n488), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n491), .A2(new_n490), .A3(new_n480), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT101), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n697), .B1(new_n706), .B2(new_n712), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n694), .B(new_n696), .C1(new_n713), .C2(KEYINPUT44), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n418), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n692), .B1(new_n715), .B2(new_n689), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n716), .B(KEYINPUT102), .Z(G1328gat));
  INV_X1    g516(.A(G36gat), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n688), .A2(new_n718), .A3(new_n425), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(KEYINPUT46), .Z(new_n720));
  NOR2_X1   g519(.A1(new_n714), .A2(new_n482), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n721), .A2(KEYINPUT103), .ZN(new_n722));
  OAI21_X1  g521(.A(G36gat), .B1(new_n721), .B2(KEYINPUT103), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n720), .B1(new_n722), .B2(new_n723), .ZN(G1329gat));
  NAND3_X1  g523(.A1(new_n688), .A2(new_n507), .A3(new_n477), .ZN(new_n725));
  OAI21_X1  g524(.A(KEYINPUT100), .B1(new_n440), .B2(new_n481), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n701), .A2(new_n704), .A3(new_n699), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n726), .A2(new_n727), .A3(new_n711), .A4(new_n707), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT44), .B1(new_n728), .B2(new_n577), .ZN(new_n729));
  NOR4_X1   g528(.A1(new_n729), .A2(new_n677), .A3(new_n693), .A4(new_n695), .ZN(new_n730));
  OAI211_X1 g529(.A(KEYINPUT47), .B(new_n725), .C1(new_n730), .C2(new_n507), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n730), .B2(new_n507), .ZN(new_n733));
  OAI211_X1 g532(.A(KEYINPUT104), .B(G43gat), .C1(new_n714), .C2(new_n677), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(new_n734), .A3(new_n725), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n736), .B1(new_n735), .B2(new_n737), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n731), .B1(new_n738), .B2(new_n739), .ZN(G1330gat));
  OAI21_X1  g539(.A(G50gat), .B1(new_n714), .B2(new_n278), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n700), .A2(new_n508), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT106), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n688), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT48), .Z(G1331gat));
  NAND3_X1  g545(.A1(new_n610), .A2(new_n686), .A3(new_n661), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(KEYINPUT107), .Z(new_n748));
  XNOR2_X1  g547(.A(new_n418), .B(KEYINPUT108), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n748), .A2(new_n728), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g550(.A(new_n482), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n748), .A2(new_n728), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n753), .B(new_n754), .Z(G1333gat));
  AND2_X1   g554(.A1(new_n679), .A2(KEYINPUT109), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n679), .A2(KEYINPUT109), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n756), .A2(new_n757), .A3(G71gat), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n748), .A2(new_n728), .A3(new_n758), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n748), .A2(new_n676), .A3(new_n728), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n760), .B2(new_n579), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(KEYINPUT50), .Z(G1334gat));
  NAND3_X1  g561(.A1(new_n748), .A2(new_n700), .A3(new_n728), .ZN(new_n763));
  XOR2_X1   g562(.A(KEYINPUT110), .B(G78gat), .Z(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(G1335gat));
  NOR2_X1   g564(.A1(new_n729), .A2(new_n693), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n686), .A2(new_n609), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n767), .B(KEYINPUT111), .Z(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n766), .A2(new_n661), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n541), .B1(new_n770), .B2(new_n418), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n713), .A2(new_n769), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT51), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n713), .A2(new_n774), .A3(new_n769), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n773), .A2(new_n661), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n416), .A2(new_n417), .A3(new_n545), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n771), .B1(new_n776), .B2(new_n777), .ZN(G1336gat));
  INV_X1    g577(.A(new_n776), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n482), .A2(G92gat), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT52), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n770), .A2(new_n482), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n782), .A2(KEYINPUT112), .ZN(new_n783));
  OAI21_X1  g582(.A(G92gat), .B1(new_n782), .B2(KEYINPUT112), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n782), .A2(new_n535), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n776), .A2(G92gat), .A3(new_n482), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT52), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(G1337gat));
  NOR3_X1   g588(.A1(new_n770), .A2(new_n525), .A3(new_n677), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n779), .A2(new_n477), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n791), .B2(new_n525), .ZN(G1338gat));
  OAI21_X1  g591(.A(G106gat), .B1(new_n770), .B2(new_n278), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n278), .A2(G106gat), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n776), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n641), .A2(new_n648), .A3(new_n640), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n799), .A2(new_n649), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n641), .A2(new_n648), .ZN(new_n802));
  INV_X1    g601(.A(new_n640), .ZN(new_n803));
  XOR2_X1   g602(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n804));
  NAND3_X1  g603(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n658), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n798), .B1(new_n801), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n641), .A2(new_n648), .A3(new_n640), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n650), .A2(KEYINPUT54), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n657), .B1(new_n649), .B2(new_n804), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(KEYINPUT55), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n807), .A2(new_n660), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n807), .A2(new_n811), .A3(KEYINPUT114), .A4(new_n660), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(new_n638), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n627), .A2(new_n611), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n620), .B1(new_n621), .B2(new_n612), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n818), .A2(new_n625), .B1(new_n819), .B2(new_n616), .ZN(new_n820));
  INV_X1    g619(.A(new_n633), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n817), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n614), .A2(new_n617), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n627), .A2(new_n611), .A3(new_n626), .ZN(new_n824));
  OAI211_X1 g623(.A(KEYINPUT115), .B(new_n633), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n822), .A2(new_n661), .A3(new_n825), .A4(new_n637), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n577), .B1(new_n816), .B2(new_n826), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n822), .A2(new_n637), .A3(new_n825), .ZN(new_n828));
  AND4_X1   g627(.A1(new_n577), .A2(new_n828), .A3(new_n814), .A4(new_n815), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n609), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NOR4_X1   g629(.A1(new_n577), .A2(new_n609), .A3(new_n638), .A4(new_n661), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n488), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n833), .A2(new_n416), .A3(new_n417), .A4(new_n482), .ZN(new_n834));
  INV_X1    g633(.A(G113gat), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n834), .A2(new_n835), .A3(new_n686), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n833), .A2(new_n749), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n837), .A2(new_n482), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n638), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n836), .B1(new_n839), .B2(new_n835), .ZN(G1340gat));
  NOR2_X1   g639(.A1(new_n662), .A2(G120gat), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT116), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G120gat), .B1(new_n834), .B2(new_n662), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(G1341gat));
  INV_X1    g644(.A(G127gat), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n838), .A2(new_n846), .A3(new_n685), .ZN(new_n847));
  OAI21_X1  g646(.A(G127gat), .B1(new_n834), .B2(new_n609), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(G1342gat));
  NAND2_X1  g648(.A1(new_n577), .A2(new_n482), .ZN(new_n850));
  XOR2_X1   g649(.A(new_n850), .B(KEYINPUT117), .Z(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n372), .A3(new_n852), .ZN(new_n853));
  XOR2_X1   g652(.A(new_n853), .B(KEYINPUT56), .Z(new_n854));
  OAI21_X1  g653(.A(G134gat), .B1(new_n834), .B2(new_n697), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(G1343gat));
  AOI21_X1  g655(.A(new_n278), .B1(new_n830), .B2(new_n832), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n826), .B1(new_n686), .B2(new_n812), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n697), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n577), .A2(new_n828), .A3(new_n814), .A4(new_n815), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n831), .B1(new_n863), .B2(new_n609), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT57), .B1(new_n864), .B2(new_n278), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n676), .A2(new_n418), .A3(new_n425), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n859), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(G141gat), .B1(new_n867), .B2(new_n686), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n857), .A2(new_n677), .A3(new_n749), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n482), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n638), .A2(new_n211), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT118), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n868), .B(KEYINPUT119), .C1(new_n870), .C2(new_n872), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(G148gat), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n859), .A2(new_n865), .A3(new_n866), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(new_n661), .ZN(new_n878));
  INV_X1    g677(.A(new_n812), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n577), .A2(new_n879), .A3(new_n828), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n685), .B1(new_n861), .B2(new_n880), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n858), .B(new_n700), .C1(new_n881), .C2(new_n831), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n866), .A2(new_n661), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n882), .B(new_n883), .C1(new_n857), .C2(new_n858), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(G148gat), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(KEYINPUT59), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(KEYINPUT120), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n885), .A2(new_n888), .A3(KEYINPUT59), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n878), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n870), .A2(G148gat), .A3(new_n662), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT121), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n893));
  INV_X1    g692(.A(new_n891), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n888), .B1(new_n885), .B2(KEYINPUT59), .ZN(new_n895));
  AOI211_X1 g694(.A(KEYINPUT120), .B(new_n875), .C1(new_n884), .C2(G148gat), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n893), .B(new_n894), .C1(new_n897), .C2(new_n878), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n892), .A2(new_n898), .ZN(G1345gat));
  OAI21_X1  g698(.A(G155gat), .B1(new_n867), .B2(new_n609), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n685), .A2(new_n203), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n870), .B2(new_n901), .ZN(G1346gat));
  OAI21_X1  g701(.A(G162gat), .B1(new_n867), .B2(new_n697), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n869), .A2(new_n204), .A3(new_n852), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1347gat));
  NAND2_X1  g704(.A1(new_n830), .A2(new_n832), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n906), .A2(new_n418), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n488), .A2(new_n482), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(G169gat), .B1(new_n909), .B2(new_n638), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n756), .A2(new_n757), .A3(new_n482), .ZN(new_n911));
  INV_X1    g710(.A(new_n749), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT122), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n913), .A2(KEYINPUT122), .ZN(new_n915));
  AND4_X1   g714(.A1(new_n278), .A2(new_n906), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n686), .A2(new_n292), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n910), .B1(new_n916), .B2(new_n917), .ZN(G1348gat));
  NAND3_X1  g717(.A1(new_n916), .A2(G176gat), .A3(new_n661), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n907), .A2(new_n661), .A3(new_n908), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n920), .A2(KEYINPUT123), .A3(new_n293), .ZN(new_n921));
  AOI21_X1  g720(.A(KEYINPUT123), .B1(new_n920), .B2(new_n293), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT124), .ZN(G1349gat));
  AOI21_X1  g723(.A(new_n281), .B1(new_n916), .B2(new_n685), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n685), .A2(new_n285), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n925), .B1(new_n909), .B2(new_n926), .ZN(new_n927));
  XOR2_X1   g726(.A(new_n927), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g727(.A(new_n282), .B1(new_n916), .B2(new_n577), .ZN(new_n929));
  XOR2_X1   g728(.A(new_n929), .B(KEYINPUT61), .Z(new_n930));
  NAND3_X1  g729(.A1(new_n909), .A2(new_n282), .A3(new_n577), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1351gat));
  NOR2_X1   g731(.A1(new_n676), .A2(new_n482), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n907), .A2(new_n700), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(G197gat), .B1(new_n934), .B2(new_n638), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n882), .B1(new_n857), .B2(new_n858), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n936), .A2(KEYINPUT125), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n912), .A2(new_n933), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n938), .B1(new_n936), .B2(KEYINPUT125), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n638), .A2(G197gat), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n935), .B1(new_n940), .B2(new_n941), .ZN(G1352gat));
  INV_X1    g741(.A(G204gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n934), .A2(new_n943), .A3(new_n661), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT62), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n943), .B1(new_n940), .B2(new_n661), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n945), .A2(new_n946), .ZN(G1353gat));
  INV_X1    g746(.A(G211gat), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n934), .A2(new_n948), .A3(new_n685), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT126), .ZN(new_n950));
  OR3_X1    g749(.A1(new_n936), .A2(new_n609), .A3(new_n938), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  OR3_X1    g751(.A1(new_n952), .A2(KEYINPUT63), .A3(new_n948), .ZN(new_n953));
  OAI21_X1  g752(.A(KEYINPUT63), .B1(new_n952), .B2(new_n948), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n950), .A2(new_n953), .A3(new_n954), .ZN(G1354gat));
  AOI21_X1  g754(.A(G218gat), .B1(new_n934), .B2(new_n577), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n577), .A2(G218gat), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT127), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n956), .B1(new_n940), .B2(new_n958), .ZN(G1355gat));
endmodule


