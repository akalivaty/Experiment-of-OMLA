//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 1 0 1 1 1 1 0 1 0 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n817, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n968, new_n969, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1027, new_n1028;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  AND2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT2), .ZN(new_n207));
  OR2_X1    g006(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G148gat), .ZN(new_n209));
  OR2_X1    g008(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(G141gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n206), .B(new_n208), .C1(new_n212), .C2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n209), .A2(G141gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n207), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n204), .A2(new_n205), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G218gat), .ZN(new_n221));
  AND2_X1   g020(.A1(KEYINPUT71), .A2(KEYINPUT22), .ZN(new_n222));
  NOR2_X1   g021(.A1(KEYINPUT71), .A2(KEYINPUT22), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT72), .B(G211gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(new_n221), .ZN(new_n226));
  INV_X1    g025(.A(G211gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(G197gat), .B(G204gat), .ZN(new_n228));
  AND3_X1   g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n227), .B1(new_n226), .B2(new_n228), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n221), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  AND2_X1   g030(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n233));
  NOR3_X1   g032(.A1(new_n232), .A2(new_n233), .A3(new_n221), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT71), .B(KEYINPUT22), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n228), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G211gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(G218gat), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT29), .B1(new_n231), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n220), .B1(new_n240), .B2(KEYINPUT3), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT73), .ZN(new_n242));
  NOR3_X1   g041(.A1(new_n229), .A2(new_n230), .A3(new_n221), .ZN(new_n243));
  AOI21_X1  g042(.A(G218gat), .B1(new_n237), .B2(new_n238), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n231), .A2(KEYINPUT73), .A3(new_n239), .ZN(new_n246));
  AND2_X1   g045(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n248));
  OAI21_X1  g047(.A(G148gat), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n218), .B1(new_n249), .B2(new_n213), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n250), .A2(new_n208), .B1(new_n218), .B2(new_n217), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT29), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n245), .A2(new_n246), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G50gat), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n241), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n257), .B1(new_n241), .B2(new_n256), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT31), .B(G22gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(G228gat), .A2(G233gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  NOR3_X1   g061(.A1(new_n258), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n262), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n245), .A2(new_n246), .A3(new_n255), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n254), .B1(new_n243), .B2(new_n244), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n251), .B1(new_n266), .B2(new_n252), .ZN(new_n267));
  OAI21_X1  g066(.A(G50gat), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n241), .A2(new_n256), .A3(new_n257), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n264), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n203), .B1(new_n263), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n262), .B1(new_n258), .B2(new_n259), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n268), .A2(new_n269), .A3(new_n264), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n272), .A2(new_n273), .A3(new_n202), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G227gat), .ZN(new_n276));
  INV_X1    g075(.A(G233gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  AND3_X1   g078(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT24), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT64), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT64), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n282), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT23), .ZN(new_n291));
  INV_X1    g090(.A(G169gat), .ZN(new_n292));
  INV_X1    g091(.A(G176gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n294), .A2(new_n295), .B1(G169gat), .B2(G176gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n290), .A2(KEYINPUT25), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT25), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(new_n295), .ZN(new_n299));
  NAND2_X1  g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR3_X1   g100(.A1(new_n280), .A2(new_n287), .A3(new_n281), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n298), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT26), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n292), .A2(new_n293), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(KEYINPUT66), .A3(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n309), .B1(new_n305), .B2(new_n300), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT66), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n311), .B1(new_n309), .B2(new_n305), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n308), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  AND2_X1   g112(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT28), .B1(new_n316), .B2(G190gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT65), .ZN(new_n318));
  INV_X1    g117(.A(G183gat), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT27), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n321));
  INV_X1    g120(.A(G190gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT27), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n323), .A2(KEYINPUT65), .A3(G183gat), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n320), .A2(new_n321), .A3(new_n322), .A4(new_n324), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n313), .A2(new_n283), .A3(new_n317), .A4(new_n325), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n304), .A2(KEYINPUT68), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT68), .B1(new_n304), .B2(new_n326), .ZN(new_n328));
  AND2_X1   g127(.A1(KEYINPUT67), .A2(G127gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(G113gat), .B(G120gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n329), .B1(new_n330), .B2(KEYINPUT1), .ZN(new_n331));
  INV_X1    g130(.A(G134gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT1), .ZN(new_n333));
  INV_X1    g132(.A(G127gat), .ZN(new_n334));
  INV_X1    g133(.A(G113gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n335), .A2(G120gat), .ZN(new_n336));
  INV_X1    g135(.A(G120gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n337), .A2(G113gat), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n333), .B(new_n334), .C1(new_n336), .C2(new_n338), .ZN(new_n339));
  AND3_X1   g138(.A1(new_n331), .A2(new_n332), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n332), .B1(new_n331), .B2(new_n339), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n327), .A2(new_n328), .A3(new_n342), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n317), .A2(new_n283), .A3(new_n325), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n344), .A2(new_n313), .B1(new_n297), .B2(new_n303), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n345), .A2(KEYINPUT68), .A3(new_n342), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n279), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT34), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT68), .ZN(new_n351));
  INV_X1    g150(.A(new_n281), .ZN(new_n352));
  NAND3_X1  g151(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(new_n285), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT25), .B1(new_n296), .B2(new_n354), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n283), .A2(new_n288), .A3(new_n284), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n288), .B1(new_n283), .B2(new_n284), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n298), .B1(new_n358), .B2(new_n282), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n355), .B1(new_n359), .B2(new_n296), .ZN(new_n360));
  AND4_X1   g159(.A1(new_n313), .A2(new_n283), .A3(new_n317), .A4(new_n325), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n351), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n341), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n331), .A2(new_n332), .A3(new_n339), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n304), .A2(new_n326), .A3(KEYINPUT68), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n362), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n346), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n368), .A2(KEYINPUT34), .A3(new_n279), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n367), .A2(new_n278), .A3(new_n346), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT32), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT33), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G71gat), .B(G99gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(KEYINPUT69), .ZN(new_n375));
  XOR2_X1   g174(.A(G15gat), .B(G43gat), .Z(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n371), .A2(new_n373), .A3(new_n378), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n370), .B(KEYINPUT32), .C1(new_n372), .C2(new_n377), .ZN(new_n380));
  AOI221_X4 g179(.A(KEYINPUT70), .B1(new_n350), .B2(new_n369), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n350), .A2(new_n369), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n379), .A2(new_n380), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT70), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n275), .B(KEYINPUT35), .C1(new_n381), .C2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n251), .B1(new_n340), .B2(new_n341), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT4), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT78), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n251), .B(KEYINPUT78), .C1(new_n340), .C2(new_n341), .ZN(new_n393));
  NAND2_X1  g192(.A1(G225gat), .A2(G233gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT4), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT77), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n215), .A2(new_n219), .A3(new_n252), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n252), .B1(new_n215), .B2(new_n219), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n397), .B1(new_n400), .B2(new_n342), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n220), .A2(KEYINPUT3), .ZN(new_n402));
  AND4_X1   g201(.A1(new_n397), .A2(new_n342), .A3(new_n253), .A4(new_n402), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n390), .B(new_n396), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT5), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n342), .A2(new_n220), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n392), .A2(new_n393), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n394), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n342), .A2(new_n253), .A3(new_n402), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT77), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n400), .A2(new_n397), .A3(new_n342), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT78), .B1(new_n365), .B2(new_n251), .ZN(new_n415));
  INV_X1    g214(.A(new_n393), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT4), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OR2_X1    g216(.A1(new_n389), .A2(KEYINPUT4), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n408), .A2(KEYINPUT5), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n414), .A2(new_n417), .A3(new_n418), .A4(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n410), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G57gat), .B(G85gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(G29gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT80), .B(G1gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  NAND2_X1  g226(.A1(new_n421), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429));
  INV_X1    g228(.A(new_n427), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n410), .A2(new_n430), .A3(new_n420), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n428), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n421), .A2(KEYINPUT6), .A3(new_n427), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n304), .A2(new_n326), .ZN(new_n434));
  NAND2_X1  g233(.A1(G226gat), .A2(G233gat), .ZN(new_n435));
  XOR2_X1   g234(.A(new_n435), .B(KEYINPUT74), .Z(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n435), .B1(new_n345), .B2(KEYINPUT29), .ZN(new_n438));
  INV_X1    g237(.A(new_n246), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT73), .B1(new_n231), .B2(new_n239), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n437), .B(new_n438), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n436), .B1(new_n434), .B2(new_n254), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n345), .A2(new_n435), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n246), .B(new_n245), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n441), .A2(new_n444), .A3(KEYINPUT30), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT30), .B1(new_n441), .B2(new_n444), .ZN(new_n446));
  XNOR2_X1  g245(.A(G64gat), .B(G92gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(G36gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n448), .B(KEYINPUT75), .ZN(new_n449));
  INV_X1    g248(.A(G8gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  OR3_X1    g250(.A1(new_n445), .A2(new_n446), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n441), .A2(new_n444), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT30), .ZN(new_n454));
  INV_X1    g253(.A(new_n451), .ZN(new_n455));
  NOR3_X1   g254(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n432), .A2(new_n433), .B1(new_n452), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT35), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n432), .A2(new_n433), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n445), .A2(new_n446), .A3(new_n451), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(new_n456), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n383), .A2(new_n382), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT34), .B1(new_n368), .B2(new_n279), .ZN(new_n465));
  AOI211_X1 g264(.A(new_n349), .B(new_n278), .C1(new_n367), .C2(new_n346), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n467), .A2(new_n379), .A3(new_n380), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n460), .A2(new_n463), .A3(new_n275), .A4(new_n469), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n387), .A2(new_n458), .B1(new_n459), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT40), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT39), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n407), .A2(new_n408), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n414), .A2(new_n417), .A3(new_n418), .ZN(new_n475));
  AOI211_X1 g274(.A(new_n473), .B(new_n474), .C1(new_n475), .C2(new_n408), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(new_n473), .A3(new_n408), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n430), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n472), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n475), .A2(new_n408), .ZN(new_n480));
  INV_X1    g279(.A(new_n474), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(KEYINPUT39), .A3(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n482), .A2(KEYINPUT40), .A3(new_n430), .A4(new_n477), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n462), .A2(new_n479), .A3(new_n428), .A4(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT37), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n441), .A2(new_n444), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT82), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT82), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n441), .A2(new_n444), .A3(new_n488), .A4(new_n485), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI22_X1  g289(.A1(new_n439), .A2(new_n440), .B1(new_n442), .B2(new_n443), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT81), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n438), .A2(new_n245), .A3(new_n246), .A4(new_n437), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n491), .A2(new_n492), .A3(new_n493), .A4(KEYINPUT37), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n494), .A2(new_n451), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT38), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n491), .A2(KEYINPUT37), .A3(new_n493), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT81), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n490), .A2(new_n495), .A3(new_n496), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n453), .A2(new_n496), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n455), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n499), .A2(new_n432), .A3(new_n433), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n453), .A2(KEYINPUT37), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n496), .B1(new_n490), .B2(new_n503), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n484), .B(new_n275), .C1(new_n502), .C2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n463), .A2(new_n460), .ZN(new_n506));
  INV_X1    g305(.A(new_n275), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT36), .B1(new_n381), .B2(new_n385), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT36), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n464), .A2(new_n510), .A3(new_n468), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n505), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n471), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G57gat), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n515), .A2(G64gat), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n515), .A2(G64gat), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT9), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G71gat), .ZN(new_n519));
  INV_X1    g318(.A(G78gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(G71gat), .A2(G78gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  XOR2_X1   g323(.A(KEYINPUT86), .B(G57gat), .Z(new_n525));
  AOI21_X1  g324(.A(new_n516), .B1(new_n525), .B2(G64gat), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n521), .B1(KEYINPUT9), .B2(new_n522), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(KEYINPUT87), .B(KEYINPUT21), .Z(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(G231gat), .A2(G233gat), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n530), .B(new_n531), .Z(new_n532));
  XOR2_X1   g331(.A(G183gat), .B(G211gat), .Z(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT89), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT20), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n532), .B(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G15gat), .B(G22gat), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n540), .A2(G1gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT16), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n540), .B1(new_n542), .B2(G1gat), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n541), .A2(new_n450), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n450), .B1(new_n541), .B2(new_n543), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT21), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n528), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT90), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NOR3_X1   g350(.A1(new_n547), .A2(KEYINPUT90), .A3(new_n549), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n539), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OR3_X1    g352(.A1(new_n547), .A2(KEYINPUT90), .A3(new_n549), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(new_n550), .A3(new_n538), .ZN(new_n555));
  XNOR2_X1  g354(.A(G127gat), .B(G155gat), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n553), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n557), .B1(new_n553), .B2(new_n555), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n537), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n553), .A2(new_n555), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(new_n556), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(new_n536), .A3(new_n558), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n257), .A2(G43gat), .ZN(new_n566));
  INV_X1    g365(.A(G43gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(G50gat), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n568), .A3(KEYINPUT15), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT83), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(G29gat), .ZN(new_n572));
  INV_X1    g371(.A(G36gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(new_n573), .A3(KEYINPUT14), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT14), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n575), .B1(G29gat), .B2(G36gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(G29gat), .A2(G36gat), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n566), .A2(new_n568), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT15), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n566), .A2(new_n568), .A3(KEYINPUT83), .A4(KEYINPUT15), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n571), .A2(new_n578), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT84), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n578), .A2(new_n569), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT15), .B1(new_n566), .B2(new_n568), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT84), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n588), .A2(new_n589), .A3(new_n571), .A4(new_n582), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n584), .A2(new_n585), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT17), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n584), .A2(KEYINPUT17), .A3(new_n585), .A4(new_n590), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT91), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT7), .ZN(new_n596));
  NAND2_X1  g395(.A1(G85gat), .A2(G92gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G99gat), .A2(G106gat), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT92), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(KEYINPUT92), .A2(G99gat), .A3(G106gat), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(KEYINPUT8), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT93), .ZN(new_n605));
  NOR2_X1   g404(.A1(G85gat), .A2(G92gat), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n605), .B1(new_n604), .B2(new_n607), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n599), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G99gat), .B(G106gat), .Z(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AND3_X1   g411(.A1(KEYINPUT92), .A2(G99gat), .A3(G106gat), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT92), .B1(G99gat), .B2(G106gat), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT8), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT93), .B1(new_n616), .B2(new_n606), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n611), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(new_n620), .A3(new_n599), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n612), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n593), .A2(new_n594), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT94), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n593), .A2(new_n622), .A3(KEYINPUT94), .A4(new_n594), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n591), .A2(new_n621), .A3(new_n612), .ZN(new_n628));
  NAND3_X1  g427(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n628), .A2(KEYINPUT95), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT95), .B1(new_n628), .B2(new_n629), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G134gat), .B(G162gat), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n627), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G190gat), .B(G218gat), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n625), .B(new_n626), .C1(new_n630), .C2(new_n631), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n633), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n635), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n638), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n634), .B1(new_n627), .B2(new_n632), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n639), .A2(new_n633), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n620), .B1(new_n619), .B2(new_n599), .ZN(new_n646));
  AOI211_X1 g445(.A(new_n611), .B(new_n598), .C1(new_n617), .C2(new_n618), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n528), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT10), .ZN(new_n649));
  INV_X1    g448(.A(new_n528), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n612), .A2(new_n621), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n648), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n612), .A2(new_n621), .A3(KEYINPUT10), .A4(new_n650), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(G230gat), .A2(G233gat), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n655), .B1(new_n648), .B2(new_n651), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G120gat), .B(G148gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(new_n293), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n660), .B(G204gat), .Z(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n656), .A2(new_n658), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n655), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n664), .B1(new_n652), .B2(new_n653), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n661), .B1(new_n665), .B2(new_n657), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n565), .A2(new_n641), .A3(new_n645), .A4(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n593), .A2(new_n546), .A3(new_n594), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n547), .A2(new_n591), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(G229gat), .A2(G233gat), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n672), .A2(KEYINPUT85), .A3(KEYINPUT18), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(KEYINPUT13), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n546), .A2(new_n585), .A3(new_n584), .A4(new_n590), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n675), .B1(new_n671), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n670), .A2(new_n671), .A3(new_n673), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT18), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n670), .A2(KEYINPUT18), .A3(new_n671), .A4(new_n673), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT85), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n674), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT11), .B(G169gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(G197gat), .ZN(new_n686));
  XOR2_X1   g485(.A(G113gat), .B(G141gat), .Z(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT12), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n684), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n674), .A2(new_n689), .A3(new_n680), .A4(new_n683), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n669), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n514), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n432), .A2(new_n433), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g498(.A1(new_n695), .A2(new_n463), .ZN(new_n700));
  NAND2_X1  g499(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n542), .A2(new_n450), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT42), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(new_n450), .B2(new_n700), .ZN(G1325gat));
  INV_X1    g504(.A(new_n512), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n696), .A2(G15gat), .A3(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n469), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n695), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n707), .B1(G15gat), .B2(new_n709), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT96), .Z(G1326gat));
  NOR2_X1   g510(.A1(new_n695), .A2(new_n275), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT43), .B(G22gat), .Z(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1327gat));
  INV_X1    g513(.A(KEYINPUT100), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n667), .B(KEYINPUT98), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n717), .A2(new_n693), .A3(new_n565), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n645), .A2(new_n641), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n719), .B1(new_n514), .B2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n720), .ZN(new_n722));
  AOI211_X1 g521(.A(KEYINPUT44), .B(new_n722), .C1(new_n471), .C2(new_n513), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n718), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT99), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI211_X1 g525(.A(KEYINPUT99), .B(new_n718), .C1(new_n721), .C2(new_n723), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n572), .B1(new_n728), .B2(new_n697), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n722), .B1(new_n471), .B2(new_n513), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n460), .A2(G29gat), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n693), .A2(new_n565), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n730), .A2(new_n668), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT97), .ZN(new_n734));
  AOI211_X1 g533(.A(new_n722), .B(new_n667), .C1(new_n471), .C2(new_n513), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT97), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n735), .A2(new_n736), .A3(new_n731), .A4(new_n732), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT45), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n734), .A2(new_n737), .A3(KEYINPUT45), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n715), .B1(new_n729), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n740), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n738), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n460), .B1(new_n726), .B2(new_n727), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n744), .B(KEYINPUT100), .C1(new_n572), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n742), .A2(new_n746), .ZN(G1328gat));
  INV_X1    g546(.A(new_n274), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n202), .B1(new_n272), .B2(new_n273), .ZN(new_n749));
  INV_X1    g548(.A(new_n468), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n467), .B1(new_n380), .B2(new_n379), .ZN(new_n751));
  OAI22_X1  g550(.A1(new_n748), .A2(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n459), .B1(new_n506), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n385), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n383), .A2(new_n384), .A3(new_n382), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n756), .A2(new_n458), .A3(KEYINPUT35), .A4(new_n275), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n508), .A2(new_n512), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n758), .B1(new_n759), .B2(new_n505), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT44), .B1(new_n760), .B2(new_n722), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n730), .A2(new_n719), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(KEYINPUT99), .B1(new_n763), .B2(new_n718), .ZN(new_n764));
  INV_X1    g563(.A(new_n727), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n462), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT101), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT101), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n728), .A2(new_n768), .A3(new_n462), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n767), .A2(G36gat), .A3(new_n769), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n735), .A2(new_n732), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n771), .A2(new_n573), .A3(new_n462), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n772), .B(KEYINPUT46), .Z(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n773), .ZN(G1329gat));
  OAI21_X1  g573(.A(G43gat), .B1(new_n724), .B2(new_n512), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n708), .A2(G43gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n771), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n775), .A2(KEYINPUT47), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n777), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n728), .A2(new_n706), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n779), .B1(new_n780), .B2(G43gat), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n778), .B1(new_n781), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g581(.A1(new_n275), .A2(G50gat), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n771), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n718), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(new_n761), .B2(new_n762), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n786), .A2(KEYINPUT102), .A3(new_n507), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G50gat), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT102), .B1(new_n786), .B2(new_n507), .ZN(new_n789));
  OAI211_X1 g588(.A(KEYINPUT48), .B(new_n784), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n784), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n728), .A2(new_n507), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n791), .B1(new_n792), .B2(G50gat), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n790), .B1(new_n793), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g593(.A(new_n565), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n760), .A2(new_n795), .A3(new_n720), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n691), .A2(new_n692), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n716), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(new_n460), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(new_n525), .ZN(G1332gat));
  NOR2_X1   g600(.A1(new_n799), .A2(new_n463), .ZN(new_n802));
  NOR2_X1   g601(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n803));
  AND2_X1   g602(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n805), .B1(new_n802), .B2(new_n803), .ZN(G1333gat));
  NAND4_X1  g605(.A1(new_n796), .A2(G71gat), .A3(new_n706), .A4(new_n798), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT103), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n469), .B(KEYINPUT104), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n519), .B1(new_n799), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT50), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n808), .A2(new_n814), .A3(new_n811), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(G1334gat));
  NOR2_X1   g615(.A1(new_n799), .A2(new_n275), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(new_n520), .ZN(G1335gat));
  NOR2_X1   g617(.A1(new_n565), .A2(new_n797), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n730), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT51), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT51), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n730), .A2(new_n822), .A3(new_n819), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n821), .A2(new_n667), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(G85gat), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(new_n825), .A3(new_n697), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n797), .A2(new_n565), .A3(new_n668), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n827), .B1(new_n721), .B2(new_n723), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT105), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT105), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n830), .B(new_n827), .C1(new_n721), .C2(new_n723), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n460), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n826), .B1(new_n832), .B2(new_n825), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT106), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI211_X1 g634(.A(KEYINPUT106), .B(new_n826), .C1(new_n832), .C2(new_n825), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(G1336gat));
  OAI21_X1  g636(.A(G92gat), .B1(new_n828), .B2(new_n463), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n716), .A2(G92gat), .A3(new_n463), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n821), .A2(new_n823), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT52), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n829), .A2(new_n831), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n462), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n842), .B1(new_n844), .B2(G92gat), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n822), .A2(KEYINPUT107), .ZN(new_n846));
  XOR2_X1   g645(.A(new_n820), .B(new_n846), .Z(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n839), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n841), .B1(new_n845), .B2(new_n848), .ZN(G1337gat));
  INV_X1    g648(.A(G99gat), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n824), .A2(new_n850), .A3(new_n469), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n512), .B1(new_n829), .B2(new_n831), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n852), .B2(new_n850), .ZN(G1338gat));
  OAI21_X1  g652(.A(G106gat), .B1(new_n828), .B2(new_n275), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n716), .A2(G106gat), .A3(new_n275), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n821), .A2(new_n823), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT53), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n507), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n858), .B1(new_n859), .B2(G106gat), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n847), .A2(new_n855), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n857), .B1(new_n860), .B2(new_n861), .ZN(G1339gat));
  NOR2_X1   g661(.A1(new_n669), .A2(new_n797), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n662), .B1(new_n665), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n652), .A2(new_n653), .A3(new_n664), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT54), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n865), .B(KEYINPUT55), .C1(new_n665), .C2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT55), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n867), .A2(new_n665), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n654), .A2(new_n864), .A3(new_n655), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n661), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n869), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n797), .A2(new_n663), .A3(new_n868), .A4(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n671), .A2(new_n676), .A3(new_n675), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT108), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n673), .B1(new_n670), .B2(new_n671), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n688), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n667), .A2(new_n692), .A3(new_n878), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n879), .A2(new_n641), .A3(new_n645), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n565), .B1(new_n874), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n873), .A2(new_n663), .A3(new_n868), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n692), .A2(new_n878), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n720), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n863), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n460), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n507), .B1(new_n755), .B2(new_n754), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n886), .A2(new_n463), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT109), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n797), .A2(new_n335), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT110), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n886), .A2(new_n463), .A3(new_n275), .A4(new_n469), .ZN(new_n893));
  OAI21_X1  g692(.A(G113gat), .B1(new_n893), .B2(new_n693), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(G1340gat));
  NAND2_X1  g694(.A1(new_n667), .A2(new_n337), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT111), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n889), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(G120gat), .B1(new_n893), .B2(new_n716), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1341gat));
  AOI21_X1  g699(.A(G127gat), .B1(new_n888), .B2(new_n565), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n893), .A2(new_n334), .A3(new_n795), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(new_n902), .ZN(G1342gat));
  XOR2_X1   g702(.A(KEYINPUT67), .B(G134gat), .Z(new_n904));
  NAND3_X1  g703(.A1(new_n888), .A2(new_n720), .A3(new_n904), .ZN(new_n905));
  XOR2_X1   g704(.A(new_n905), .B(KEYINPUT56), .Z(new_n906));
  OAI21_X1  g705(.A(G134gat), .B1(new_n893), .B2(new_n722), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1343gat));
  NOR2_X1   g707(.A1(new_n885), .A2(new_n275), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n460), .B1(new_n509), .B2(new_n511), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT114), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n909), .A2(KEYINPUT114), .A3(new_n910), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n913), .A2(new_n463), .A3(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n693), .A2(G141gat), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT58), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n910), .A2(new_n463), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n693), .A2(new_n882), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n879), .A2(new_n641), .A3(new_n645), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n884), .B(new_n795), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n669), .A2(new_n797), .ZN(new_n923));
  AOI211_X1 g722(.A(new_n919), .B(new_n275), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT113), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n918), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  XOR2_X1   g725(.A(KEYINPUT112), .B(KEYINPUT57), .Z(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n928), .B1(new_n885), .B2(new_n275), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n922), .A2(new_n923), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(KEYINPUT57), .A3(new_n507), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n929), .A2(KEYINPUT113), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n926), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n210), .B(new_n211), .C1(new_n933), .C2(new_n693), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n917), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT115), .ZN(new_n936));
  INV_X1    g735(.A(new_n934), .ZN(new_n937));
  NOR4_X1   g736(.A1(new_n911), .A2(G141gat), .A3(new_n462), .A4(new_n693), .ZN(new_n938));
  OAI21_X1  g737(.A(KEYINPUT58), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT115), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n917), .A2(new_n940), .A3(new_n934), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n936), .A2(new_n939), .A3(new_n941), .ZN(G1344gat));
  NAND3_X1  g741(.A1(new_n926), .A2(new_n932), .A3(new_n667), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT59), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n943), .A2(new_n944), .A3(G148gat), .ZN(new_n945));
  OAI21_X1  g744(.A(KEYINPUT57), .B1(new_n885), .B2(new_n275), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT116), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n512), .A2(new_n947), .A3(new_n697), .A4(new_n463), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n667), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n947), .B1(new_n910), .B2(new_n463), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n930), .A2(new_n507), .A3(new_n928), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n946), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G148gat), .ZN(new_n954));
  AOI21_X1  g753(.A(KEYINPUT117), .B1(new_n954), .B2(KEYINPUT59), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT117), .ZN(new_n956));
  AOI211_X1 g755(.A(new_n956), .B(new_n944), .C1(new_n953), .C2(G148gat), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n945), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n915), .A2(new_n209), .A3(new_n667), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT118), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n958), .A2(KEYINPUT118), .A3(new_n959), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1345gat));
  AOI21_X1  g763(.A(G155gat), .B1(new_n915), .B2(new_n565), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n933), .A2(new_n795), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n965), .B1(new_n966), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g766(.A(G162gat), .B1(new_n915), .B2(new_n720), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n933), .A2(new_n722), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n969), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g769(.A1(new_n697), .A2(new_n463), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT119), .ZN(new_n972));
  NOR4_X1   g771(.A1(new_n972), .A2(new_n885), .A3(new_n507), .A4(new_n810), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g773(.A(G169gat), .B1(new_n974), .B2(new_n693), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n930), .A2(new_n460), .A3(new_n462), .A4(new_n887), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n977), .A2(new_n292), .A3(new_n797), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n975), .A2(new_n978), .ZN(G1348gat));
  NAND3_X1  g778(.A1(new_n973), .A2(G176gat), .A3(new_n717), .ZN(new_n980));
  XOR2_X1   g779(.A(new_n980), .B(KEYINPUT120), .Z(new_n981));
  AOI21_X1  g780(.A(G176gat), .B1(new_n977), .B2(new_n667), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n981), .A2(new_n982), .ZN(G1349gat));
  AOI21_X1  g782(.A(new_n319), .B1(new_n973), .B2(new_n565), .ZN(new_n984));
  NOR3_X1   g783(.A1(new_n976), .A2(new_n316), .A3(new_n795), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g785(.A(new_n986), .B(KEYINPUT60), .Z(G1350gat));
  OAI21_X1  g786(.A(G190gat), .B1(new_n974), .B2(new_n722), .ZN(new_n988));
  OR3_X1    g787(.A1(new_n988), .A2(KEYINPUT122), .A3(KEYINPUT61), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(KEYINPUT61), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(KEYINPUT121), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT121), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n988), .A2(new_n992), .A3(KEYINPUT61), .ZN(new_n993));
  OAI21_X1  g792(.A(KEYINPUT122), .B1(new_n988), .B2(KEYINPUT61), .ZN(new_n994));
  NAND4_X1  g793(.A1(new_n989), .A2(new_n991), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n977), .A2(new_n322), .A3(new_n720), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(G1351gat));
  XNOR2_X1  g796(.A(KEYINPUT123), .B(G197gat), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT124), .ZN(new_n999));
  OR3_X1    g798(.A1(new_n972), .A2(new_n999), .A3(new_n706), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n999), .B1(new_n972), .B2(new_n706), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AND2_X1   g801(.A1(new_n946), .A2(new_n952), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n998), .B1(new_n1004), .B2(new_n693), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n909), .A2(new_n512), .A3(new_n971), .ZN(new_n1006));
  OR2_X1    g805(.A1(new_n693), .A2(new_n998), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(G1352gat));
  OR3_X1    g807(.A1(new_n1004), .A2(KEYINPUT125), .A3(new_n716), .ZN(new_n1009));
  OAI21_X1  g808(.A(KEYINPUT125), .B1(new_n1004), .B2(new_n716), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1009), .A2(G204gat), .A3(new_n1010), .ZN(new_n1011));
  NOR3_X1   g810(.A1(new_n1006), .A2(G204gat), .A3(new_n668), .ZN(new_n1012));
  XNOR2_X1  g811(.A(new_n1012), .B(KEYINPUT62), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1011), .A2(new_n1013), .ZN(G1353gat));
  NAND3_X1  g813(.A1(new_n1002), .A2(new_n565), .A3(new_n1003), .ZN(new_n1015));
  INV_X1    g814(.A(KEYINPUT127), .ZN(new_n1016));
  OR2_X1    g815(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1018));
  NAND3_X1  g817(.A1(new_n1017), .A2(G211gat), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1019), .A2(KEYINPUT63), .ZN(new_n1020));
  INV_X1    g819(.A(KEYINPUT63), .ZN(new_n1021));
  NAND4_X1  g820(.A1(new_n1017), .A2(new_n1021), .A3(G211gat), .A4(new_n1018), .ZN(new_n1022));
  INV_X1    g821(.A(new_n225), .ZN(new_n1023));
  NOR3_X1   g822(.A1(new_n1006), .A2(new_n1023), .A3(new_n795), .ZN(new_n1024));
  XNOR2_X1  g823(.A(new_n1024), .B(KEYINPUT126), .ZN(new_n1025));
  NAND3_X1  g824(.A1(new_n1020), .A2(new_n1022), .A3(new_n1025), .ZN(G1354gat));
  OAI21_X1  g825(.A(G218gat), .B1(new_n1004), .B2(new_n722), .ZN(new_n1027));
  NAND2_X1  g826(.A1(new_n720), .A2(new_n221), .ZN(new_n1028));
  OAI21_X1  g827(.A(new_n1027), .B1(new_n1006), .B2(new_n1028), .ZN(G1355gat));
endmodule


