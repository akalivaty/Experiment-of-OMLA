//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 1 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 1 0 1 0 0 0 0 1 1 1 0 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1313, new_n1314, new_n1315,
    new_n1316, new_n1317, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1372, new_n1373, new_n1374, new_n1375;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT64), .B(G244), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n217), .A2(G77), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G107), .A2(G264), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n208), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XOR2_X1   g0036(.A(G107), .B(G116), .Z(new_n237));
  XOR2_X1   g0037(.A(new_n236), .B(new_n237), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  INV_X1    g0042(.A(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G351));
  NAND3_X1  g0044(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n245), .A2(G50), .ZN(new_n246));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n214), .ZN(new_n248));
  AOI21_X1  g0048(.A(new_n248), .B1(new_n205), .B2(G20), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n246), .B1(new_n249), .B2(G50), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n206), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT69), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n206), .A2(KEYINPUT69), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G58), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(KEYINPUT8), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT68), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n258), .B(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(KEYINPUT8), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n261), .B(KEYINPUT67), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n256), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n264));
  INV_X1    g0064(.A(G150), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n264), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n248), .B1(new_n263), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n251), .B1(new_n269), .B2(KEYINPUT70), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT70), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n271), .B(new_n248), .C1(new_n263), .C2(new_n268), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(KEYINPUT9), .A3(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  OAI21_X1  g0074(.A(KEYINPUT66), .B1(new_n274), .B2(new_n214), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT66), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n276), .A2(new_n277), .A3(G1), .A4(G13), .ZN(new_n278));
  INV_X1    g0078(.A(G41), .ZN(new_n279));
  INV_X1    g0079(.A(G45), .ZN(new_n280));
  AOI21_X1  g0080(.A(G1), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n275), .A2(G274), .A3(new_n278), .A4(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n275), .A2(new_n278), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G226), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT3), .ZN(new_n287));
  INV_X1    g0087(.A(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  AOI21_X1  g0090(.A(G1698), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G222), .ZN(new_n292));
  INV_X1    g0092(.A(G77), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n289), .A2(new_n290), .ZN(new_n294));
  INV_X1    g0094(.A(G1698), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(new_n289), .B2(new_n290), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G223), .ZN(new_n298));
  OAI221_X1 g0098(.A(new_n292), .B1(new_n293), .B2(new_n294), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n276), .A2(G1), .A3(G13), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n286), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G190), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n273), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(KEYINPUT9), .B1(new_n270), .B2(new_n272), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G200), .ZN(new_n307));
  OR2_X1    g0107(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n306), .B(new_n308), .C1(KEYINPUT72), .C2(KEYINPUT10), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n270), .A2(new_n272), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT9), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n312), .A2(new_n308), .A3(new_n273), .A4(new_n303), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n312), .A2(KEYINPUT72), .A3(new_n273), .A4(new_n303), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT10), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n310), .ZN(new_n317));
  INV_X1    g0117(.A(G179), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n302), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(G169), .B2(new_n302), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n309), .A2(new_n316), .A3(new_n321), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n205), .B(G274), .C1(G41), .C2(G45), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n281), .B2(new_n228), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n324), .A2(new_n275), .A3(new_n278), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n298), .A2(new_n295), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n285), .A2(G1698), .ZN(new_n327));
  AND2_X1   g0127(.A1(KEYINPUT3), .A2(G33), .ZN(new_n328));
  NOR2_X1   g0128(.A1(KEYINPUT3), .A2(G33), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n326), .B(new_n327), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G33), .A2(G87), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n300), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n325), .A2(new_n318), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G169), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n330), .A2(new_n331), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n301), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n324), .A2(new_n275), .A3(new_n278), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(KEYINPUT76), .B1(new_n333), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(G169), .B1(new_n325), .B2(new_n332), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT76), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n336), .A2(G179), .A3(new_n337), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n249), .B1(new_n260), .B2(new_n262), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n260), .A2(new_n262), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n345), .B1(new_n347), .B2(new_n245), .ZN(new_n348));
  INV_X1    g0148(.A(new_n248), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n328), .A2(new_n329), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT7), .B1(new_n350), .B2(new_n206), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n289), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n290), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(G68), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G159), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n267), .A2(new_n355), .ZN(new_n356));
  AND2_X1   g0156(.A1(G58), .A2(G68), .ZN(new_n357));
  OAI21_X1  g0157(.A(G20), .B1(new_n357), .B2(new_n201), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT75), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT75), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n360), .B(G20), .C1(new_n357), .C2(new_n201), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n356), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n354), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT16), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n349), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n354), .A2(new_n362), .A3(KEYINPUT16), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n348), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT18), .B1(new_n344), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n356), .ZN(new_n369));
  XNOR2_X1  g0169(.A(G58), .B(G68), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n360), .B1(new_n370), .B2(G20), .ZN(new_n371));
  INV_X1    g0171(.A(new_n361), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G68), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n289), .A2(new_n206), .A3(new_n290), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n374), .B1(new_n377), .B2(new_n352), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n364), .B1(new_n373), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n379), .A2(new_n248), .A3(new_n366), .ZN(new_n380));
  INV_X1    g0180(.A(new_n345), .ZN(new_n381));
  INV_X1    g0181(.A(new_n245), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n381), .B1(new_n346), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n307), .B1(new_n325), .B2(new_n332), .ZN(new_n384));
  INV_X1    g0184(.A(G190), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n336), .A2(new_n385), .A3(new_n337), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n380), .A2(new_n383), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT17), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n367), .A2(KEYINPUT17), .A3(new_n387), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n380), .A2(new_n383), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT18), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n392), .A2(new_n393), .A3(new_n339), .A4(new_n343), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n368), .A2(new_n390), .A3(new_n391), .A4(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G20), .A2(G77), .ZN(new_n396));
  XNOR2_X1  g0196(.A(KEYINPUT15), .B(G87), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT8), .B(G58), .ZN(new_n398));
  OAI221_X1 g0198(.A(new_n396), .B1(new_n397), .B2(new_n252), .C1(new_n267), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n248), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n382), .A2(new_n293), .ZN(new_n401));
  INV_X1    g0201(.A(new_n249), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n400), .B(new_n401), .C1(new_n293), .C2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n294), .A2(G232), .A3(new_n295), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n350), .A2(G107), .ZN(new_n405));
  INV_X1    g0205(.A(G238), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n404), .B(new_n405), .C1(new_n297), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n301), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n275), .A2(new_n217), .A3(new_n278), .A4(new_n283), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n409), .A2(new_n282), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n403), .B(KEYINPUT71), .C1(new_n411), .C2(G169), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT71), .ZN(new_n413));
  AOI21_X1  g0213(.A(G169), .B1(new_n408), .B2(new_n410), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n401), .B1(new_n402), .B2(new_n293), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n248), .B2(new_n399), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n413), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n411), .A2(new_n318), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n412), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n411), .A2(G190), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n420), .B(new_n416), .C1(new_n307), .C2(new_n411), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n395), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n275), .A2(G238), .A3(new_n278), .A4(new_n283), .ZN(new_n424));
  NAND2_X1  g0224(.A1(G33), .A2(G97), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(G226), .A2(G1698), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n228), .B2(G1698), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n426), .B1(new_n428), .B2(new_n294), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n282), .B(new_n424), .C1(new_n429), .C2(new_n300), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT13), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n285), .A2(new_n295), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n228), .A2(G1698), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n432), .B(new_n433), .C1(new_n328), .C2(new_n329), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n301), .B1(new_n435), .B2(new_n426), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT13), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(new_n282), .A4(new_n424), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n431), .A2(new_n438), .A3(KEYINPUT73), .ZN(new_n439));
  OR3_X1    g0239(.A1(new_n430), .A2(KEYINPUT73), .A3(KEYINPUT13), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(new_n440), .A3(G169), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT14), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT14), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n439), .A2(new_n440), .A3(new_n443), .A4(G169), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n431), .A2(new_n438), .A3(G179), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n442), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n254), .A2(G77), .A3(new_n255), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n266), .A2(G50), .B1(G20), .B2(new_n374), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n248), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT11), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(KEYINPUT11), .A3(new_n248), .ZN(new_n453));
  OR3_X1    g0253(.A1(new_n245), .A2(KEYINPUT12), .A3(G68), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT12), .B1(new_n245), .B2(G68), .ZN(new_n455));
  AOI22_X1  g0255(.A1(G68), .A2(new_n249), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n452), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT74), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT74), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n452), .A2(new_n459), .A3(new_n453), .A4(new_n456), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n446), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n439), .A2(new_n440), .A3(G200), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n385), .B1(new_n430), .B2(KEYINPUT13), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n457), .B1(new_n438), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n322), .A2(new_n423), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  OAI211_X1 g0269(.A(G264), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT82), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n294), .A2(KEYINPUT82), .A3(G264), .A4(G1698), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n291), .A2(G257), .B1(new_n350), .B2(G303), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n474), .A2(KEYINPUT83), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT83), .B1(new_n474), .B2(new_n475), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n301), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n280), .A2(G1), .ZN(new_n479));
  AND2_X1   g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  NOR2_X1   g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n482), .A2(new_n275), .A3(G270), .A4(new_n278), .ZN(new_n483));
  XNOR2_X1  g0283(.A(KEYINPUT5), .B(G41), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n205), .A2(G45), .A3(G274), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n275), .A2(new_n484), .A3(new_n486), .A4(new_n278), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n478), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n205), .A2(G33), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n245), .A2(new_n491), .A3(new_n214), .A4(new_n247), .ZN(new_n492));
  INV_X1    g0292(.A(G116), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT80), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT80), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G116), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OAI22_X1  g0297(.A1(new_n492), .A2(new_n493), .B1(new_n245), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n494), .A2(new_n496), .A3(G20), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n248), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT84), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT84), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n500), .A2(new_n503), .A3(new_n248), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G283), .ZN(new_n506));
  INV_X1    g0306(.A(G97), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n506), .B(new_n206), .C1(G33), .C2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT20), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n500), .A2(new_n503), .A3(new_n248), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n503), .B1(new_n500), .B2(new_n248), .ZN(new_n511));
  OAI211_X1 g0311(.A(KEYINPUT20), .B(new_n508), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n499), .B1(new_n509), .B2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n490), .A2(KEYINPUT21), .A3(G169), .A4(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT82), .B1(new_n296), .B2(G264), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n470), .A2(new_n471), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n475), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT83), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n474), .A2(KEYINPUT83), .A3(new_n475), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n488), .B1(new_n522), .B2(new_n301), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(G179), .A3(new_n514), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n515), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g0325(.A(KEYINPUT85), .B(KEYINPUT21), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n508), .B1(new_n510), .B2(new_n511), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT20), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n498), .B1(new_n530), .B2(new_n512), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(new_n334), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n527), .B1(new_n532), .B2(new_n490), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n525), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n514), .B1(new_n490), .B2(G200), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n385), .B2(new_n490), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n349), .A2(KEYINPUT78), .A3(new_n245), .A4(new_n491), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT78), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n492), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n397), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n538), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT19), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n206), .B1(new_n425), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(G87), .ZN(new_n545));
  INV_X1    g0345(.A(G107), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n507), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n206), .B(G68), .C1(new_n328), .C2(new_n329), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n543), .B1(new_n252), .B2(new_n507), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n248), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n397), .A2(new_n382), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n542), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n497), .A2(G33), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n406), .A2(new_n295), .ZN(new_n556));
  INV_X1    g0356(.A(G244), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G1698), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n556), .B(new_n558), .C1(new_n328), .C2(new_n329), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n300), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(G250), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n485), .B1(new_n479), .B2(new_n561), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n562), .A2(new_n275), .A3(new_n278), .ZN(new_n563));
  OAI21_X1  g0363(.A(G169), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n275), .A3(new_n278), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n556), .A2(new_n558), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n566), .A2(new_n294), .B1(new_n497), .B2(G33), .ZN(new_n567));
  OAI211_X1 g0367(.A(G179), .B(new_n565), .C1(new_n567), .C2(new_n300), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n554), .A2(KEYINPUT81), .B1(new_n564), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT81), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n542), .A2(new_n552), .A3(new_n570), .A4(new_n553), .ZN(new_n571));
  OAI21_X1  g0371(.A(G200), .B1(new_n560), .B2(new_n563), .ZN(new_n572));
  OAI211_X1 g0372(.A(G190), .B(new_n565), .C1(new_n567), .C2(new_n300), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n538), .A2(new_n540), .A3(G87), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n575), .A2(new_n552), .A3(new_n553), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n569), .A2(new_n571), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(G250), .A2(G1698), .ZN(new_n579));
  INV_X1    g0379(.A(G257), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n579), .B1(new_n580), .B2(G1698), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n294), .ZN(new_n582));
  NAND2_X1  g0382(.A1(G33), .A2(G294), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n301), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n482), .A2(new_n275), .A3(G264), .A4(new_n278), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n585), .A2(new_n318), .A3(new_n487), .A4(new_n586), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n581), .A2(new_n294), .B1(G33), .B2(G294), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n487), .B(new_n586), .C1(new_n588), .C2(new_n300), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n334), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n206), .B(G87), .C1(new_n328), .C2(new_n329), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT22), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT22), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n294), .A2(new_n594), .A3(new_n206), .A4(G87), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n497), .A2(new_n206), .A3(G33), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT23), .ZN(new_n598));
  OAI211_X1 g0398(.A(G20), .B(new_n546), .C1(new_n598), .C2(KEYINPUT86), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n206), .A2(G107), .ZN(new_n600));
  XNOR2_X1  g0400(.A(KEYINPUT86), .B(KEYINPUT23), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n597), .B(new_n599), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(KEYINPUT24), .B1(new_n596), .B2(new_n602), .ZN(new_n603));
  XNOR2_X1  g0403(.A(KEYINPUT80), .B(G116), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n604), .A2(G20), .A3(new_n288), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n599), .B1(new_n601), .B2(new_n600), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT24), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n593), .A2(new_n595), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n349), .B1(new_n603), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n538), .A2(new_n540), .A3(G107), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n245), .A2(G107), .ZN(new_n613));
  XNOR2_X1  g0413(.A(new_n613), .B(KEYINPUT25), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n591), .B1(new_n611), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(G107), .B1(new_n351), .B2(new_n353), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n507), .A2(new_n546), .A3(KEYINPUT6), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT6), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(G97), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n546), .A2(KEYINPUT77), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT77), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(G107), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n618), .A2(new_n620), .A3(new_n621), .A4(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n618), .A2(new_n620), .B1(new_n621), .B2(new_n623), .ZN(new_n625));
  OAI21_X1  g0425(.A(G20), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n266), .A2(G77), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n617), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n248), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n538), .A2(new_n540), .A3(G97), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n382), .A2(new_n507), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(G244), .B(new_n295), .C1(new_n328), .C2(new_n329), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT4), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n294), .A2(KEYINPUT4), .A3(G244), .A4(new_n295), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n294), .A2(G250), .A3(G1698), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n637), .A2(new_n638), .A3(new_n506), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n301), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n482), .A2(new_n275), .A3(G257), .A4(new_n278), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n487), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n334), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT79), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n642), .A2(new_n487), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n647), .B1(new_n642), .B2(new_n487), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n641), .B(new_n318), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n634), .A2(new_n646), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n632), .B1(new_n628), .B2(new_n248), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n643), .B1(new_n640), .B2(new_n301), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(G190), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n643), .A2(KEYINPUT79), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n656), .A2(new_n648), .B1(new_n301), .B2(new_n640), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n653), .B(new_n655), .C1(new_n657), .C2(new_n307), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n608), .B1(new_n607), .B2(new_n609), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n248), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n589), .A2(new_n307), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(G190), .B2(new_n589), .ZN(new_n663));
  INV_X1    g0463(.A(new_n615), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n661), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n616), .A2(new_n652), .A3(new_n658), .A4(new_n665), .ZN(new_n666));
  NOR4_X1   g0466(.A1(new_n469), .A2(new_n537), .A3(new_n578), .A4(new_n666), .ZN(G372));
  INV_X1    g0467(.A(new_n321), .ZN(new_n668));
  AOI221_X4 g0468(.A(KEYINPUT18), .B1(new_n340), .B2(new_n342), .C1(new_n380), .C2(new_n383), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n340), .A2(new_n342), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n393), .B1(new_n392), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n412), .A2(new_n417), .A3(new_n418), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n446), .A2(new_n461), .B1(new_n673), .B2(new_n466), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n674), .A2(KEYINPUT89), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n388), .B(KEYINPUT17), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n674), .B2(KEYINPUT89), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n672), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n309), .A2(new_n316), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n668), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n634), .A2(new_n646), .A3(new_n651), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n681), .A2(KEYINPUT26), .A3(new_n577), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT26), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n576), .A2(new_n573), .A3(new_n572), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n564), .A2(new_n568), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n554), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n683), .B1(new_n652), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n682), .A2(KEYINPUT88), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT88), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n681), .A2(new_n577), .A3(new_n690), .A4(KEYINPUT26), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n689), .A2(new_n686), .A3(new_n691), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n684), .A2(new_n686), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n693), .A2(new_n652), .A3(new_n658), .A4(new_n665), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n514), .A2(G169), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n526), .B1(new_n695), .B2(new_n523), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n696), .A2(new_n515), .A3(new_n524), .A4(new_n616), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n694), .B1(new_n697), .B2(KEYINPUT87), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n515), .A2(new_n524), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT87), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n699), .A2(new_n700), .A3(new_n696), .A4(new_n616), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n692), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n680), .B1(new_n469), .B2(new_n702), .ZN(G369));
  NAND3_X1  g0503(.A1(new_n696), .A2(new_n515), .A3(new_n524), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(G213), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(G343), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n531), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n704), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n537), .B2(new_n712), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n710), .B1(new_n611), .B2(new_n615), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n616), .A2(new_n717), .A3(new_n665), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n661), .A2(new_n664), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(new_n591), .A3(new_n710), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT90), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT90), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n718), .A2(new_n723), .A3(new_n720), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n716), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n616), .A2(new_n710), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n711), .B1(new_n525), .B2(new_n533), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT91), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT91), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n730), .B(new_n711), .C1(new_n525), .C2(new_n533), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n727), .B1(new_n732), .B2(new_n725), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n726), .A2(new_n733), .ZN(G399));
  INV_X1    g0534(.A(new_n209), .ZN(new_n735));
  OR3_X1    g0535(.A1(new_n735), .A2(KEYINPUT92), .A3(G41), .ZN(new_n736));
  OAI21_X1  g0536(.A(KEYINPUT92), .B1(new_n735), .B2(G41), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n547), .A2(G116), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n739), .A2(new_n205), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n742), .B1(new_n213), .B2(new_n739), .ZN(new_n743));
  XOR2_X1   g0543(.A(new_n743), .B(KEYINPUT28), .Z(new_n744));
  INV_X1    g0544(.A(new_n694), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n697), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n681), .A2(new_n683), .A3(new_n577), .ZN(new_n747));
  OAI21_X1  g0547(.A(KEYINPUT26), .B1(new_n652), .B2(new_n687), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n747), .A2(new_n748), .A3(new_n686), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n710), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(KEYINPUT29), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n698), .A2(new_n701), .ZN(new_n752));
  INV_X1    g0552(.A(new_n692), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n710), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n751), .B1(new_n754), .B2(KEYINPUT29), .ZN(new_n755));
  INV_X1    g0555(.A(G330), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n710), .A2(KEYINPUT31), .ZN(new_n757));
  INV_X1    g0557(.A(new_n568), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n586), .B1(new_n588), .B2(new_n300), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n488), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n758), .A2(new_n654), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n300), .B1(new_n520), .B2(new_n521), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n589), .B(new_n318), .C1(new_n560), .C2(new_n563), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n657), .A2(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n763), .A2(KEYINPUT30), .B1(new_n490), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT30), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(new_n761), .B2(new_n762), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n757), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  OAI211_X1 g0569(.A(KEYINPUT93), .B(new_n767), .C1(new_n761), .C2(new_n762), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT93), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n766), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n710), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT31), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n769), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n666), .A2(new_n578), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n534), .A2(new_n777), .A3(new_n536), .A4(new_n711), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n756), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n755), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n744), .B1(new_n781), .B2(G1), .ZN(G364));
  AND2_X1   g0582(.A1(new_n206), .A2(G13), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n205), .B1(new_n783), .B2(G45), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n739), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G13), .A2(G33), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(G20), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n214), .B1(G20), .B2(new_n334), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT94), .Z(new_n792));
  NAND2_X1  g0592(.A1(new_n209), .A2(new_n294), .ZN(new_n793));
  INV_X1    g0593(.A(G355), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n793), .A2(new_n794), .B1(G116), .B2(new_n209), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n735), .A2(new_n294), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n280), .B2(new_n213), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n243), .A2(G45), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n385), .A2(G20), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT97), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n803), .A2(G179), .A3(new_n307), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n546), .ZN(new_n806));
  NAND2_X1  g0606(.A1(G20), .A2(G179), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT95), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n385), .A2(new_n307), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n806), .B1(G50), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n307), .A2(G179), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n813), .A2(G20), .A3(G190), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n350), .B1(new_n815), .B2(G87), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n385), .A2(G200), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n808), .A2(new_n817), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n812), .B(new_n816), .C1(new_n257), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n808), .A2(new_n385), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(new_n307), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n374), .ZN(new_n823));
  NOR2_X1   g0623(.A1(G179), .A2(G200), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n206), .B1(new_n824), .B2(G190), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT98), .Z(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n507), .ZN(new_n828));
  NOR3_X1   g0628(.A1(new_n803), .A2(G179), .A3(G200), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(G159), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT32), .ZN(new_n831));
  NOR4_X1   g0631(.A1(new_n819), .A2(new_n823), .A3(new_n828), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n820), .A2(G200), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n834), .A2(KEYINPUT96), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n834), .A2(KEYINPUT96), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(G77), .ZN(new_n839));
  INV_X1    g0639(.A(new_n825), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n811), .A2(G326), .B1(G294), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(G311), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n841), .B1(new_n842), .B2(new_n834), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT99), .ZN(new_n844));
  INV_X1    g0644(.A(G283), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n350), .B1(new_n805), .B2(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n814), .B(KEYINPUT100), .ZN(new_n847));
  AOI22_X1  g0647(.A1(G329), .A2(new_n829), .B1(new_n847), .B2(G303), .ZN(new_n848));
  INV_X1    g0648(.A(G322), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n848), .B1(new_n849), .B2(new_n818), .ZN(new_n850));
  XNOR2_X1  g0650(.A(KEYINPUT33), .B(G317), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n846), .B(new_n850), .C1(new_n821), .C2(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n832), .A2(new_n839), .B1(new_n844), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n790), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n786), .B1(new_n792), .B2(new_n800), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT101), .ZN(new_n856));
  INV_X1    g0656(.A(new_n789), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n856), .B1(new_n714), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n716), .A2(new_n786), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(G330), .B2(new_n714), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(G396));
  NAND2_X1  g0662(.A1(new_n403), .A2(new_n710), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n673), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n422), .B2(new_n864), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n419), .A2(new_n421), .A3(new_n711), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n754), .A2(new_n866), .B1(new_n702), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n786), .B1(new_n868), .B2(new_n780), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n780), .B2(new_n868), .ZN(new_n870));
  INV_X1    g0670(.A(new_n786), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n790), .A2(new_n787), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(new_n293), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n818), .ZN(new_n874));
  AOI22_X1  g0674(.A1(G294), .A2(new_n874), .B1(new_n811), .B2(G303), .ZN(new_n875));
  INV_X1    g0675(.A(new_n829), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n875), .B1(new_n545), .B2(new_n805), .C1(new_n842), .C2(new_n876), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n294), .B(new_n828), .C1(G107), .C2(new_n847), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n845), .B2(new_n822), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n877), .B(new_n879), .C1(new_n497), .C2(new_n838), .ZN(new_n880));
  AOI22_X1  g0680(.A1(G137), .A2(new_n811), .B1(new_n874), .B2(G143), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n265), .B2(new_n822), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n838), .B2(G159), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n883), .A2(KEYINPUT34), .ZN(new_n884));
  INV_X1    g0684(.A(G132), .ZN(new_n885));
  OAI221_X1 g0685(.A(new_n294), .B1(new_n825), .B2(new_n257), .C1(new_n876), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n804), .A2(G68), .ZN(new_n887));
  INV_X1    g0687(.A(new_n847), .ZN(new_n888));
  INV_X1    g0688(.A(G50), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT102), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n886), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n891), .B2(new_n890), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n883), .B2(KEYINPUT34), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n880), .B1(new_n884), .B2(new_n894), .ZN(new_n895));
  OAI221_X1 g0695(.A(new_n873), .B1(new_n788), .B2(new_n866), .C1(new_n895), .C2(new_n854), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n870), .A2(new_n896), .ZN(G384));
  NOR2_X1   g0697(.A1(new_n624), .A2(new_n625), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n899), .A2(KEYINPUT35), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(KEYINPUT35), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n900), .A2(G116), .A3(new_n215), .A4(new_n901), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n902), .B(KEYINPUT36), .Z(new_n903));
  OR3_X1    g0703(.A1(new_n212), .A2(new_n293), .A3(new_n357), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n889), .A2(G68), .ZN(new_n905));
  AOI211_X1 g0705(.A(new_n205), .B(G13), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n446), .A2(new_n461), .A3(new_n711), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n708), .B1(new_n380), .B2(new_n383), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n395), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n388), .B1(new_n367), .B2(new_n708), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n380), .A2(new_n383), .B1(new_n340), .B2(new_n342), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT37), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n333), .A2(new_n338), .A3(KEYINPUT76), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n341), .B1(new_n340), .B2(new_n342), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n392), .ZN(new_n918));
  INV_X1    g0718(.A(new_n708), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n392), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT37), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n918), .A2(new_n920), .A3(new_n921), .A4(new_n388), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n914), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n911), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT38), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT104), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n911), .A2(new_n923), .A3(KEYINPUT38), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n924), .A2(KEYINPUT104), .A3(new_n925), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n929), .A2(KEYINPUT39), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n920), .B1(new_n672), .B2(new_n676), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n392), .A2(new_n670), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n933), .A2(new_n920), .A3(new_n388), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT37), .B1(new_n917), .B2(new_n392), .ZN(new_n935));
  AND3_X1   g0735(.A1(new_n380), .A2(new_n383), .A3(new_n387), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n936), .A2(new_n910), .ZN(new_n937));
  AOI22_X1  g0737(.A1(KEYINPUT37), .A2(new_n934), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n925), .B1(new_n932), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT39), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n939), .A2(new_n940), .A3(new_n928), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT105), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n939), .A2(KEYINPUT105), .A3(new_n928), .A4(new_n940), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n909), .B1(new_n931), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n673), .A2(new_n711), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT103), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n702), .B2(new_n867), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n458), .A2(new_n460), .A3(new_n710), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n462), .B2(new_n466), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n463), .A2(new_n465), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n950), .B(new_n953), .C1(new_n446), .C2(new_n461), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n949), .A2(new_n930), .A3(new_n929), .A4(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n672), .A2(new_n919), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n946), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n468), .B(new_n751), .C1(new_n754), .C2(KEYINPUT29), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n960), .A2(new_n680), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n959), .B(new_n961), .Z(new_n962));
  INV_X1    g0762(.A(KEYINPUT40), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n929), .A2(new_n930), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n774), .A2(new_n775), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n773), .A2(KEYINPUT31), .A3(new_n710), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n965), .A2(new_n778), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n955), .A2(new_n967), .A3(new_n866), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n963), .B1(new_n964), .B2(new_n968), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n955), .A2(new_n967), .A3(new_n866), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n963), .B1(new_n939), .B2(new_n928), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n468), .A2(new_n967), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n974), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n975), .A2(G330), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n962), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n205), .B2(new_n783), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n962), .A2(new_n977), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n907), .B1(new_n979), .B2(new_n980), .ZN(G367));
  NOR2_X1   g0781(.A1(new_n576), .A2(new_n711), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n982), .A2(new_n554), .A3(new_n685), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n687), .B2(new_n982), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT43), .Z(new_n985));
  NAND2_X1  g0785(.A1(new_n634), .A2(new_n710), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n652), .A2(new_n658), .A3(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT106), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n681), .A2(new_n710), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n987), .A2(new_n988), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n731), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n730), .B1(new_n704), .B2(new_n711), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n725), .B(new_n992), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(KEYINPUT107), .B1(new_n995), .B2(KEYINPUT42), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n729), .A2(new_n731), .B1(new_n724), .B2(new_n722), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT107), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT42), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .A4(new_n992), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n989), .A2(new_n991), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1002), .A2(new_n719), .A3(new_n591), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n710), .B1(new_n1003), .B2(new_n652), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(KEYINPUT42), .B2(new_n995), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT108), .ZN(new_n1006));
  AND3_X1   g0806(.A1(new_n1001), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1006), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n985), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(KEYINPUT110), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT110), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1011), .B(new_n985), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(KEYINPUT108), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1001), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT109), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1015), .A2(KEYINPUT109), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1013), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n726), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n992), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT111), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1023), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1013), .A2(new_n1022), .A3(new_n1026), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n738), .B(KEYINPUT41), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(KEYINPUT113), .B(KEYINPUT44), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n725), .B1(new_n993), .B2(new_n994), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n727), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n992), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1032), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n992), .B(new_n1031), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n733), .A2(new_n992), .A3(new_n1040), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1024), .B1(new_n1039), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n732), .A2(new_n725), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n716), .A2(new_n1047), .A3(new_n1033), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n715), .B1(new_n1046), .B2(new_n997), .ZN(new_n1049));
  AND4_X1   g0849(.A1(new_n780), .A2(new_n1048), .A3(new_n755), .A4(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1031), .B1(new_n733), .B2(new_n992), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1035), .A2(new_n1036), .A3(new_n1032), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1053), .A2(new_n726), .A3(new_n1043), .A4(new_n1042), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1045), .A2(new_n1050), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT114), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1045), .A2(new_n1050), .A3(new_n1054), .A4(KEYINPUT114), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1030), .B1(new_n1059), .B2(new_n781), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1028), .B(new_n1029), .C1(new_n1060), .C2(new_n785), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n837), .A2(new_n889), .B1(new_n355), .B2(new_n822), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1062), .A2(KEYINPUT116), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1062), .A2(KEYINPUT116), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n804), .A2(G77), .ZN(new_n1065));
  INV_X1    g0865(.A(G143), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1065), .B1(new_n810), .B2(new_n1066), .C1(new_n265), .C2(new_n818), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n826), .A2(G68), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n829), .A2(G137), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n350), .B1(new_n815), .B2(G58), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  NOR4_X1   g0871(.A1(new_n1063), .A2(new_n1064), .A3(new_n1067), .A4(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n805), .A2(new_n507), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(G311), .B2(new_n811), .ZN(new_n1074));
  INV_X1    g0874(.A(G317), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n876), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n837), .A2(new_n845), .ZN(new_n1077));
  INV_X1    g0877(.A(G294), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n822), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n847), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1080));
  XOR2_X1   g0880(.A(KEYINPUT115), .B(KEYINPUT46), .Z(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n814), .B2(new_n604), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n294), .B1(new_n840), .B2(G107), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n874), .A2(G303), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1080), .A2(new_n1082), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  NOR4_X1   g0885(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .A4(new_n1085), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n1072), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT47), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n854), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n1088), .B2(new_n1087), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n796), .A2(new_n234), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n790), .B(new_n789), .C1(new_n735), .C2(new_n541), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n871), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1090), .B(new_n1093), .C1(new_n857), .C2(new_n984), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1061), .A2(new_n1094), .ZN(G387));
  OAI22_X1  g0895(.A1(new_n793), .A2(new_n740), .B1(G107), .B2(new_n209), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n231), .A2(G45), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT117), .ZN(new_n1098));
  AOI211_X1 g0898(.A(G45), .B(new_n741), .C1(G68), .C2(G77), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n398), .A2(G50), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT50), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n797), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1096), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n786), .B1(new_n1103), .B2(new_n792), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G317), .A2(new_n874), .B1(new_n811), .B2(G322), .ZN(new_n1105));
  INV_X1    g0905(.A(G303), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1105), .B1(new_n842), .B2(new_n822), .C1(new_n837), .C2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT48), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n815), .A2(G294), .B1(new_n840), .B2(G283), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT49), .Z(new_n1113));
  AOI21_X1  g0913(.A(new_n294), .B1(new_n829), .B2(G326), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n604), .B2(new_n805), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G50), .A2(new_n874), .B1(new_n811), .B2(G159), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n265), .B2(new_n876), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n814), .A2(new_n293), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n1073), .A2(new_n350), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n826), .A2(new_n541), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(G68), .A2(new_n833), .B1(new_n821), .B2(new_n346), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1113), .A2(new_n1115), .B1(new_n1117), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1104), .B1(new_n1123), .B2(new_n790), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n722), .A2(new_n724), .A3(new_n789), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1124), .A2(new_n1125), .B1(new_n1126), .B2(new_n785), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1050), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n739), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1126), .A2(new_n781), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1127), .B1(new_n1129), .B2(new_n1130), .ZN(G393));
  NAND3_X1  g0931(.A1(new_n1045), .A2(new_n785), .A3(new_n1054), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n791), .B1(new_n507), .B2(new_n209), .C1(new_n797), .C2(new_n238), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n786), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n827), .A2(new_n293), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n350), .B1(new_n815), .B2(G68), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1136), .B1(new_n876), .B2(new_n1066), .C1(new_n545), .C2(new_n805), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1135), .B(new_n1137), .C1(G50), .C2(new_n821), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n265), .A2(new_n810), .B1(new_n818), .B2(new_n355), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT51), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1138), .B(new_n1140), .C1(new_n398), .C2(new_n837), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n350), .B1(new_n825), .B2(new_n604), .C1(new_n845), .C2(new_n814), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1142), .B(new_n806), .C1(G322), .C2(new_n829), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n842), .A2(new_n818), .B1(new_n810), .B2(new_n1075), .ZN(new_n1144));
  XOR2_X1   g0944(.A(KEYINPUT118), .B(KEYINPUT52), .Z(new_n1145));
  XNOR2_X1  g0945(.A(new_n1144), .B(new_n1145), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G294), .A2(new_n833), .B1(new_n821), .B2(G303), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1143), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1141), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1134), .B1(new_n1149), .B2(new_n790), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n992), .B2(new_n857), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1132), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT119), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1045), .A2(new_n1054), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n738), .B1(new_n1155), .B2(new_n1128), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1059), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1154), .B1(new_n1059), .B2(new_n1156), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1153), .B1(new_n1157), .B2(new_n1158), .ZN(G390));
  INV_X1    g0959(.A(KEYINPUT121), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n952), .A2(new_n954), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n746), .A2(new_n749), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1162), .A2(new_n711), .A3(new_n866), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1161), .B1(new_n1163), .B2(new_n948), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n939), .A2(new_n928), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n909), .A2(KEYINPUT120), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT120), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n908), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1165), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1160), .B1(new_n1164), .B2(new_n1170), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n939), .A2(new_n928), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT103), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n947), .B(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n750), .B2(new_n866), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1172), .B(KEYINPUT121), .C1(new_n1175), .C2(new_n1161), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1171), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n779), .A2(new_n866), .A3(new_n955), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n944), .B(new_n943), .C1(new_n964), .C2(new_n940), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n909), .B1(new_n949), .B2(new_n955), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1177), .B(new_n1178), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n931), .A2(new_n945), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n949), .A2(new_n955), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n908), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1182), .A2(new_n1184), .B1(new_n1171), .B2(new_n1176), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n967), .A2(G330), .A3(new_n866), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1186), .A2(new_n1161), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1181), .B(new_n785), .C1(new_n1185), .C2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n815), .A2(G150), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n294), .B1(new_n1190), .B2(KEYINPUT53), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n829), .A2(G125), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n805), .B2(new_n889), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1191), .B(new_n1193), .C1(KEYINPUT53), .C2(new_n1190), .ZN(new_n1194));
  XOR2_X1   g0994(.A(KEYINPUT54), .B(G143), .Z(new_n1195));
  NAND2_X1  g0995(.A1(new_n838), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(G128), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n1197), .A2(new_n810), .B1(new_n818), .B2(new_n885), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT123), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G159), .A2(new_n826), .B1(new_n821), .B2(G137), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1194), .A2(new_n1196), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n887), .A2(new_n350), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1202), .B(new_n1135), .C1(G107), .C2(new_n821), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n876), .A2(new_n1078), .B1(new_n845), .B2(new_n810), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n888), .A2(new_n545), .B1(new_n818), .B2(new_n493), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1203), .B(new_n1206), .C1(new_n507), .C2(new_n837), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n854), .B1(new_n1201), .B2(new_n1207), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n871), .B(new_n1208), .C1(new_n347), .C2(new_n872), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1179), .B2(new_n788), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1189), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n468), .A2(G330), .A3(new_n967), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n960), .A2(new_n680), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n955), .B1(new_n779), .B2(new_n866), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n949), .B1(new_n1187), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1186), .A2(new_n1161), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1217), .A2(new_n1175), .A3(new_n1178), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1214), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1181), .B(new_n1219), .C1(new_n1185), .C2(new_n1188), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1220), .A2(KEYINPUT122), .A3(new_n739), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1181), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1219), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1221), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(KEYINPUT122), .B1(new_n1220), .B2(new_n739), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1212), .B1(new_n1225), .B2(new_n1226), .ZN(G378));
  AOI21_X1  g1027(.A(new_n756), .B1(new_n970), .B2(new_n971), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1228), .A2(new_n969), .A3(KEYINPUT124), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n317), .A2(new_n708), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n322), .B(new_n1230), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1231), .B(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1229), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT124), .B1(new_n1228), .B2(new_n969), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n959), .A2(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n959), .A2(new_n1235), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1234), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n957), .B1(new_n1179), .B2(new_n909), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1228), .A2(new_n969), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1239), .B(new_n956), .C1(new_n1240), .C2(KEYINPUT124), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1234), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n959), .A2(new_n1235), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1238), .A2(new_n785), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1233), .A2(new_n787), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n810), .A2(new_n493), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n805), .A2(new_n257), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1247), .B(new_n1248), .C1(G283), .C2(new_n829), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n350), .A2(new_n279), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1118), .B(new_n1250), .C1(new_n874), .C2(G107), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(G97), .A2(new_n821), .B1(new_n833), .B2(new_n541), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1249), .A2(new_n1068), .A3(new_n1251), .A4(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT58), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(G33), .A2(G41), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1255), .A2(G50), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1253), .A2(new_n1254), .B1(new_n1250), .B2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1255), .B1(new_n805), .B2(new_n355), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(G124), .B2(new_n829), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n811), .A2(G125), .B1(new_n815), .B2(new_n1195), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n1197), .B2(new_n818), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n827), .A2(new_n265), .B1(new_n822), .B2(new_n885), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n1261), .B(new_n1262), .C1(G137), .C2(new_n833), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT59), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1259), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1263), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1266), .A2(KEYINPUT59), .ZN(new_n1267));
  OAI221_X1 g1067(.A(new_n1257), .B1(new_n1254), .B2(new_n1253), .C1(new_n1265), .C2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n790), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n872), .A2(new_n889), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1246), .A2(new_n786), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1245), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1214), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1220), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1238), .A2(new_n1244), .A3(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT57), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1238), .A2(new_n1274), .A3(KEYINPUT57), .A4(new_n1244), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n739), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1272), .B1(new_n1277), .B2(new_n1279), .ZN(G375));
  NAND2_X1  g1080(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n785), .ZN(new_n1282));
  AOI211_X1 g1082(.A(new_n350), .B(new_n1248), .C1(new_n821), .C2(new_n1195), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(G132), .A2(new_n811), .B1(new_n874), .B2(G137), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(G128), .A2(new_n829), .B1(new_n847), .B2(G159), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(G50), .A2(new_n826), .B1(new_n833), .B2(G150), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .A4(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1120), .A2(new_n1065), .A3(new_n350), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(new_n497), .B2(new_n821), .ZN(new_n1289));
  OAI22_X1  g1089(.A1(new_n876), .A2(new_n1106), .B1(new_n1078), .B2(new_n810), .ZN(new_n1290));
  OAI22_X1  g1090(.A1(new_n888), .A2(new_n507), .B1(new_n818), .B2(new_n845), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1289), .B(new_n1292), .C1(new_n546), .C2(new_n837), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n854), .B1(new_n1287), .B2(new_n1293), .ZN(new_n1294));
  AOI211_X1 g1094(.A(new_n871), .B(new_n1294), .C1(new_n374), .C2(new_n872), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1295), .B1(new_n955), .B2(new_n788), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1282), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1030), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1223), .A2(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1281), .A2(new_n1273), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1298), .B1(new_n1300), .B2(new_n1301), .ZN(G381));
  NAND2_X1  g1102(.A1(new_n1245), .A2(new_n1271), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1279), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1303), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1221), .A2(new_n1224), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1226), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1211), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1306), .A2(new_n1309), .ZN(new_n1310));
  OR4_X1    g1110(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1311));
  OR4_X1    g1111(.A1(G387), .A2(new_n1310), .A3(G390), .A4(new_n1311), .ZN(G407));
  NOR2_X1   g1112(.A1(G375), .A2(G378), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n709), .A2(G213), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1316));
  XNOR2_X1  g1116(.A(new_n1316), .B(KEYINPUT125), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1317), .A2(G213), .A3(G407), .ZN(G409));
  XNOR2_X1  g1118(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1238), .A2(new_n1274), .A3(new_n1299), .A4(new_n1244), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1320), .A2(new_n1245), .A3(new_n1271), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1315), .B1(new_n1321), .B2(new_n1309), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1322), .B1(new_n1306), .B2(new_n1309), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1301), .B1(KEYINPUT60), .B2(new_n1223), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1216), .A2(new_n1214), .A3(KEYINPUT60), .A4(new_n1218), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n739), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1298), .B1(new_n1324), .B2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(G384), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  OAI211_X1 g1129(.A(G384), .B(new_n1298), .C1(new_n1324), .C2(new_n1326), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1315), .A2(KEYINPUT126), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1329), .A2(new_n1330), .A3(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1315), .A2(G2897), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1333), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1329), .A2(new_n1330), .A3(new_n1335), .A4(new_n1331), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1334), .A2(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1319), .B1(new_n1323), .B2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(G375), .A2(G378), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1339), .A2(new_n1322), .A3(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(KEYINPUT62), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1320), .A2(new_n1245), .A3(new_n1271), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1314), .B1(new_n1344), .B2(G378), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1345), .B1(G378), .B2(G375), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT62), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1346), .A2(new_n1347), .A3(new_n1341), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1338), .A2(new_n1343), .A3(new_n1348), .ZN(new_n1349));
  XNOR2_X1  g1149(.A(G393), .B(new_n861), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1350), .ZN(new_n1351));
  AND3_X1   g1151(.A1(new_n1061), .A2(G390), .A3(new_n1094), .ZN(new_n1352));
  AOI21_X1  g1152(.A(G390), .B1(new_n1094), .B2(new_n1061), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1351), .B1(new_n1352), .B2(new_n1353), .ZN(new_n1354));
  INV_X1    g1154(.A(G390), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(G387), .A2(new_n1355), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1061), .A2(G390), .A3(new_n1094), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1356), .A2(new_n1350), .A3(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1354), .A2(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1349), .A2(new_n1359), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT61), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1305), .A2(new_n739), .A3(new_n1278), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1309), .B1(new_n1362), .B2(new_n1272), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1337), .B1(new_n1363), .B2(new_n1345), .ZN(new_n1364));
  AND4_X1   g1164(.A1(new_n1361), .A2(new_n1354), .A3(new_n1364), .A4(new_n1358), .ZN(new_n1365));
  AOI21_X1  g1165(.A(KEYINPUT63), .B1(new_n1346), .B2(new_n1341), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT63), .ZN(new_n1367));
  NOR4_X1   g1167(.A1(new_n1363), .A2(new_n1345), .A3(new_n1367), .A4(new_n1340), .ZN(new_n1368));
  NOR2_X1   g1168(.A1(new_n1366), .A2(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1365), .A2(new_n1369), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1360), .A2(new_n1370), .ZN(G405));
  INV_X1    g1171(.A(new_n1359), .ZN(new_n1372));
  OAI21_X1  g1172(.A(new_n1341), .B1(new_n1313), .B2(new_n1363), .ZN(new_n1373));
  NAND3_X1  g1173(.A1(new_n1310), .A2(new_n1339), .A3(new_n1340), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1373), .A2(new_n1374), .ZN(new_n1375));
  XNOR2_X1  g1175(.A(new_n1372), .B(new_n1375), .ZN(G402));
endmodule


