//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n999, new_n1000;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n204), .A2(KEYINPUT92), .A3(KEYINPUT16), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT92), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(G1gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n202), .A2(new_n205), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT95), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT95), .ZN(new_n211));
  NAND4_X1  g010(.A1(new_n202), .A2(new_n211), .A3(new_n205), .A4(new_n208), .ZN(new_n212));
  AOI21_X1  g011(.A(G8gat), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G8gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n214), .A2(KEYINPUT94), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n203), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT93), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n209), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT94), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(new_n203), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n209), .A2(new_n217), .ZN(new_n221));
  OAI21_X1  g020(.A(G8gat), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT96), .B1(new_n216), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT90), .B(G29gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G36gat), .ZN(new_n226));
  OR3_X1    g025(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(G43gat), .B(G50gat), .Z(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT91), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT15), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT15), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(KEYINPUT91), .A3(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n230), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT89), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n227), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n228), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n227), .B1(new_n239), .B2(new_n237), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n238), .A2(new_n240), .B1(G36gat), .B2(new_n225), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n231), .A2(new_n234), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n236), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n216), .A2(new_n222), .A3(KEYINPUT96), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n224), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n238), .A2(new_n240), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(new_n226), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n242), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT17), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n250), .A3(new_n236), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n250), .B1(new_n249), .B2(new_n236), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n216), .B(new_n222), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(G229gat), .A2(G233gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n246), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT18), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n256), .A2(KEYINPUT97), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT97), .B1(new_n256), .B2(new_n257), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n255), .B(KEYINPUT13), .Z(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n244), .ZN(new_n264));
  INV_X1    g063(.A(new_n245), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n264), .B1(new_n265), .B2(new_n223), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n263), .B1(new_n246), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G113gat), .B(G141gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(G169gat), .B(G197gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT12), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n268), .B(new_n274), .C1(new_n257), .C2(new_n256), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n261), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n256), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n267), .B1(new_n277), .B2(KEYINPUT18), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n256), .A2(new_n257), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n274), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n282));
  INV_X1    g081(.A(G120gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n282), .B1(new_n283), .B2(G113gat), .ZN(new_n284));
  INV_X1    g083(.A(G113gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(KEYINPUT71), .A3(G120gat), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n284), .B(new_n286), .C1(new_n285), .C2(G120gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n288));
  INV_X1    g087(.A(G127gat), .ZN(new_n289));
  AND2_X1   g088(.A1(new_n289), .A2(G134gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(G134gat), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n288), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G127gat), .B(G134gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT72), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT1), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n287), .A2(new_n292), .A3(new_n294), .A4(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n293), .A2(KEYINPUT70), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n285), .A2(G120gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n283), .A2(G113gat), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n295), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n290), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n297), .B(new_n300), .C1(KEYINPUT70), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT66), .ZN(new_n305));
  NOR2_X1   g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT23), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT23), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n308), .B1(G169gat), .B2(G176gat), .ZN(new_n309));
  OAI211_X1 g108(.A(KEYINPUT25), .B(new_n307), .C1(new_n309), .C2(new_n306), .ZN(new_n310));
  INV_X1    g109(.A(G183gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT64), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT64), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G183gat), .ZN(new_n314));
  INV_X1    g113(.A(G190gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n312), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT24), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT24), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n319), .A2(G183gat), .A3(G190gat), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n316), .A2(KEYINPUT65), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT65), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n312), .A2(new_n314), .A3(new_n322), .A4(new_n315), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n310), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n318), .A2(new_n320), .B1(new_n311), .B2(new_n315), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n308), .A2(G169gat), .A3(G176gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n306), .ZN(new_n328));
  INV_X1    g127(.A(G169gat), .ZN(new_n329));
  INV_X1    g128(.A(G176gat), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT23), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n327), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT25), .B1(new_n326), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n305), .B1(new_n324), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n316), .A2(KEYINPUT65), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(new_n336), .A3(new_n323), .ZN(new_n337));
  INV_X1    g136(.A(new_n310), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT25), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n307), .B1(new_n309), .B2(new_n306), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n340), .B1(new_n341), .B2(new_n325), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n339), .A2(KEYINPUT66), .A3(new_n342), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n334), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT69), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n345), .B1(new_n346), .B2(new_n306), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT26), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n306), .A2(new_n348), .ZN(new_n349));
  MUX2_X1   g148(.A(new_n345), .B(new_n347), .S(new_n349), .Z(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n317), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n312), .A2(new_n314), .A3(KEYINPUT27), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT67), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n312), .A2(new_n314), .A3(KEYINPUT67), .A4(KEYINPUT27), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n315), .B1(new_n311), .B2(KEYINPUT27), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n354), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT68), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT28), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n354), .A2(KEYINPUT68), .A3(new_n355), .A4(new_n357), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT27), .B(G183gat), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(KEYINPUT28), .A3(new_n315), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n351), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n304), .B1(new_n344), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(G227gat), .ZN(new_n368));
  INV_X1    g167(.A(G233gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n362), .A2(new_n361), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n356), .B1(new_n352), .B2(new_n353), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT68), .B1(new_n372), .B2(new_n355), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n365), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n351), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n334), .A2(new_n343), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n303), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n367), .A2(new_n370), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT73), .B1(new_n379), .B2(KEYINPUT32), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(KEYINPUT73), .A3(KEYINPUT32), .ZN(new_n382));
  XNOR2_X1  g181(.A(G15gat), .B(G43gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(G71gat), .B(G99gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT33), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n385), .B1(new_n379), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n381), .A2(new_n382), .A3(new_n387), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n379), .B(KEYINPUT32), .C1(new_n386), .C2(new_n385), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT34), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n367), .A2(new_n378), .ZN(new_n391));
  INV_X1    g190(.A(new_n370), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AOI211_X1 g192(.A(KEYINPUT34), .B(new_n370), .C1(new_n367), .C2(new_n378), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n388), .A2(new_n389), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n387), .A2(new_n382), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n389), .B1(new_n397), .B2(new_n380), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT74), .B1(new_n393), .B2(new_n394), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n376), .A2(new_n303), .A3(new_n377), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n303), .B1(new_n376), .B2(new_n377), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n392), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT34), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT74), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n391), .A2(new_n390), .A3(new_n392), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n399), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT75), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n398), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n408), .B1(new_n398), .B2(new_n407), .ZN(new_n410));
  OAI211_X1 g209(.A(KEYINPUT36), .B(new_n396), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  XOR2_X1   g210(.A(KEYINPUT76), .B(KEYINPUT36), .Z(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n396), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n395), .B1(new_n388), .B2(new_n389), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(G225gat), .A2(G233gat), .ZN(new_n417));
  XOR2_X1   g216(.A(G155gat), .B(G162gat), .Z(new_n418));
  XNOR2_X1  g217(.A(G141gat), .B(G148gat), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n418), .B1(KEYINPUT2), .B2(new_n419), .ZN(new_n420));
  XOR2_X1   g219(.A(G141gat), .B(G148gat), .Z(new_n421));
  XNOR2_X1  g220(.A(G155gat), .B(G162gat), .ZN(new_n422));
  INV_X1    g221(.A(G155gat), .ZN(new_n423));
  INV_X1    g222(.A(G162gat), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT2), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n421), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n296), .A2(new_n302), .A3(new_n420), .A4(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT4), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n420), .A2(new_n426), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT3), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT3), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n420), .A2(new_n426), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n431), .A2(new_n303), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n430), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n435), .A2(KEYINPUT4), .A3(new_n302), .A4(new_n296), .ZN(new_n436));
  AND4_X1   g235(.A1(new_n417), .A2(new_n429), .A3(new_n434), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(KEYINPUT81), .A2(KEYINPUT5), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n303), .A2(new_n430), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n427), .ZN(new_n441));
  INV_X1    g240(.A(new_n417), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n442), .A2(KEYINPUT5), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n437), .A2(new_n439), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G1gat), .B(G29gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n445), .B(KEYINPUT0), .ZN(new_n446));
  XNOR2_X1  g245(.A(G57gat), .B(G85gat), .ZN(new_n447));
  XOR2_X1   g246(.A(new_n446), .B(new_n447), .Z(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n429), .A2(new_n434), .A3(new_n436), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n438), .B1(new_n450), .B2(new_n442), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n444), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT6), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n444), .A2(new_n451), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT6), .B1(new_n455), .B2(new_n448), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT82), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n452), .B1(new_n456), .B2(new_n457), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n454), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(G226gat), .A2(G233gat), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n376), .A2(new_n462), .A3(new_n377), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n324), .A2(new_n333), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n464), .B1(new_n374), .B2(new_n375), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n462), .A2(KEYINPUT29), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(G197gat), .B(G204gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT22), .ZN(new_n469));
  XNOR2_X1  g268(.A(G211gat), .B(G218gat), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT22), .ZN(new_n473));
  INV_X1    g272(.A(G211gat), .ZN(new_n474));
  INV_X1    g273(.A(G218gat), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n470), .A2(new_n468), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n467), .A2(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(G8gat), .B(G36gat), .Z(new_n480));
  XNOR2_X1  g279(.A(new_n480), .B(KEYINPUT79), .ZN(new_n481));
  XOR2_X1   g280(.A(G64gat), .B(G92gat), .Z(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT78), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n465), .B2(new_n461), .ZN(new_n485));
  OAI211_X1 g284(.A(KEYINPUT78), .B(new_n462), .C1(new_n366), .C2(new_n464), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT77), .B(KEYINPUT29), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(new_n344), .B2(new_n366), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n485), .A2(new_n486), .B1(new_n489), .B2(new_n461), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n479), .B(new_n483), .C1(new_n490), .C2(new_n478), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT80), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT30), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n491), .A2(new_n492), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n479), .B1(new_n490), .B2(new_n478), .ZN(new_n496));
  INV_X1    g295(.A(new_n483), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n495), .A2(KEYINPUT30), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n460), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT85), .ZN(new_n500));
  INV_X1    g299(.A(G22gat), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n432), .B1(new_n420), .B2(new_n426), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n477), .A2(KEYINPUT83), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT83), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n470), .A2(new_n468), .A3(new_n504), .A4(new_n476), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n472), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n487), .B1(new_n420), .B2(new_n426), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n508), .A2(KEYINPUT84), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n478), .B1(new_n433), .B2(new_n488), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n510), .B1(new_n508), .B2(KEYINPUT84), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n509), .A2(new_n511), .B1(G228gat), .B2(G233gat), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n478), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n432), .B1(new_n514), .B2(KEYINPUT29), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n430), .ZN(new_n516));
  INV_X1    g315(.A(new_n510), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n516), .A2(G228gat), .A3(G233gat), .A4(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n501), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n518), .ZN(new_n520));
  NOR3_X1   g319(.A1(new_n512), .A2(new_n520), .A3(G22gat), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n500), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G78gat), .B(G106gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT31), .B(G50gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n513), .A2(new_n501), .A3(new_n518), .ZN(new_n527));
  OAI21_X1  g326(.A(G22gat), .B1(new_n512), .B2(new_n520), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT85), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n522), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n500), .B(new_n525), .C1(new_n519), .C2(new_n521), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n411), .A2(new_n416), .B1(new_n499), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT86), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n534), .B1(new_n444), .B2(new_n451), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n420), .A2(new_n426), .A3(new_n432), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n536), .A2(new_n502), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n537), .A2(new_n303), .B1(new_n428), .B2(new_n427), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n538), .A2(new_n417), .A3(new_n436), .A4(new_n439), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n441), .A2(new_n443), .ZN(new_n540));
  AND4_X1   g339(.A1(new_n534), .A2(new_n451), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n449), .B1(new_n535), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n542), .A2(new_n456), .B1(KEYINPUT6), .B2(new_n453), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT37), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n544), .B(new_n479), .C1(new_n490), .C2(new_n478), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n544), .B1(new_n467), .B2(new_n514), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n546), .B1(new_n490), .B2(new_n514), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT38), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n545), .A2(new_n547), .A3(new_n548), .A4(new_n497), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n543), .A2(new_n549), .A3(new_n491), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n496), .A2(KEYINPUT37), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n545), .A2(new_n497), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT38), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n532), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n450), .A2(new_n442), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n555), .B(KEYINPUT39), .C1(new_n442), .C2(new_n441), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n556), .B(new_n448), .C1(KEYINPUT39), .C2(new_n555), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT40), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n558), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n559), .A2(new_n542), .A3(new_n560), .ZN(new_n561));
  AOI211_X1 g360(.A(KEYINPUT87), .B(new_n561), .C1(new_n498), .C2(new_n494), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT87), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n495), .A2(KEYINPUT30), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n496), .A2(new_n497), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n564), .A2(new_n494), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n561), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n563), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n554), .B1(new_n562), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n533), .A2(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n530), .A2(new_n531), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n396), .B(new_n571), .C1(new_n409), .C2(new_n410), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT35), .B1(new_n572), .B2(new_n499), .ZN(new_n573));
  NOR3_X1   g372(.A1(new_n532), .A2(KEYINPUT35), .A3(new_n543), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n414), .A2(new_n415), .ZN(new_n575));
  INV_X1    g374(.A(new_n566), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n281), .B1(new_n570), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G183gat), .B(G211gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT102), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT99), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G57gat), .B(G64gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(G71gat), .ZN(new_n589));
  INV_X1    g388(.A(G78gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n591), .A2(KEYINPUT98), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(KEYINPUT98), .ZN(new_n593));
  AOI22_X1  g392(.A1(new_n592), .A2(new_n593), .B1(G71gat), .B2(G78gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n586), .A2(KEYINPUT100), .ZN(new_n596));
  XNOR2_X1  g395(.A(G71gat), .B(G78gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n586), .A2(KEYINPUT100), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n596), .A2(new_n585), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT21), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G127gat), .B(G155gat), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n609), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n606), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  OAI22_X1  g412(.A1(new_n265), .A2(new_n223), .B1(new_n601), .B2(new_n600), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT101), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n613), .A2(new_n615), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n582), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n618), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n620), .A2(new_n616), .A3(new_n581), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G232gat), .A2(G233gat), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n625), .A2(KEYINPUT41), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT103), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G99gat), .A2(G106gat), .ZN(new_n629));
  INV_X1    g428(.A(G85gat), .ZN(new_n630));
  INV_X1    g429(.A(G92gat), .ZN(new_n631));
  AOI22_X1  g430(.A1(KEYINPUT8), .A2(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT7), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n630), .B2(new_n631), .ZN(new_n634));
  NAND3_X1  g433(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n632), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(G99gat), .B(G106gat), .Z(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT104), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n636), .A2(KEYINPUT104), .A3(new_n637), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n636), .A2(new_n637), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n643), .B1(new_n252), .B2(new_n253), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n244), .A2(new_n645), .B1(KEYINPUT41), .B2(new_n625), .ZN(new_n646));
  XNOR2_X1  g445(.A(G190gat), .B(G218gat), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n644), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n244), .A2(KEYINPUT17), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n645), .B1(new_n650), .B2(new_n251), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n625), .A2(KEYINPUT41), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n652), .B1(new_n264), .B2(new_n643), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n647), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(G134gat), .B(G162gat), .Z(new_n655));
  AND3_X1   g454(.A1(new_n649), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n655), .B1(new_n649), .B2(new_n654), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n628), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n655), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n648), .B1(new_n644), .B2(new_n646), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n651), .A2(new_n653), .A3(new_n647), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n649), .A2(new_n654), .A3(new_n655), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n662), .A2(new_n627), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT105), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n643), .A2(new_n600), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT10), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n595), .A2(new_n599), .A3(new_n638), .A4(new_n642), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n645), .A2(KEYINPUT10), .A3(new_n595), .A4(new_n599), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(G230gat), .A2(G233gat), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n666), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n673), .ZN(new_n675));
  AOI211_X1 g474(.A(KEYINPUT105), .B(new_n675), .C1(new_n670), .C2(new_n671), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n673), .B1(new_n667), .B2(new_n669), .ZN(new_n678));
  XNOR2_X1  g477(.A(G120gat), .B(G148gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(G176gat), .B(G204gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n672), .A2(new_n673), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n681), .B1(new_n685), .B2(new_n678), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n579), .A2(new_n623), .A3(new_n665), .A4(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(new_n460), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(new_n204), .ZN(G1324gat));
  NOR2_X1   g490(.A1(new_n689), .A2(new_n576), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT42), .B1(new_n692), .B2(new_n214), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT16), .B(G8gat), .Z(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  MUX2_X1   g494(.A(KEYINPUT42), .B(new_n693), .S(new_n695), .Z(G1325gat));
  NAND2_X1  g495(.A1(new_n411), .A2(new_n416), .ZN(new_n697));
  OAI21_X1  g496(.A(G15gat), .B1(new_n689), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n575), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n699), .A2(G15gat), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n689), .B2(new_n700), .ZN(G1326gat));
  NOR2_X1   g500(.A1(new_n689), .A2(new_n571), .ZN(new_n702));
  XOR2_X1   g501(.A(KEYINPUT43), .B(G22gat), .Z(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1327gat));
  NOR3_X1   g503(.A1(new_n623), .A2(new_n665), .A3(new_n687), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n579), .A2(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n706), .A2(new_n460), .A3(new_n225), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT45), .Z(new_n708));
  XNOR2_X1  g507(.A(new_n687), .B(KEYINPUT106), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n623), .A2(new_n281), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n570), .A2(new_n578), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT107), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n570), .A2(new_n578), .A3(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n665), .A2(KEYINPUT44), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n714), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n658), .A2(new_n664), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n713), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT44), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n712), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n225), .B1(new_n723), .B2(new_n460), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n724), .ZN(G1328gat));
  OAI21_X1  g524(.A(G36gat), .B1(new_n723), .B2(new_n576), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n706), .A2(G36gat), .A3(new_n576), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT46), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(G1329gat));
  INV_X1    g528(.A(new_n697), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n722), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(G43gat), .ZN(new_n732));
  OAI21_X1  g531(.A(KEYINPUT108), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n579), .A2(new_n732), .A3(new_n575), .A4(new_n705), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(new_n731), .B2(new_n732), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n733), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  OAI221_X1 g536(.A(new_n734), .B1(KEYINPUT108), .B2(KEYINPUT47), .C1(new_n731), .C2(new_n732), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(G1330gat));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n706), .A2(G50gat), .A3(new_n571), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n570), .A2(new_n578), .A3(new_n715), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n715), .B1(new_n570), .B2(new_n578), .ZN(new_n743));
  INV_X1    g542(.A(new_n717), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n665), .B1(new_n570), .B2(new_n578), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n532), .B(new_n711), .C1(new_n745), .C2(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n741), .B1(new_n749), .B2(G50gat), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n740), .B1(new_n750), .B2(KEYINPUT48), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT48), .ZN(new_n752));
  INV_X1    g551(.A(G50gat), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n753), .B1(new_n722), .B2(new_n532), .ZN(new_n754));
  OAI211_X1 g553(.A(KEYINPUT109), .B(new_n752), .C1(new_n754), .C2(new_n741), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n749), .A2(KEYINPUT110), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n758), .B1(new_n722), .B2(new_n532), .ZN(new_n759));
  OAI21_X1  g558(.A(G50gat), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n741), .A2(new_n752), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n756), .A2(new_n762), .ZN(G1331gat));
  NOR2_X1   g562(.A1(new_n742), .A2(new_n743), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n619), .A2(new_n621), .A3(new_n665), .ZN(new_n765));
  INV_X1    g564(.A(new_n281), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n765), .A2(new_n766), .A3(new_n709), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n460), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g571(.A(new_n576), .B(new_n768), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n773));
  NOR2_X1   g572(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1333gat));
  OAI21_X1  g574(.A(G71gat), .B1(new_n768), .B2(new_n697), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n575), .A2(new_n589), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n768), .B2(new_n777), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n778), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g578(.A1(new_n768), .A2(new_n571), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(new_n590), .ZN(G1335gat));
  NOR2_X1   g580(.A1(new_n623), .A2(new_n766), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n783), .A2(new_n688), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(new_n718), .B2(new_n721), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(G85gat), .B1(new_n787), .B2(new_n460), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n746), .A2(KEYINPUT51), .A3(new_n782), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT51), .B1(new_n746), .B2(new_n782), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n790), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n794), .A2(KEYINPUT112), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT112), .B1(new_n794), .B2(new_n795), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n687), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n770), .A2(new_n630), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n788), .B1(new_n798), .B2(new_n799), .ZN(G1336gat));
  NAND2_X1  g599(.A1(new_n794), .A2(new_n795), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n576), .A2(new_n709), .A3(G92gat), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT52), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n786), .A2(new_n804), .A3(new_n566), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(G92gat), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n804), .B1(new_n786), .B2(new_n566), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n803), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n631), .B1(new_n786), .B2(new_n566), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n746), .A2(KEYINPUT113), .A3(new_n782), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT51), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(KEYINPUT51), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n746), .A2(new_n782), .B1(KEYINPUT113), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n809), .B1(new_n802), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n808), .B1(new_n816), .B2(new_n817), .ZN(G1337gat));
  OAI21_X1  g617(.A(G99gat), .B1(new_n787), .B2(new_n697), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n699), .A2(G99gat), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(new_n798), .B2(new_n820), .ZN(G1338gat));
  NOR3_X1   g620(.A1(new_n709), .A2(new_n571), .A3(G106gat), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n794), .B2(new_n795), .ZN(new_n824));
  INV_X1    g623(.A(G106gat), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(new_n786), .B2(new_n532), .ZN(new_n826));
  OR3_X1    g625(.A1(new_n824), .A2(new_n826), .A3(KEYINPUT53), .ZN(new_n827));
  AOI21_X1  g626(.A(KEYINPUT116), .B1(new_n815), .B2(new_n822), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n829));
  NOR4_X1   g628(.A1(new_n812), .A2(new_n829), .A3(new_n814), .A4(new_n823), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n828), .A2(new_n830), .A3(new_n826), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n827), .B1(new_n831), .B2(new_n832), .ZN(G1339gat));
  NOR2_X1   g632(.A1(new_n566), .A2(new_n460), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n681), .B1(new_n684), .B2(KEYINPUT54), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837));
  INV_X1    g636(.A(new_n672), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n837), .B1(new_n838), .B2(new_n675), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n836), .B1(new_n677), .B2(new_n839), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n840), .A2(KEYINPUT55), .ZN(new_n841));
  AOI22_X1  g640(.A1(new_n840), .A2(KEYINPUT55), .B1(new_n677), .B2(new_n682), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n719), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n246), .A2(new_n266), .A3(new_n263), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n246), .A2(new_n254), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n844), .B1(new_n845), .B2(new_n255), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n273), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(new_n261), .B2(new_n275), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n835), .B1(new_n843), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n275), .ZN(new_n850));
  INV_X1    g649(.A(new_n260), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n258), .ZN(new_n852));
  AOI22_X1  g651(.A1(new_n850), .A2(new_n852), .B1(new_n273), .B2(new_n846), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n840), .A2(KEYINPUT55), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n665), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n853), .A2(KEYINPUT117), .A3(new_n855), .A4(new_n842), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n849), .A2(new_n856), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n841), .B(new_n842), .C1(new_n276), .C2(new_n280), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n853), .A2(new_n687), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n665), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n623), .B1(new_n857), .B2(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n765), .A2(new_n766), .A3(new_n687), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n834), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(new_n572), .ZN(new_n865));
  XOR2_X1   g664(.A(new_n865), .B(KEYINPUT118), .Z(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n285), .A3(new_n766), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n864), .A2(new_n532), .A3(new_n699), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G113gat), .B1(new_n869), .B2(new_n281), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n867), .A2(new_n870), .ZN(G1340gat));
  NAND3_X1  g670(.A1(new_n866), .A2(new_n283), .A3(new_n687), .ZN(new_n872));
  OAI21_X1  g671(.A(G120gat), .B1(new_n869), .B2(new_n709), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1341gat));
  AOI21_X1  g673(.A(new_n289), .B1(new_n868), .B2(new_n623), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n622), .A2(G127gat), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n875), .B1(new_n865), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT119), .ZN(G1342gat));
  NOR2_X1   g677(.A1(new_n864), .A2(new_n665), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n572), .A2(G134gat), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n881), .B(KEYINPUT56), .Z(new_n882));
  OAI21_X1  g681(.A(G134gat), .B1(new_n869), .B2(new_n665), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1343gat));
  NAND2_X1  g683(.A1(new_n697), .A2(new_n834), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n849), .A2(new_n856), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n719), .B1(new_n858), .B2(new_n859), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n622), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n623), .A2(new_n281), .A3(new_n665), .A4(new_n688), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n571), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n885), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n840), .A2(KEYINPUT55), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n683), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n850), .A2(new_n852), .ZN(new_n895));
  INV_X1    g694(.A(new_n274), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n268), .B1(new_n257), .B2(new_n256), .ZN(new_n897));
  INV_X1    g696(.A(new_n279), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n894), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT55), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n840), .A2(KEYINPUT120), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n840), .A2(KEYINPUT120), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI22_X1  g703(.A1(new_n900), .A2(new_n904), .B1(new_n853), .B2(new_n687), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n849), .B(new_n856), .C1(new_n905), .C2(new_n719), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n863), .B1(new_n906), .B2(new_n622), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT57), .B1(new_n907), .B2(new_n571), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n892), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(G141gat), .A3(new_n766), .ZN(new_n910));
  INV_X1    g709(.A(new_n864), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n730), .A2(new_n571), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n913), .A2(new_n281), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n910), .B1(G141gat), .B2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT58), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n915), .B(new_n916), .ZN(G1344gat));
  NAND3_X1  g716(.A1(new_n892), .A2(new_n908), .A3(new_n687), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n919), .A2(G148gat), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n900), .A2(new_n904), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n719), .B1(new_n922), .B2(new_n859), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n843), .A2(new_n848), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n622), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n889), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT57), .B1(new_n926), .B2(new_n532), .ZN(new_n927));
  OAI211_X1 g726(.A(KEYINPUT57), .B(new_n532), .C1(new_n862), .C2(new_n863), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n890), .A2(KEYINPUT121), .A3(KEYINPUT57), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n885), .A2(new_n688), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(G148gat), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n921), .B1(new_n935), .B2(KEYINPUT59), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n913), .A2(G148gat), .A3(new_n688), .ZN(new_n937));
  OAI21_X1  g736(.A(KEYINPUT122), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT122), .ZN(new_n939));
  INV_X1    g738(.A(new_n937), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n926), .A2(new_n532), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n891), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n890), .A2(KEYINPUT121), .A3(KEYINPUT57), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT121), .B1(new_n890), .B2(KEYINPUT57), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n933), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n919), .B1(new_n946), .B2(G148gat), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n939), .B(new_n940), .C1(new_n947), .C2(new_n921), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n938), .A2(new_n948), .ZN(G1345gat));
  INV_X1    g748(.A(new_n909), .ZN(new_n950));
  OAI21_X1  g749(.A(G155gat), .B1(new_n950), .B2(new_n622), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n623), .A2(new_n423), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n913), .B2(new_n952), .ZN(G1346gat));
  INV_X1    g752(.A(KEYINPUT123), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n954), .B1(new_n950), .B2(new_n665), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n909), .A2(KEYINPUT123), .A3(new_n719), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n955), .A2(G162gat), .A3(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n879), .A2(new_n424), .A3(new_n912), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1347gat));
  AOI21_X1  g758(.A(new_n770), .B1(new_n888), .B2(new_n889), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n572), .A2(new_n576), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(G169gat), .B1(new_n962), .B2(new_n766), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n699), .A2(new_n532), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n960), .A2(new_n566), .A3(new_n964), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n965), .A2(new_n329), .A3(new_n281), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n963), .A2(new_n966), .ZN(G1348gat));
  NAND3_X1  g766(.A1(new_n962), .A2(new_n330), .A3(new_n687), .ZN(new_n968));
  OAI21_X1  g767(.A(G176gat), .B1(new_n965), .B2(new_n709), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(G1349gat));
  NAND3_X1  g769(.A1(new_n962), .A2(new_n364), .A3(new_n623), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n312), .A2(new_n314), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n972), .B1(new_n965), .B2(new_n622), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n975));
  XOR2_X1   g774(.A(new_n974), .B(new_n975), .Z(G1350gat));
  OAI21_X1  g775(.A(G190gat), .B1(new_n965), .B2(new_n665), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(KEYINPUT61), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n962), .A2(new_n315), .A3(new_n719), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(G1351gat));
  AND3_X1   g779(.A1(new_n960), .A2(new_n566), .A3(new_n912), .ZN(new_n981));
  INV_X1    g780(.A(G197gat), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n981), .A2(new_n982), .A3(new_n766), .ZN(new_n983));
  XOR2_X1   g782(.A(new_n983), .B(KEYINPUT125), .Z(new_n984));
  NOR2_X1   g783(.A1(new_n576), .A2(new_n770), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n945), .A2(new_n697), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g785(.A(G197gat), .B1(new_n986), .B2(new_n281), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n984), .A2(new_n987), .ZN(G1352gat));
  XNOR2_X1  g787(.A(KEYINPUT126), .B(G204gat), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n981), .A2(new_n687), .A3(new_n989), .ZN(new_n990));
  XOR2_X1   g789(.A(new_n990), .B(KEYINPUT62), .Z(new_n991));
  NOR2_X1   g790(.A1(new_n986), .A2(new_n709), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n991), .B1(new_n992), .B2(new_n989), .ZN(G1353gat));
  NAND3_X1  g792(.A1(new_n981), .A2(new_n474), .A3(new_n623), .ZN(new_n994));
  NAND4_X1  g793(.A1(new_n945), .A2(new_n697), .A3(new_n623), .A4(new_n985), .ZN(new_n995));
  AND3_X1   g794(.A1(new_n995), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n996));
  AOI21_X1  g795(.A(KEYINPUT63), .B1(new_n995), .B2(G211gat), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n994), .B1(new_n996), .B2(new_n997), .ZN(G1354gat));
  OAI21_X1  g797(.A(G218gat), .B1(new_n986), .B2(new_n665), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n981), .A2(new_n475), .A3(new_n719), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(G1355gat));
endmodule


