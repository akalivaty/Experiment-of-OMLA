

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577;

  XOR2_X1 U323 ( .A(KEYINPUT95), .B(n441), .Z(n540) );
  INV_X1 U324 ( .A(KEYINPUT76), .ZN(n346) );
  XNOR2_X1 U325 ( .A(KEYINPUT45), .B(KEYINPUT65), .ZN(n497) );
  XNOR2_X1 U326 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U327 ( .A(n498), .B(n497), .ZN(n501) );
  XNOR2_X1 U328 ( .A(n349), .B(n348), .ZN(n350) );
  NOR2_X1 U329 ( .A1(n507), .A2(n506), .ZN(n508) );
  XOR2_X1 U330 ( .A(n359), .B(n358), .Z(n519) );
  NOR2_X1 U331 ( .A1(n547), .A2(n546), .ZN(n558) );
  NOR2_X1 U332 ( .A1(n459), .A2(n474), .ZN(n452) );
  XNOR2_X1 U333 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n447) );
  XOR2_X1 U334 ( .A(KEYINPUT6), .B(KEYINPUT94), .Z(n296) );
  XOR2_X1 U335 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n292) );
  XNOR2_X1 U336 ( .A(G85GAT), .B(KEYINPUT5), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n294) );
  XNOR2_X1 U338 ( .A(G120GAT), .B(G148GAT), .ZN(n293) );
  XNOR2_X1 U339 ( .A(n293), .B(G57GAT), .ZN(n329) );
  XNOR2_X1 U340 ( .A(n294), .B(n329), .ZN(n295) );
  XNOR2_X1 U341 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U342 ( .A(G29GAT), .B(G134GAT), .Z(n355) );
  XOR2_X1 U343 ( .A(G1GAT), .B(G127GAT), .Z(n373) );
  XOR2_X1 U344 ( .A(n355), .B(n373), .Z(n298) );
  NAND2_X1 U345 ( .A1(G225GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U347 ( .A(n300), .B(n299), .Z(n306) );
  XOR2_X1 U348 ( .A(G113GAT), .B(KEYINPUT0), .Z(n421) );
  XNOR2_X1 U349 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n301), .B(KEYINPUT92), .ZN(n302) );
  XOR2_X1 U351 ( .A(n302), .B(KEYINPUT3), .Z(n304) );
  XNOR2_X1 U352 ( .A(G141GAT), .B(G162GAT), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n304), .B(n303), .ZN(n383) );
  XNOR2_X1 U354 ( .A(n421), .B(n383), .ZN(n305) );
  XNOR2_X1 U355 ( .A(n306), .B(n305), .ZN(n441) );
  XOR2_X1 U356 ( .A(G141GAT), .B(G197GAT), .Z(n308) );
  XNOR2_X1 U357 ( .A(G36GAT), .B(G29GAT), .ZN(n307) );
  XNOR2_X1 U358 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U359 ( .A(n309), .B(G113GAT), .Z(n311) );
  XOR2_X1 U360 ( .A(G22GAT), .B(G15GAT), .Z(n374) );
  XNOR2_X1 U361 ( .A(G169GAT), .B(n374), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n317) );
  XOR2_X1 U363 ( .A(G43GAT), .B(G50GAT), .Z(n313) );
  XNOR2_X1 U364 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n313), .B(n312), .ZN(n349) );
  XOR2_X1 U366 ( .A(n349), .B(KEYINPUT67), .Z(n315) );
  NAND2_X1 U367 ( .A1(G229GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U369 ( .A(n317), .B(n316), .Z(n325) );
  XOR2_X1 U370 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n319) );
  XNOR2_X1 U371 ( .A(G1GAT), .B(G8GAT), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U373 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n321) );
  XNOR2_X1 U374 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n320) );
  XNOR2_X1 U375 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n563) );
  XOR2_X1 U378 ( .A(KEYINPUT72), .B(KEYINPUT33), .Z(n331) );
  XOR2_X1 U379 ( .A(KEYINPUT73), .B(KEYINPUT31), .Z(n327) );
  XNOR2_X1 U380 ( .A(KEYINPUT74), .B(KEYINPUT32), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U384 ( .A(G71GAT), .B(KEYINPUT13), .Z(n366) );
  XOR2_X1 U385 ( .A(G99GAT), .B(G85GAT), .Z(n343) );
  XOR2_X1 U386 ( .A(n366), .B(n343), .Z(n333) );
  NAND2_X1 U387 ( .A1(G230GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U389 ( .A(n335), .B(n334), .Z(n340) );
  XOR2_X1 U390 ( .A(G106GAT), .B(G78GAT), .Z(n393) );
  XOR2_X1 U391 ( .A(G92GAT), .B(G64GAT), .Z(n337) );
  XNOR2_X1 U392 ( .A(G204GAT), .B(KEYINPUT75), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U394 ( .A(G176GAT), .B(n338), .Z(n407) );
  XNOR2_X1 U395 ( .A(n393), .B(n407), .ZN(n339) );
  XNOR2_X1 U396 ( .A(n340), .B(n339), .ZN(n499) );
  NAND2_X1 U397 ( .A1(n563), .A2(n499), .ZN(n459) );
  XOR2_X1 U398 ( .A(KEYINPUT66), .B(KEYINPUT11), .Z(n342) );
  XNOR2_X1 U399 ( .A(KEYINPUT10), .B(KEYINPUT9), .ZN(n341) );
  XNOR2_X1 U400 ( .A(n342), .B(n341), .ZN(n359) );
  XOR2_X1 U401 ( .A(G36GAT), .B(G190GAT), .Z(n403) );
  XOR2_X1 U402 ( .A(n343), .B(n403), .Z(n345) );
  XNOR2_X1 U403 ( .A(G218GAT), .B(G92GAT), .ZN(n344) );
  XNOR2_X1 U404 ( .A(n345), .B(n344), .ZN(n351) );
  NAND2_X1 U405 ( .A1(G232GAT), .A2(G233GAT), .ZN(n347) );
  XOR2_X1 U406 ( .A(n351), .B(n350), .Z(n357) );
  XOR2_X1 U407 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n353) );
  XNOR2_X1 U408 ( .A(G162GAT), .B(G106GAT), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U410 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U412 ( .A(G64GAT), .B(G57GAT), .Z(n361) );
  XNOR2_X1 U413 ( .A(G183GAT), .B(G78GAT), .ZN(n360) );
  XNOR2_X1 U414 ( .A(n361), .B(n360), .ZN(n365) );
  XOR2_X1 U415 ( .A(KEYINPUT82), .B(KEYINPUT80), .Z(n363) );
  XNOR2_X1 U416 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U418 ( .A(n365), .B(n364), .ZN(n378) );
  XOR2_X1 U419 ( .A(G8GAT), .B(KEYINPUT79), .Z(n402) );
  XOR2_X1 U420 ( .A(n366), .B(n402), .Z(n368) );
  XNOR2_X1 U421 ( .A(G211GAT), .B(G155GAT), .ZN(n367) );
  XNOR2_X1 U422 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U423 ( .A(KEYINPUT15), .B(KEYINPUT81), .Z(n370) );
  NAND2_X1 U424 ( .A1(G231GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U425 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U426 ( .A(n372), .B(n371), .Z(n376) );
  XNOR2_X1 U427 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U428 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U429 ( .A(n378), .B(n377), .ZN(n570) );
  NAND2_X1 U430 ( .A1(n519), .A2(n570), .ZN(n379) );
  XOR2_X1 U431 ( .A(KEYINPUT16), .B(n379), .Z(n445) );
  XOR2_X1 U432 ( .A(KEYINPUT91), .B(G218GAT), .Z(n381) );
  XNOR2_X1 U433 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n380) );
  XNOR2_X1 U434 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U435 ( .A(G197GAT), .B(n382), .Z(n411) );
  XNOR2_X1 U436 ( .A(n411), .B(n383), .ZN(n397) );
  XOR2_X1 U437 ( .A(KEYINPUT90), .B(KEYINPUT93), .Z(n385) );
  XNOR2_X1 U438 ( .A(G50GAT), .B(G22GAT), .ZN(n384) );
  XNOR2_X1 U439 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U440 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n387) );
  XNOR2_X1 U441 ( .A(G204GAT), .B(G148GAT), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U443 ( .A(n389), .B(n388), .Z(n395) );
  XOR2_X1 U444 ( .A(KEYINPUT89), .B(KEYINPUT22), .Z(n391) );
  NAND2_X1 U445 ( .A1(G228GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U446 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U447 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U448 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U449 ( .A(n397), .B(n396), .ZN(n543) );
  XOR2_X1 U450 ( .A(n543), .B(KEYINPUT28), .Z(n492) );
  XNOR2_X1 U451 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n398) );
  XNOR2_X1 U452 ( .A(n398), .B(KEYINPUT86), .ZN(n399) );
  XOR2_X1 U453 ( .A(n399), .B(KEYINPUT18), .Z(n401) );
  XNOR2_X1 U454 ( .A(G169GAT), .B(G183GAT), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n431) );
  XOR2_X1 U456 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n405) );
  XNOR2_X1 U457 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U458 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U459 ( .A(n407), .B(n406), .Z(n409) );
  NAND2_X1 U460 ( .A1(G226GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U461 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U462 ( .A(n431), .B(n410), .ZN(n412) );
  XOR2_X1 U463 ( .A(n412), .B(n411), .Z(n536) );
  XNOR2_X1 U464 ( .A(KEYINPUT27), .B(n536), .ZN(n437) );
  NAND2_X1 U465 ( .A1(n540), .A2(n437), .ZN(n525) );
  NOR2_X1 U466 ( .A1(n492), .A2(n525), .ZN(n509) );
  XNOR2_X1 U467 ( .A(n509), .B(KEYINPUT98), .ZN(n432) );
  XOR2_X1 U468 ( .A(KEYINPUT87), .B(G120GAT), .Z(n414) );
  XNOR2_X1 U469 ( .A(G15GAT), .B(KEYINPUT83), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U471 ( .A(KEYINPUT20), .B(G176GAT), .Z(n416) );
  XNOR2_X1 U472 ( .A(G43GAT), .B(G134GAT), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U474 ( .A(n418), .B(n417), .ZN(n429) );
  XOR2_X1 U475 ( .A(KEYINPUT84), .B(G127GAT), .Z(n420) );
  XNOR2_X1 U476 ( .A(KEYINPUT85), .B(KEYINPUT88), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n425) );
  XOR2_X1 U478 ( .A(G190GAT), .B(G99GAT), .Z(n423) );
  XNOR2_X1 U479 ( .A(G71GAT), .B(n421), .ZN(n422) );
  XNOR2_X1 U480 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U481 ( .A(n425), .B(n424), .Z(n427) );
  NAND2_X1 U482 ( .A1(G227GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U484 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U485 ( .A(n431), .B(n430), .ZN(n546) );
  NAND2_X1 U486 ( .A1(n432), .A2(n546), .ZN(n444) );
  INV_X1 U487 ( .A(n546), .ZN(n489) );
  NAND2_X1 U488 ( .A1(n489), .A2(n536), .ZN(n433) );
  XOR2_X1 U489 ( .A(KEYINPUT99), .B(n433), .Z(n434) );
  NAND2_X1 U490 ( .A1(n543), .A2(n434), .ZN(n435) );
  XNOR2_X1 U491 ( .A(n435), .B(KEYINPUT25), .ZN(n439) );
  NOR2_X1 U492 ( .A1(n543), .A2(n489), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n436), .B(KEYINPUT26), .ZN(n561) );
  AND2_X1 U494 ( .A1(n437), .A2(n561), .ZN(n438) );
  NOR2_X1 U495 ( .A1(n439), .A2(n438), .ZN(n440) );
  NOR2_X1 U496 ( .A1(n441), .A2(n440), .ZN(n442) );
  XOR2_X1 U497 ( .A(KEYINPUT100), .B(n442), .Z(n443) );
  NAND2_X1 U498 ( .A1(n444), .A2(n443), .ZN(n455) );
  NAND2_X1 U499 ( .A1(n445), .A2(n455), .ZN(n474) );
  NAND2_X1 U500 ( .A1(n540), .A2(n452), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n447), .B(n446), .ZN(G1324GAT) );
  XOR2_X1 U502 ( .A(G8GAT), .B(KEYINPUT101), .Z(n449) );
  NAND2_X1 U503 ( .A1(n452), .A2(n536), .ZN(n448) );
  XNOR2_X1 U504 ( .A(n449), .B(n448), .ZN(G1325GAT) );
  XOR2_X1 U505 ( .A(G15GAT), .B(KEYINPUT35), .Z(n451) );
  NAND2_X1 U506 ( .A1(n452), .A2(n489), .ZN(n450) );
  XNOR2_X1 U507 ( .A(n451), .B(n450), .ZN(G1326GAT) );
  NAND2_X1 U508 ( .A1(n452), .A2(n492), .ZN(n453) );
  XNOR2_X1 U509 ( .A(n453), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U510 ( .A(G29GAT), .B(KEYINPUT102), .Z(n462) );
  XNOR2_X1 U511 ( .A(n519), .B(KEYINPUT103), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n454), .B(KEYINPUT36), .ZN(n574) );
  NAND2_X1 U513 ( .A1(n574), .A2(n455), .ZN(n456) );
  NOR2_X1 U514 ( .A1(n570), .A2(n456), .ZN(n458) );
  XNOR2_X1 U515 ( .A(KEYINPUT104), .B(KEYINPUT37), .ZN(n457) );
  XNOR2_X1 U516 ( .A(n458), .B(n457), .ZN(n485) );
  NOR2_X1 U517 ( .A1(n459), .A2(n485), .ZN(n460) );
  XNOR2_X1 U518 ( .A(n460), .B(KEYINPUT38), .ZN(n470) );
  NAND2_X1 U519 ( .A1(n540), .A2(n470), .ZN(n461) );
  XNOR2_X1 U520 ( .A(n462), .B(n461), .ZN(n464) );
  XOR2_X1 U521 ( .A(KEYINPUT39), .B(KEYINPUT105), .Z(n463) );
  XNOR2_X1 U522 ( .A(n464), .B(n463), .ZN(G1328GAT) );
  NAND2_X1 U523 ( .A1(n470), .A2(n536), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n465), .B(KEYINPUT106), .ZN(n466) );
  XNOR2_X1 U525 ( .A(G36GAT), .B(n466), .ZN(G1329GAT) );
  XOR2_X1 U526 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n468) );
  NAND2_X1 U527 ( .A1(n489), .A2(n470), .ZN(n467) );
  XNOR2_X1 U528 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U529 ( .A(G43GAT), .B(n469), .ZN(G1330GAT) );
  NAND2_X1 U530 ( .A1(n470), .A2(n492), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n471), .B(KEYINPUT108), .ZN(n472) );
  XNOR2_X1 U532 ( .A(G50GAT), .B(n472), .ZN(G1331GAT) );
  XOR2_X1 U533 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n477) );
  INV_X1 U534 ( .A(n563), .ZN(n473) );
  XNOR2_X1 U535 ( .A(n499), .B(KEYINPUT41), .ZN(n550) );
  NAND2_X1 U536 ( .A1(n473), .A2(n550), .ZN(n484) );
  NOR2_X1 U537 ( .A1(n484), .A2(n474), .ZN(n475) );
  XOR2_X1 U538 ( .A(KEYINPUT109), .B(n475), .Z(n481) );
  NAND2_X1 U539 ( .A1(n481), .A2(n540), .ZN(n476) );
  XNOR2_X1 U540 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U541 ( .A(G57GAT), .B(n478), .Z(G1332GAT) );
  NAND2_X1 U542 ( .A1(n536), .A2(n481), .ZN(n479) );
  XNOR2_X1 U543 ( .A(n479), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U544 ( .A1(n481), .A2(n489), .ZN(n480) );
  XNOR2_X1 U545 ( .A(n480), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U546 ( .A(G78GAT), .B(KEYINPUT43), .Z(n483) );
  NAND2_X1 U547 ( .A1(n481), .A2(n492), .ZN(n482) );
  XNOR2_X1 U548 ( .A(n483), .B(n482), .ZN(G1335GAT) );
  XOR2_X1 U549 ( .A(G85GAT), .B(KEYINPUT111), .Z(n487) );
  NOR2_X1 U550 ( .A1(n485), .A2(n484), .ZN(n493) );
  NAND2_X1 U551 ( .A1(n493), .A2(n540), .ZN(n486) );
  XNOR2_X1 U552 ( .A(n487), .B(n486), .ZN(G1336GAT) );
  NAND2_X1 U553 ( .A1(n536), .A2(n493), .ZN(n488) );
  XNOR2_X1 U554 ( .A(n488), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U555 ( .A1(n493), .A2(n489), .ZN(n490) );
  XNOR2_X1 U556 ( .A(n490), .B(KEYINPUT112), .ZN(n491) );
  XNOR2_X1 U557 ( .A(G99GAT), .B(n491), .ZN(G1338GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n495) );
  NAND2_X1 U559 ( .A1(n493), .A2(n492), .ZN(n494) );
  XNOR2_X1 U560 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U561 ( .A(G106GAT), .B(n496), .ZN(G1339GAT) );
  NAND2_X1 U562 ( .A1(n574), .A2(n570), .ZN(n498) );
  INV_X1 U563 ( .A(n499), .ZN(n567) );
  NOR2_X1 U564 ( .A1(n567), .A2(n563), .ZN(n500) );
  AND2_X1 U565 ( .A1(n501), .A2(n500), .ZN(n507) );
  NAND2_X1 U566 ( .A1(n563), .A2(n550), .ZN(n502) );
  XOR2_X1 U567 ( .A(KEYINPUT46), .B(n502), .Z(n503) );
  NOR2_X1 U568 ( .A1(n570), .A2(n503), .ZN(n504) );
  NAND2_X1 U569 ( .A1(n519), .A2(n504), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n505), .B(KEYINPUT47), .ZN(n506) );
  XOR2_X1 U571 ( .A(KEYINPUT48), .B(n508), .Z(n537) );
  NAND2_X1 U572 ( .A1(n537), .A2(n509), .ZN(n510) );
  NOR2_X1 U573 ( .A1(n546), .A2(n510), .ZN(n520) );
  NAND2_X1 U574 ( .A1(n520), .A2(n563), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n511), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n513) );
  NAND2_X1 U577 ( .A1(n520), .A2(n550), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G120GAT), .B(n514), .ZN(G1341GAT) );
  NAND2_X1 U580 ( .A1(n520), .A2(n570), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n515), .B(KEYINPUT50), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G127GAT), .B(n516), .ZN(G1342GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n518) );
  XNOR2_X1 U584 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(n523) );
  INV_X1 U586 ( .A(n519), .ZN(n557) );
  NAND2_X1 U587 ( .A1(n557), .A2(n520), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n521), .B(KEYINPUT115), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(G1343GAT) );
  NAND2_X1 U590 ( .A1(n537), .A2(n561), .ZN(n524) );
  NOR2_X1 U591 ( .A1(n525), .A2(n524), .ZN(n534) );
  NAND2_X1 U592 ( .A1(n534), .A2(n563), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n526), .B(G141GAT), .ZN(G1344GAT) );
  NAND2_X1 U594 ( .A1(n550), .A2(n534), .ZN(n532) );
  XOR2_X1 U595 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n528) );
  XNOR2_X1 U596 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n527) );
  XNOR2_X1 U597 ( .A(n528), .B(n527), .ZN(n530) );
  XOR2_X1 U598 ( .A(G148GAT), .B(KEYINPUT52), .Z(n529) );
  XNOR2_X1 U599 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U600 ( .A(n532), .B(n531), .ZN(G1345GAT) );
  NAND2_X1 U601 ( .A1(n534), .A2(n570), .ZN(n533) );
  XNOR2_X1 U602 ( .A(n533), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U603 ( .A1(n557), .A2(n534), .ZN(n535) );
  XNOR2_X1 U604 ( .A(n535), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U605 ( .A(KEYINPUT55), .B(KEYINPUT122), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n537), .A2(n536), .ZN(n539) );
  XOR2_X1 U607 ( .A(KEYINPUT121), .B(KEYINPUT54), .Z(n538) );
  XNOR2_X1 U608 ( .A(n539), .B(n538), .ZN(n541) );
  NOR2_X1 U609 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n542), .B(KEYINPUT64), .ZN(n562) );
  AND2_X1 U611 ( .A1(n543), .A2(n562), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n547) );
  NAND2_X1 U613 ( .A1(n558), .A2(n563), .ZN(n549) );
  XOR2_X1 U614 ( .A(G169GAT), .B(KEYINPUT123), .Z(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(G1348GAT) );
  NAND2_X1 U616 ( .A1(n558), .A2(n550), .ZN(n555) );
  XOR2_X1 U617 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n552) );
  XNOR2_X1 U618 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U620 ( .A(KEYINPUT56), .B(n553), .Z(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1349GAT) );
  NAND2_X1 U622 ( .A1(n558), .A2(n570), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U624 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1351GAT) );
  AND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n573) );
  NAND2_X1 U628 ( .A1(n573), .A2(n563), .ZN(n565) );
  XOR2_X1 U629 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(G197GAT), .ZN(G1352GAT) );
  XOR2_X1 U632 ( .A(G204GAT), .B(KEYINPUT61), .Z(n569) );
  NAND2_X1 U633 ( .A1(n573), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1353GAT) );
  NAND2_X1 U635 ( .A1(n573), .A2(n570), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(KEYINPUT126), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G211GAT), .B(n572), .ZN(G1354GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n576) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(G218GAT), .ZN(G1355GAT) );
endmodule

