//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1191, new_n1192, new_n1193, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n207), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT66), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n210), .B1(new_n212), .B2(new_n216), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT1), .Z(new_n218));
  NOR2_X1   g0018(.A1(new_n210), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT0), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  OR2_X1    g0025(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n226), .A2(G50), .A3(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n218), .B(new_n221), .C1(new_n225), .C2(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT67), .Z(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT68), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n235), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G50), .B(G68), .Z(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(G97), .B(G107), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G274), .ZN(new_n249));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n250), .B1(G41), .B2(G45), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT71), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n252), .B1(new_n254), .B2(new_n222), .ZN(new_n255));
  INV_X1    g0055(.A(new_n222), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(KEYINPUT71), .A3(new_n253), .ZN(new_n257));
  AOI211_X1 g0057(.A(new_n249), .B(new_n251), .C1(new_n255), .C2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT3), .B(G33), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(G222), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G77), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(G1698), .ZN(new_n263));
  INV_X1    g0063(.A(G223), .ZN(new_n264));
  OAI221_X1 g0064(.A(new_n261), .B1(new_n262), .B2(new_n259), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n254), .A2(new_n222), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n258), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NOR3_X1   g0067(.A1(new_n254), .A2(new_n252), .A3(new_n222), .ZN(new_n268));
  AOI21_X1  g0068(.A(KEYINPUT71), .B1(new_n256), .B2(new_n253), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n251), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT72), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n255), .A2(new_n257), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT72), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(new_n273), .A3(new_n251), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n271), .A2(G226), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n267), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(G179), .ZN(new_n277));
  AOI21_X1  g0077(.A(G169), .B1(new_n267), .B2(new_n275), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n250), .A2(G20), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G50), .ZN(new_n280));
  XNOR2_X1  g0080(.A(new_n280), .B(KEYINPUT73), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n250), .A2(G13), .A3(G20), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n222), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G50), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n281), .A2(new_n286), .B1(new_n287), .B2(new_n283), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n223), .B1(new_n206), .B2(new_n287), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT8), .B(G58), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n223), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(G150), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G20), .A2(G33), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI22_X1  g0094(.A1(new_n290), .A2(new_n291), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n285), .B1(new_n289), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n288), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n277), .A2(new_n278), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n297), .B(KEYINPUT9), .ZN(new_n300));
  INV_X1    g0100(.A(G200), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(new_n267), .B2(new_n275), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G190), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n300), .B(new_n303), .C1(new_n304), .C2(new_n276), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n299), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G33), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT3), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT3), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G33), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n310), .A2(new_n312), .A3(G226), .A4(G1698), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n310), .A2(new_n312), .A3(G223), .A4(new_n260), .ZN(new_n314));
  INV_X1    g0114(.A(G87), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n313), .B(new_n314), .C1(new_n309), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n266), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n249), .B1(new_n255), .B2(new_n257), .ZN(new_n318));
  INV_X1    g0118(.A(new_n251), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n272), .A2(G232), .A3(new_n251), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n317), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n301), .ZN(new_n323));
  AND3_X1   g0123(.A1(new_n316), .A2(KEYINPUT78), .A3(new_n266), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT78), .B1(new_n316), .B2(new_n266), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n320), .A2(new_n304), .A3(new_n321), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n323), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n202), .A2(new_n203), .ZN(new_n329));
  OAI21_X1  g0129(.A(G20), .B1(new_n206), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n293), .A2(G159), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n310), .A2(new_n312), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(KEYINPUT7), .A3(new_n223), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n310), .A2(new_n312), .A3(KEYINPUT77), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT77), .B1(new_n310), .B2(new_n312), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n223), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT7), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n336), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(KEYINPUT16), .B(new_n333), .C1(new_n341), .C2(new_n203), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT16), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n340), .B1(new_n259), .B2(G20), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n203), .B1(new_n344), .B2(new_n335), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n343), .B1(new_n345), .B2(new_n332), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n342), .A2(new_n285), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n285), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n279), .ZN(new_n349));
  INV_X1    g0149(.A(new_n290), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n283), .B2(new_n350), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n328), .A2(new_n347), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT17), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT17), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n328), .A2(new_n347), .A3(new_n355), .A4(new_n352), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G169), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n322), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G179), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n320), .A2(new_n360), .A3(new_n321), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n359), .B1(new_n326), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n347), .B2(new_n352), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(KEYINPUT18), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n347), .A2(new_n352), .ZN(new_n365));
  INV_X1    g0165(.A(new_n362), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n365), .A2(new_n366), .A3(KEYINPUT18), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n357), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n310), .A2(new_n312), .A3(G226), .A4(new_n260), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT75), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n259), .A2(KEYINPUT75), .A3(G226), .A4(new_n260), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G33), .A2(G97), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n259), .A2(G232), .A3(G1698), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n372), .A2(new_n373), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n258), .B1(new_n376), .B2(new_n266), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n271), .A2(G238), .A3(new_n274), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT13), .ZN(new_n379));
  AND3_X1   g0179(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n379), .B1(new_n377), .B2(new_n378), .ZN(new_n381));
  OAI21_X1  g0181(.A(G200), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n377), .A2(new_n378), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT13), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(G190), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n291), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n387), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n293), .A2(G50), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n348), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g0190(.A(new_n390), .B(KEYINPUT11), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT76), .B1(new_n283), .B2(new_n203), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n392), .B(KEYINPUT12), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n203), .B2(new_n349), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n382), .A2(new_n386), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(G169), .B1(new_n380), .B2(new_n381), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT14), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT14), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n400), .B(G169), .C1(new_n380), .C2(new_n381), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n384), .A2(G179), .A3(new_n385), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n395), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n397), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n283), .A2(new_n262), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n349), .B2(new_n262), .ZN(new_n407));
  OAI22_X1  g0207(.A1(new_n290), .A2(new_n294), .B1(new_n223), .B2(new_n262), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT74), .ZN(new_n409));
  XOR2_X1   g0209(.A(KEYINPUT15), .B(G87), .Z(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n387), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n408), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n409), .B2(new_n411), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n407), .B1(new_n413), .B2(new_n285), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n259), .A2(G232), .A3(new_n260), .ZN(new_n415));
  INV_X1    g0215(.A(G107), .ZN(new_n416));
  INV_X1    g0216(.A(G238), .ZN(new_n417));
  OAI221_X1 g0217(.A(new_n415), .B1(new_n416), .B2(new_n259), .C1(new_n263), .C2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n258), .B1(new_n418), .B2(new_n266), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n271), .A2(G244), .A3(new_n274), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n414), .B1(new_n421), .B2(new_n358), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n419), .A2(new_n360), .A3(new_n420), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n421), .A2(G200), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n425), .B(new_n414), .C1(new_n304), .C2(new_n421), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n308), .A2(new_n369), .A3(new_n405), .A4(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G41), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n250), .B(G45), .C1(new_n429), .C2(KEYINPUT5), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT81), .ZN(new_n431));
  INV_X1    g0231(.A(G45), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n432), .A2(G1), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT81), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT5), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G41), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n433), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT82), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n435), .B2(G41), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n429), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n431), .A2(new_n437), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n259), .A2(G257), .A3(new_n260), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n259), .A2(G264), .A3(G1698), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n334), .A2(G303), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n442), .A2(new_n318), .B1(new_n446), .B2(new_n266), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n441), .A2(G270), .A3(new_n272), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT84), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT84), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n441), .A2(new_n450), .A3(G270), .A4(new_n272), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n447), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G283), .ZN(new_n453));
  INV_X1    g0253(.A(G97), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n453), .B(new_n223), .C1(G33), .C2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n455), .B(new_n285), .C1(new_n223), .C2(G116), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT20), .ZN(new_n457));
  XNOR2_X1  g0257(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n282), .A2(G116), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n309), .A2(G1), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n283), .A2(new_n285), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n459), .B1(new_n461), .B2(G116), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n358), .B1(new_n458), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n452), .A2(KEYINPUT21), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT21), .B1(new_n452), .B2(new_n463), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n447), .A2(new_n449), .A3(G179), .A4(new_n451), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n458), .A2(new_n462), .ZN(new_n469));
  OR3_X1    g0269(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT85), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT85), .B1(new_n468), .B2(new_n469), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT25), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n282), .A2(new_n472), .A3(G107), .ZN(new_n473));
  OR2_X1    g0273(.A1(new_n473), .A2(KEYINPUT87), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(KEYINPUT87), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n472), .B1(new_n282), .B2(G107), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n461), .A2(G107), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT23), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n480), .A2(new_n223), .A3(G107), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT23), .B1(new_n416), .B2(G20), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G116), .ZN(new_n483));
  OAI22_X1  g0283(.A1(new_n481), .A2(new_n482), .B1(G20), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n259), .A2(new_n223), .A3(G87), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT22), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(KEYINPUT86), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n487), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n259), .A2(new_n489), .A3(new_n223), .A4(G87), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n484), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n491), .A2(KEYINPUT24), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n285), .B1(new_n491), .B2(KEYINPUT24), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n479), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n442), .A2(new_n318), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n441), .A2(G264), .A3(new_n272), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n259), .A2(G250), .A3(new_n260), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n259), .A2(G257), .A3(G1698), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G294), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n266), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n495), .A2(new_n496), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n358), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n501), .A2(new_n496), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(new_n360), .A3(new_n495), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n494), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n467), .A2(new_n470), .A3(new_n471), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n502), .A2(G200), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n495), .A2(new_n501), .A3(G190), .A4(new_n496), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(new_n494), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT19), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(new_n291), .B2(new_n454), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT83), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n259), .A2(new_n223), .A3(G68), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT83), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n516), .B(new_n512), .C1(new_n291), .C2(new_n454), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n223), .B1(new_n374), .B2(new_n512), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n315), .A2(new_n454), .A3(new_n416), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n514), .A2(new_n515), .A3(new_n517), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n285), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n461), .A2(G87), .ZN(new_n523));
  INV_X1    g0323(.A(new_n410), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n283), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n259), .A2(G238), .A3(new_n260), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n259), .A2(G244), .A3(G1698), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(new_n529), .A3(new_n483), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n266), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n433), .A2(new_n249), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n272), .B(new_n532), .C1(G250), .C2(new_n433), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n301), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n531), .A2(G190), .A3(new_n533), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n527), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n531), .A2(new_n533), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n358), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n461), .A2(new_n410), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n522), .A2(new_n525), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n531), .A2(new_n360), .A3(new_n533), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n511), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n461), .A2(G97), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT80), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n282), .B2(G97), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n283), .A2(KEYINPUT80), .A3(new_n454), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT6), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n551), .A2(new_n454), .A3(G107), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(new_n551), .B2(new_n246), .ZN(new_n553));
  OAI22_X1  g0353(.A1(new_n553), .A2(new_n223), .B1(new_n262), .B2(new_n294), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n416), .B1(new_n344), .B2(new_n335), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n285), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(KEYINPUT79), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(KEYINPUT79), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n550), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n441), .A2(G257), .A3(new_n272), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n495), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n259), .A2(G244), .A3(new_n260), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT4), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n259), .A2(KEYINPUT4), .A3(G244), .A4(new_n260), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n259), .A2(G250), .A3(G1698), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n566), .A2(new_n453), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n266), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n563), .A2(new_n304), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n562), .B1(new_n266), .B2(new_n569), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n571), .B1(new_n572), .B2(G200), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n560), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n550), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n294), .A2(new_n262), .ZN(new_n576));
  INV_X1    g0376(.A(new_n552), .ZN(new_n577));
  INV_X1    g0377(.A(new_n246), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n577), .B1(new_n578), .B2(KEYINPUT6), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n576), .B1(new_n579), .B2(G20), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n344), .A2(new_n335), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G107), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n348), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT79), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n575), .B1(new_n585), .B2(new_n557), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n572), .A2(new_n360), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n563), .A2(new_n570), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n358), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n452), .A2(G200), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n447), .A2(new_n449), .A3(G190), .A4(new_n451), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n469), .A3(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n545), .A2(new_n574), .A3(new_n590), .A4(new_n593), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n428), .A2(new_n507), .A3(new_n594), .ZN(G372));
  NOR2_X1   g0395(.A1(new_n364), .A2(new_n367), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n424), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n403), .B2(new_n404), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n357), .A2(new_n396), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n597), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n306), .A2(new_n307), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n299), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n574), .A2(new_n590), .ZN(new_n607));
  INV_X1    g0407(.A(new_n511), .ZN(new_n608));
  INV_X1    g0408(.A(new_n543), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n526), .A2(new_n534), .ZN(new_n610));
  INV_X1    g0410(.A(new_n538), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n610), .A2(KEYINPUT88), .B1(G190), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT88), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n526), .B2(new_n534), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n609), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n607), .A2(new_n507), .A3(new_n608), .A4(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n617), .A2(new_n615), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT26), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(KEYINPUT26), .B1(new_n590), .B2(new_n544), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n616), .A2(new_n620), .A3(new_n543), .A4(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n606), .B1(new_n428), .B2(new_n623), .ZN(G369));
  INV_X1    g0424(.A(G13), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n625), .A2(G20), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n250), .ZN(new_n627));
  OR2_X1    g0427(.A1(new_n627), .A2(KEYINPUT27), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(KEYINPUT27), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(G213), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(G343), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n469), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n633), .B(KEYINPUT89), .ZN(new_n634));
  INV_X1    g0434(.A(new_n466), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n470), .A2(new_n635), .A3(new_n471), .A4(new_n464), .ZN(new_n636));
  INV_X1    g0436(.A(new_n593), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n636), .B2(new_n634), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n639), .B(KEYINPUT90), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n640), .A2(G330), .ZN(new_n641));
  INV_X1    g0441(.A(new_n632), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n506), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n494), .A2(new_n642), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n506), .B1(new_n645), .B2(new_n511), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n641), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n636), .A2(new_n632), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n649), .A2(new_n644), .A3(new_n651), .ZN(G399));
  INV_X1    g0452(.A(new_n219), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(G41), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n519), .A2(G116), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(G1), .A3(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n228), .B2(new_n655), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(KEYINPUT28), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n615), .A2(new_n574), .A3(new_n590), .A4(new_n608), .ZN(new_n660));
  INV_X1    g0460(.A(new_n506), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n636), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n543), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n617), .A2(new_n619), .A3(new_n537), .A4(new_n543), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n618), .B2(new_n619), .ZN(new_n665));
  OAI211_X1 g0465(.A(KEYINPUT29), .B(new_n632), .C1(new_n663), .C2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(KEYINPUT29), .B1(new_n622), .B2(new_n632), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT91), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT91), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n637), .A2(new_n511), .A3(new_n544), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n662), .A2(new_n607), .A3(new_n673), .A4(new_n632), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT31), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT30), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n563), .A2(new_n611), .A3(new_n504), .A4(new_n570), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n676), .B1(new_n677), .B2(new_n468), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n611), .A2(new_n504), .ZN(new_n679));
  INV_X1    g0479(.A(new_n468), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n679), .A2(new_n680), .A3(KEYINPUT30), .A4(new_n572), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n611), .A2(G179), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n588), .A2(new_n682), .A3(new_n452), .A4(new_n502), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n678), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n675), .B1(new_n684), .B2(new_n642), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n674), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n684), .A2(new_n675), .A3(new_n642), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G330), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n672), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n659), .B1(new_n690), .B2(G1), .ZN(G364));
  NOR2_X1   g0491(.A1(new_n640), .A2(G330), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n250), .B1(new_n626), .B2(G45), .ZN(new_n693));
  AOI211_X1 g0493(.A(new_n692), .B(new_n641), .C1(new_n655), .C2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n653), .A2(new_n334), .ZN(new_n695));
  INV_X1    g0495(.A(G116), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n695), .A2(G355), .B1(new_n696), .B2(new_n653), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n228), .A2(G45), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT77), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n311), .A2(G33), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n309), .A2(KEYINPUT3), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n310), .A2(new_n312), .A3(KEYINPUT77), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n653), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n244), .B2(new_n432), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n697), .B1(new_n698), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(G20), .B1(KEYINPUT92), .B2(G169), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(KEYINPUT92), .A2(G169), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n222), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(G13), .A2(G33), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G20), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n708), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n693), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n654), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n223), .A2(new_n304), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n360), .A2(new_n301), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n223), .A2(G190), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI22_X1  g0526(.A1(G50), .A2(new_n723), .B1(new_n726), .B2(G68), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n360), .A2(G200), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n720), .A2(new_n728), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT93), .Z(new_n731));
  OAI221_X1 g0531(.A(new_n727), .B1(new_n262), .B2(new_n729), .C1(new_n731), .C2(new_n202), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G179), .A2(G200), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G190), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n454), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT32), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n724), .A2(new_n733), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n738), .B1(new_n740), .B2(G159), .ZN(new_n741));
  INV_X1    g0541(.A(G159), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n739), .A2(KEYINPUT32), .A3(new_n742), .ZN(new_n743));
  NOR4_X1   g0543(.A1(new_n732), .A2(new_n737), .A3(new_n741), .A4(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n301), .A2(G179), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n724), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n720), .A2(new_n745), .ZN(new_n747));
  OAI221_X1 g0547(.A(new_n259), .B1(new_n746), .B2(new_n416), .C1(new_n315), .C2(new_n747), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT94), .ZN(new_n749));
  INV_X1    g0549(.A(new_n746), .ZN(new_n750));
  AOI22_X1  g0550(.A1(G283), .A2(new_n750), .B1(new_n740), .B2(G329), .ZN(new_n751));
  INV_X1    g0551(.A(G322), .ZN(new_n752));
  XOR2_X1   g0552(.A(KEYINPUT33), .B(G317), .Z(new_n753));
  OAI221_X1 g0553(.A(new_n751), .B1(new_n752), .B2(new_n730), .C1(new_n725), .C2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n747), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n259), .B1(new_n755), .B2(G303), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n757), .A2(KEYINPUT96), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(KEYINPUT96), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n754), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G326), .ZN(new_n761));
  INV_X1    g0561(.A(G311), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n722), .A2(new_n761), .B1(new_n729), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(G294), .B2(new_n735), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT95), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n744), .A2(new_n749), .B1(new_n760), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n712), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n719), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n715), .B(KEYINPUT97), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n717), .B(new_n768), .C1(new_n639), .C2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n694), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(G396));
  INV_X1    g0572(.A(G132), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n705), .B1(new_n773), .B2(new_n739), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n750), .A2(G68), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(new_n287), .B2(new_n747), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT99), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n774), .B(new_n777), .C1(G58), .C2(new_n735), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT100), .Z(new_n779));
  INV_X1    g0579(.A(new_n729), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G137), .A2(new_n723), .B1(new_n780), .B2(G159), .ZN(new_n781));
  INV_X1    g0581(.A(G143), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n781), .B1(new_n292), .B2(new_n725), .C1(new_n731), .C2(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT34), .Z(new_n784));
  NOR2_X1   g0584(.A1(new_n779), .A2(new_n784), .ZN(new_n785));
  AOI22_X1  g0585(.A1(G87), .A2(new_n750), .B1(new_n740), .B2(G311), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n786), .B1(new_n416), .B2(new_n747), .C1(new_n696), .C2(new_n729), .ZN(new_n787));
  INV_X1    g0587(.A(G294), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n334), .B1(new_n730), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G303), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n722), .A2(new_n790), .B1(new_n725), .B2(new_n791), .ZN(new_n792));
  NOR4_X1   g0592(.A1(new_n787), .A2(new_n737), .A3(new_n789), .A4(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n712), .B1(new_n785), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n712), .A2(new_n713), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT98), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n794), .B(new_n719), .C1(G77), .C2(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n426), .B1(new_n414), .B2(new_n632), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n424), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n424), .A2(new_n642), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n797), .B1(new_n713), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n802), .B1(new_n623), .B2(new_n642), .ZN(new_n804));
  INV_X1    g0604(.A(new_n802), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n622), .A2(new_n632), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n719), .B1(new_n807), .B2(new_n688), .ZN(new_n808));
  INV_X1    g0608(.A(new_n688), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n804), .A2(new_n809), .A3(new_n806), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n803), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(G384));
  NOR2_X1   g0612(.A1(new_n626), .A2(new_n250), .ZN(new_n813));
  INV_X1    g0613(.A(new_n428), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n809), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT103), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(new_n365), .B2(new_n631), .ZN(new_n817));
  AOI211_X1 g0617(.A(KEYINPUT103), .B(new_n630), .C1(new_n347), .C2(new_n352), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n368), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT37), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n817), .A2(new_n818), .ZN(new_n822));
  INV_X1    g0622(.A(new_n353), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(new_n363), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n821), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n365), .A2(new_n366), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n353), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n819), .A2(KEYINPUT37), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n820), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT104), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT38), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(KEYINPUT37), .B1(new_n819), .B2(new_n827), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n824), .B(new_n821), .C1(new_n818), .C2(new_n817), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n833), .A2(new_n834), .B1(new_n368), .B2(new_n819), .ZN(new_n835));
  OAI21_X1  g0635(.A(KEYINPUT104), .B1(new_n835), .B2(KEYINPUT38), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT101), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n342), .A2(new_n285), .ZN(new_n838));
  AOI21_X1  g0638(.A(KEYINPUT7), .B1(new_n704), .B2(new_n223), .ZN(new_n839));
  OAI21_X1  g0639(.A(G68), .B1(new_n839), .B2(new_n336), .ZN(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT16), .B1(new_n840), .B2(new_n333), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n837), .B(new_n352), .C1(new_n838), .C2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n352), .B1(new_n838), .B2(new_n841), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(KEYINPUT101), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n368), .A2(new_n631), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n362), .A2(new_n630), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n844), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n821), .B1(new_n847), .B2(new_n353), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT102), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n834), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI211_X1 g0650(.A(KEYINPUT102), .B(new_n821), .C1(new_n847), .C2(new_n353), .ZN(new_n851));
  OAI211_X1 g0651(.A(KEYINPUT38), .B(new_n845), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n832), .A2(new_n836), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n395), .A2(new_n632), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n854), .B(new_n397), .C1(new_n403), .C2(new_n404), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n403), .A2(new_n404), .A3(new_n642), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n805), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n594), .A2(new_n507), .A3(new_n642), .ZN(new_n859));
  INV_X1    g0659(.A(new_n685), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n687), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n853), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n854), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n405), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n802), .B1(new_n865), .B2(new_n856), .ZN(new_n866));
  INV_X1    g0666(.A(new_n687), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n674), .B2(new_n685), .ZN(new_n868));
  OR2_X1    g0668(.A1(KEYINPUT106), .A2(KEYINPUT40), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT106), .B1(new_n866), .B2(new_n868), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n845), .B1(new_n850), .B2(new_n851), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n831), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n852), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n863), .A2(KEYINPUT40), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(G330), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n815), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n814), .A2(new_n868), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n878), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n669), .A2(new_n814), .A3(new_n671), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n606), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n880), .B(new_n882), .Z(new_n883));
  NOR2_X1   g0683(.A1(new_n855), .A2(new_n857), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n806), .B2(new_n801), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n875), .A2(new_n885), .B1(new_n596), .B2(new_n630), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT105), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n832), .A2(new_n836), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT39), .B1(new_n889), .B2(new_n875), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n888), .A2(KEYINPUT39), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n853), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n403), .A2(new_n404), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n894), .A2(new_n642), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n887), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n813), .B1(new_n883), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n896), .B2(new_n883), .ZN(new_n898));
  OAI211_X1 g0698(.A(G116), .B(new_n224), .C1(new_n579), .C2(KEYINPUT35), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(KEYINPUT35), .B2(new_n579), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n900), .B(KEYINPUT36), .Z(new_n901));
  NOR3_X1   g0701(.A1(new_n228), .A2(new_n262), .A3(new_n329), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n287), .B2(G68), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n625), .A2(G1), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n898), .B(new_n901), .C1(new_n903), .C2(new_n904), .ZN(G367));
  INV_X1    g0705(.A(new_n706), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n240), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n716), .B1(new_n219), .B2(new_n524), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n719), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(G317), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n746), .A2(new_n454), .B1(new_n739), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n747), .A2(new_n696), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT46), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n911), .B(new_n913), .C1(G283), .C2(new_n780), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n722), .A2(new_n762), .B1(new_n725), .B2(new_n788), .ZN(new_n915));
  AOI211_X1 g0715(.A(new_n915), .B(new_n705), .C1(G107), .C2(new_n735), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n914), .B(new_n916), .C1(new_n790), .C2(new_n731), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n746), .A2(new_n262), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n918), .A2(new_n334), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n919), .B(KEYINPUT107), .Z(new_n920));
  NOR2_X1   g0720(.A1(new_n736), .A2(new_n203), .ZN(new_n921));
  OAI22_X1  g0721(.A1(new_n722), .A2(new_n782), .B1(new_n725), .B2(new_n742), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n202), .A2(new_n747), .B1(new_n730), .B2(new_n292), .ZN(new_n923));
  INV_X1    g0723(.A(G137), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n729), .A2(new_n287), .B1(new_n739), .B2(new_n924), .ZN(new_n925));
  NOR4_X1   g0725(.A1(new_n921), .A2(new_n922), .A3(new_n923), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n920), .A2(new_n926), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n927), .A2(KEYINPUT108), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(KEYINPUT108), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n917), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT47), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n767), .B1(new_n930), .B2(new_n931), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n909), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n769), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n642), .A2(new_n526), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n615), .A2(new_n936), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n543), .A2(new_n936), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n934), .B1(new_n935), .B2(new_n939), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n650), .B(new_n647), .Z(new_n941));
  XNOR2_X1  g0741(.A(new_n641), .B(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n690), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n607), .B1(new_n560), .B2(new_n632), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n617), .A2(new_n642), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n651), .A2(new_n644), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT44), .Z(new_n951));
  NOR2_X1   g0751(.A1(new_n948), .A2(new_n949), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT45), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n951), .A2(new_n649), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(new_n953), .ZN(new_n955));
  INV_X1    g0755(.A(new_n649), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n944), .A2(new_n954), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n690), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n654), .B(KEYINPUT41), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n718), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n651), .A2(new_n945), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n962), .A2(KEYINPUT42), .B1(new_n617), .B2(new_n632), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n945), .B1(KEYINPUT42), .B2(new_n644), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n949), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n963), .A2(new_n965), .B1(KEYINPUT43), .B2(new_n939), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n649), .A2(new_n948), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n968), .B(new_n969), .Z(new_n970));
  OAI21_X1  g0770(.A(new_n940), .B1(new_n961), .B2(new_n970), .ZN(G387));
  INV_X1    g0771(.A(new_n656), .ZN(new_n972));
  AOI211_X1 g0772(.A(G45), .B(new_n972), .C1(G68), .C2(G77), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(KEYINPUT110), .ZN(new_n975));
  OAI21_X1  g0775(.A(KEYINPUT50), .B1(new_n290), .B2(G50), .ZN(new_n976));
  OR3_X1    g0776(.A1(new_n290), .A2(KEYINPUT50), .A3(G50), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT110), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n976), .B(new_n977), .C1(new_n973), .C2(new_n978), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n706), .B1(new_n432), .B2(new_n235), .C1(new_n975), .C2(new_n979), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n695), .A2(new_n972), .B1(new_n416), .B2(new_n653), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT109), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n716), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n719), .B(new_n984), .C1(new_n648), .C2(new_n935), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G68), .A2(new_n780), .B1(new_n750), .B2(G97), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n287), .B2(new_n730), .C1(new_n290), .C2(new_n725), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G159), .A2(new_n723), .B1(new_n755), .B2(G77), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n292), .B2(new_n739), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n736), .A2(new_n524), .ZN(new_n990));
  NOR4_X1   g0790(.A1(new_n987), .A2(new_n989), .A3(new_n704), .A4(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT111), .Z(new_n992));
  AOI22_X1  g0792(.A1(G116), .A2(new_n750), .B1(new_n740), .B2(G326), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n731), .A2(new_n910), .B1(new_n790), .B2(new_n729), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT113), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n762), .B2(new_n725), .C1(new_n752), .C2(new_n722), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT48), .Z(new_n997));
  AOI22_X1  g0797(.A1(new_n755), .A2(G294), .B1(new_n735), .B2(G283), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT112), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n704), .B(new_n993), .C1(new_n1000), .C2(KEYINPUT49), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n1000), .A2(KEYINPUT49), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n992), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT114), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n767), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n985), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(new_n942), .B2(new_n718), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n690), .A2(new_n942), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n943), .A2(new_n654), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1008), .B1(new_n1009), .B2(new_n1010), .ZN(G393));
  INV_X1    g0811(.A(KEYINPUT115), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n957), .A2(new_n1012), .A3(new_n954), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n955), .A2(KEYINPUT115), .A3(new_n956), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n958), .B(new_n654), .C1(new_n944), .C2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n948), .A2(new_n715), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n716), .B1(new_n454), .B2(new_n219), .C1(new_n906), .C2(new_n247), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n719), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G68), .A2(new_n755), .B1(new_n750), .B2(G87), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n735), .A2(G77), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1020), .A2(new_n705), .A3(new_n1021), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n722), .A2(new_n292), .B1(new_n730), .B2(new_n742), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT51), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n780), .A2(new_n350), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G50), .A2(new_n726), .B1(new_n740), .B2(G143), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n722), .A2(new_n910), .B1(new_n730), .B2(new_n762), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT52), .Z(new_n1031));
  AOI22_X1  g0831(.A1(G283), .A2(new_n755), .B1(new_n726), .B2(G303), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G294), .A2(new_n780), .B1(new_n740), .B2(G322), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n735), .A2(G116), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n259), .B1(new_n750), .B2(G107), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n1022), .A2(new_n1029), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1019), .B1(new_n1037), .B2(new_n712), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1015), .A2(new_n718), .B1(new_n1017), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1016), .A2(new_n1039), .ZN(G390));
  NAND4_X1  g0840(.A1(new_n686), .A2(G330), .A3(new_n687), .A4(new_n805), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n884), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT117), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT116), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n688), .B2(new_n858), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n866), .A2(new_n868), .A3(KEYINPUT116), .A4(G330), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1041), .A2(KEYINPUT117), .A3(new_n884), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1044), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n806), .A2(new_n801), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n809), .A2(new_n866), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n632), .B(new_n799), .C1(new_n663), .C2(new_n665), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1054), .A2(new_n801), .ZN(new_n1055));
  AND3_X1   g0855(.A1(new_n1053), .A2(new_n1055), .A3(new_n1042), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1052), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n881), .A2(new_n606), .A3(new_n815), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(KEYINPUT118), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1056), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT118), .ZN(new_n1063));
  NOR3_X1   g0863(.A1(new_n1062), .A2(new_n1059), .A3(new_n1063), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n885), .A2(new_n895), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n890), .A2(new_n892), .A3(new_n1065), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n853), .B1(new_n894), .B2(new_n642), .C1(new_n1055), .C2(new_n884), .ZN(new_n1067));
  AND3_X1   g0867(.A1(new_n1066), .A2(new_n1067), .A3(new_n1053), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n1061), .A2(new_n1064), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1066), .A2(new_n1067), .A3(new_n1053), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1062), .A2(new_n1059), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1073), .B(new_n1074), .C1(new_n1075), .C2(new_n1070), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1072), .A2(new_n654), .A3(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n890), .A2(new_n713), .A3(new_n892), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n719), .B1(new_n796), .B2(new_n350), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n747), .A2(new_n292), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT53), .ZN(new_n1082));
  XOR2_X1   g0882(.A(KEYINPUT54), .B(G143), .Z(new_n1083));
  AOI22_X1  g0883(.A1(new_n780), .A2(new_n1083), .B1(new_n750), .B2(G50), .ZN(new_n1084));
  INV_X1    g0884(.A(G128), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1082), .B(new_n1084), .C1(new_n1085), .C2(new_n722), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n730), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(G132), .A2(new_n1087), .B1(new_n726), .B2(G137), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n334), .B1(new_n740), .B2(G125), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1088), .B(new_n1089), .C1(new_n742), .C2(new_n736), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G283), .A2(new_n723), .B1(new_n780), .B2(G97), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1091), .B1(new_n416), .B2(new_n725), .C1(new_n696), .C2(new_n730), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n259), .B1(new_n755), .B2(G87), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n740), .A2(G294), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1093), .A2(new_n1094), .A3(new_n775), .A4(new_n1021), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n1086), .A2(new_n1090), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1080), .B1(new_n1096), .B2(new_n712), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1078), .A2(new_n718), .B1(new_n1079), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1077), .A2(new_n1098), .ZN(G378));
  INV_X1    g0899(.A(KEYINPUT123), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n298), .A2(new_n630), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n308), .A2(KEYINPUT121), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n308), .A2(KEYINPUT121), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1101), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1104), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1101), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1106), .A2(new_n1107), .A3(new_n1102), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1105), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n876), .B2(new_n877), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n872), .A2(new_n875), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT40), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n853), .B2(new_n862), .ZN(new_n1120));
  OAI211_X1 g0920(.A(G330), .B(new_n1116), .C1(new_n1118), .C2(new_n1120), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n896), .A2(new_n1115), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n893), .A2(new_n895), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1115), .A2(new_n1121), .B1(new_n1123), .B2(new_n886), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1100), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1115), .A2(new_n1121), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1123), .A2(new_n886), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n896), .A2(new_n1115), .A3(new_n1121), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1128), .A2(KEYINPUT123), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1076), .A2(new_n1060), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1125), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT57), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1059), .B1(new_n1078), .B2(new_n1058), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1128), .A2(KEYINPUT57), .A3(new_n1129), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n654), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1125), .A2(new_n718), .A3(new_n1130), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n1085), .A2(new_n730), .B1(new_n725), .B2(new_n773), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n723), .A2(G125), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1083), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1142), .B1(new_n924), .B2(new_n729), .C1(new_n747), .C2(new_n1143), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1141), .B(new_n1144), .C1(G150), .C2(new_n735), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT59), .ZN(new_n1146));
  OR2_X1    g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n750), .A2(G159), .ZN(new_n1149));
  AOI211_X1 g0949(.A(G33), .B(G41), .C1(new_n740), .C2(G124), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n921), .B1(G116), .B2(new_n723), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT119), .Z(new_n1153));
  NOR2_X1   g0953(.A1(new_n705), .A2(G41), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(G77), .A2(new_n755), .B1(new_n740), .B2(G283), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G97), .A2(new_n726), .B1(new_n780), .B2(new_n410), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G107), .A2(new_n1087), .B1(new_n750), .B2(G58), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1153), .A2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g0959(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1151), .A2(new_n1161), .ZN(new_n1162));
  AOI211_X1 g0962(.A(G50), .B(new_n1154), .C1(new_n309), .C2(new_n429), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n719), .B1(G50), .B2(new_n796), .C1(new_n1165), .C2(new_n767), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n1116), .B2(new_n713), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT122), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1140), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1139), .A2(new_n1170), .ZN(G375));
  NAND2_X1  g0971(.A1(new_n1062), .A2(new_n1059), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n960), .B(new_n1172), .C1(new_n1061), .C2(new_n1064), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n731), .A2(new_n924), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n722), .A2(new_n773), .B1(new_n739), .B2(new_n1085), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n1143), .A2(new_n725), .B1(new_n742), .B2(new_n747), .ZN(new_n1176));
  NOR3_X1   g0976(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n202), .A2(new_n746), .B1(new_n729), .B2(new_n292), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n704), .B(new_n1178), .C1(G50), .C2(new_n735), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n722), .A2(new_n788), .B1(new_n725), .B2(new_n696), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n730), .A2(new_n791), .B1(new_n739), .B2(new_n790), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n747), .A2(new_n454), .B1(new_n729), .B2(new_n416), .ZN(new_n1183));
  NOR4_X1   g0983(.A1(new_n990), .A2(new_n1183), .A3(new_n259), .A4(new_n918), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1177), .A2(new_n1179), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n719), .B1(G68), .B2(new_n796), .C1(new_n1185), .C2(new_n767), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1186), .B(KEYINPUT124), .Z(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n884), .B2(new_n713), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n1058), .B2(new_n718), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1173), .A2(new_n1189), .ZN(G381));
  NOR2_X1   g0990(.A1(G375), .A2(G378), .ZN(new_n1191));
  OR2_X1    g0991(.A1(G393), .A2(G396), .ZN(new_n1192));
  NOR4_X1   g0992(.A1(G387), .A2(G390), .A3(G384), .A4(new_n1192), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1191), .A2(new_n1189), .A3(new_n1173), .A4(new_n1193), .ZN(G407));
  INV_X1    g0994(.A(G343), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(G213), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT125), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1191), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(G407), .A2(new_n1198), .A3(G213), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT126), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1199), .B(new_n1200), .ZN(G409));
  NAND3_X1  g1001(.A1(G387), .A2(new_n1016), .A3(new_n1039), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(G393), .B(new_n771), .ZN(new_n1203));
  OAI211_X1 g1003(.A(G390), .B(new_n940), .C1(new_n961), .C2(new_n970), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1203), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1074), .A2(new_n655), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1062), .A2(KEYINPUT60), .A3(new_n1059), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT60), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1172), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1209), .A2(new_n1210), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n1189), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n811), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1214), .A2(new_n811), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1128), .A2(new_n718), .A3(new_n1129), .ZN(new_n1219));
  AND4_X1   g1019(.A1(new_n1077), .A2(new_n1098), .A3(new_n1168), .A4(new_n1219), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1125), .A2(new_n1131), .A3(new_n1130), .A4(new_n960), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1197), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1169), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1223));
  INV_X1    g1023(.A(G378), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1218), .B(new_n1222), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(KEYINPUT127), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT62), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1137), .B1(new_n1133), .B2(new_n1132), .ZN(new_n1228));
  OAI21_X1  g1028(.A(G378), .B1(new_n1228), .B2(new_n1169), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT127), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1229), .A2(new_n1230), .A3(new_n1218), .A4(new_n1222), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1226), .A2(new_n1227), .A3(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1222), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1197), .A2(G2897), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1217), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1237), .A2(new_n1215), .A3(new_n1234), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1236), .A2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT61), .B1(new_n1233), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1225), .A2(KEYINPUT62), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1208), .B1(new_n1232), .B2(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1229), .A2(KEYINPUT63), .A3(new_n1218), .A4(new_n1222), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1240), .A2(new_n1244), .A3(new_n1207), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1226), .A2(new_n1231), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT63), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1245), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1243), .A2(new_n1249), .ZN(G405));
  NAND2_X1  g1050(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1229), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n1252), .A2(new_n1218), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1218), .ZN(new_n1254));
  AND3_X1   g1054(.A1(new_n1253), .A2(new_n1207), .A3(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1207), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1255), .A2(new_n1256), .ZN(G402));
endmodule


