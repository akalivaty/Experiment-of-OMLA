//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT76), .B(G902), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT83), .A3(G104), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT3), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n198), .A2(new_n195), .A3(KEYINPUT83), .A4(G104), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n195), .A2(G104), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n197), .A2(new_n199), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G101), .ZN(new_n203));
  INV_X1    g017(.A(G101), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n197), .A2(new_n201), .A3(new_n204), .A4(new_n199), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(KEYINPUT4), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT4), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n202), .A2(new_n207), .A3(G101), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  AND2_X1   g025(.A1(KEYINPUT64), .A2(G146), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT64), .A2(G146), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n211), .B1(new_n214), .B2(G143), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n215), .A2(KEYINPUT65), .A3(KEYINPUT0), .A4(G128), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(new_n210), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT64), .A2(G146), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(G143), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n211), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n220), .A2(KEYINPUT0), .A3(G128), .A4(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n210), .A2(G143), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n225), .B1(new_n214), .B2(G143), .ZN(new_n226));
  XOR2_X1   g040(.A(KEYINPUT0), .B(G128), .Z(new_n227));
  AOI22_X1  g041(.A1(new_n216), .A2(new_n224), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G104), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(G107), .ZN(new_n230));
  OAI21_X1  g044(.A(G101), .B1(new_n230), .B2(new_n200), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n205), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT1), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n220), .A2(new_n233), .A3(G128), .A4(new_n221), .ZN(new_n234));
  INV_X1    g048(.A(G143), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT1), .B1(new_n235), .B2(G146), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n220), .A2(new_n221), .B1(G128), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n234), .B1(new_n237), .B2(KEYINPUT84), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT84), .ZN(new_n239));
  INV_X1    g053(.A(G128), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(new_n225), .B2(KEYINPUT1), .ZN(new_n241));
  NOR3_X1   g055(.A1(new_n215), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n232), .B1(new_n238), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT10), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n209), .A2(new_n228), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n240), .B1(new_n220), .B2(KEYINPUT1), .ZN(new_n246));
  INV_X1    g060(.A(new_n225), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n218), .A2(new_n219), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n247), .B1(new_n248), .B2(new_n235), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT71), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT71), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n233), .B1(new_n214), .B2(G143), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n251), .B(new_n226), .C1(new_n252), .C2(new_n240), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n253), .A3(new_n234), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n205), .A2(new_n231), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(new_n244), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n245), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G134), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT11), .B1(new_n259), .B2(G137), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT11), .ZN(new_n261));
  INV_X1    g075(.A(G137), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(new_n262), .A3(G134), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G131), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT66), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n266), .B1(new_n262), .B2(G134), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n259), .A2(KEYINPUT66), .A3(G137), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n264), .A2(new_n265), .A3(new_n267), .A4(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT67), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n267), .A2(new_n268), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n272), .A2(KEYINPUT67), .A3(new_n265), .A4(new_n264), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n264), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G131), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n258), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n243), .A2(new_n244), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n271), .A2(new_n273), .B1(G131), .B2(new_n275), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n216), .A2(new_n224), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n226), .A2(new_n227), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n281), .A2(new_n282), .A3(new_n206), .A4(new_n208), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n279), .A2(new_n257), .A3(new_n280), .A4(new_n283), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n284), .A2(KEYINPUT85), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n284), .A2(KEYINPUT85), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n278), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G953), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G227), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n289), .B(KEYINPUT82), .ZN(new_n290));
  XNOR2_X1  g104(.A(G110), .B(G140), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n290), .B(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n243), .B1(new_n254), .B2(new_n232), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(KEYINPUT12), .A3(new_n277), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT86), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n294), .A2(new_n277), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT12), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n294), .A2(KEYINPUT86), .A3(KEYINPUT12), .A4(new_n277), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n297), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n292), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT85), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n245), .A2(new_n304), .A3(new_n280), .A4(new_n257), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n284), .A2(KEYINPUT85), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n302), .A2(new_n303), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n194), .B1(new_n293), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n192), .B1(new_n309), .B2(new_n190), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n307), .A2(new_n303), .A3(new_n278), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n302), .A2(new_n307), .ZN(new_n312));
  OAI211_X1 g126(.A(G469), .B(new_n311), .C1(new_n312), .C2(new_n303), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n189), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(G210), .B1(G237), .B2(G902), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT90), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n253), .A2(new_n234), .ZN(new_n318));
  INV_X1    g132(.A(G125), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n318), .A2(KEYINPUT88), .A3(new_n319), .A4(new_n250), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n250), .A2(new_n253), .A3(new_n319), .A4(new_n234), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT88), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G224), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(G953), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT87), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n328), .B1(new_n228), .B2(new_n319), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n222), .A2(new_n223), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n222), .A2(new_n223), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n282), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(KEYINPUT87), .A3(G125), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n324), .A2(new_n327), .A3(new_n329), .A4(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT7), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G119), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT73), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT73), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G119), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n340), .A3(G116), .ZN(new_n341));
  INV_X1    g155(.A(G116), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G119), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT2), .B(G113), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n345), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(new_n341), .A3(new_n343), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n206), .A2(new_n349), .A3(new_n208), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n341), .A2(KEYINPUT5), .A3(new_n343), .ZN(new_n351));
  OAI21_X1  g165(.A(G113), .B1(new_n341), .B2(KEYINPUT5), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n232), .B(new_n348), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(G110), .B(G122), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n354), .B(KEYINPUT8), .ZN(new_n356));
  INV_X1    g170(.A(new_n353), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n348), .B1(new_n351), .B2(new_n352), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n358), .A2(new_n255), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n356), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n320), .A2(new_n323), .B1(G125), .B2(new_n332), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n326), .A2(new_n335), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n355), .B(new_n360), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n317), .B(new_n191), .C1(new_n336), .C2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n321), .B(KEYINPUT88), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n329), .A2(new_n333), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n326), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n334), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT89), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n355), .A2(KEYINPUT6), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n354), .B1(new_n350), .B2(new_n353), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI211_X1 g186(.A(KEYINPUT6), .B(new_n354), .C1(new_n350), .C2(new_n353), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n368), .A2(new_n369), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n369), .B1(new_n368), .B2(new_n374), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n364), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n191), .B1(new_n336), .B2(new_n363), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n378), .A2(KEYINPUT90), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n316), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n368), .A2(new_n374), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT89), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n368), .A2(new_n374), .A3(new_n369), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n378), .A2(KEYINPUT90), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n384), .A2(new_n315), .A3(new_n385), .A4(new_n364), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(G214), .B1(G237), .B2(G902), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n314), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n235), .A2(G128), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT94), .B1(new_n391), .B2(KEYINPUT13), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n240), .A2(G143), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT94), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT13), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n390), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n392), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n397), .A2(KEYINPUT95), .B1(KEYINPUT13), .B2(new_n391), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT95), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n392), .A2(new_n399), .A3(new_n393), .A4(new_n396), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n259), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  OR2_X1    g215(.A1(new_n342), .A2(G122), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n342), .A2(G122), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n195), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n390), .A2(new_n393), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n259), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n403), .A3(G107), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n405), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n401), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n406), .B(G134), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT96), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n411), .A2(KEYINPUT96), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n195), .B1(new_n402), .B2(KEYINPUT14), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(new_n404), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n413), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G217), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n187), .A2(new_n418), .A3(G953), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n410), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT97), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OR2_X1    g237(.A1(new_n414), .A2(new_n416), .ZN(new_n424));
  OAI221_X1 g238(.A(new_n419), .B1(new_n401), .B2(new_n409), .C1(new_n424), .C2(new_n413), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT97), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n420), .B1(new_n410), .B2(new_n417), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n423), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n193), .ZN(new_n429));
  INV_X1    g243(.A(G478), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(KEYINPUT15), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n429), .B(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G237), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT75), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT75), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(G237), .ZN(new_n438));
  AOI21_X1  g252(.A(G953), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(G143), .A3(G214), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(G143), .B1(new_n439), .B2(G214), .ZN(new_n442));
  OAI211_X1 g256(.A(KEYINPUT18), .B(G131), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G125), .B(G140), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n214), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(new_n210), .B2(new_n444), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n439), .A2(G214), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n235), .ZN(new_n448));
  NAND2_X1  g262(.A1(KEYINPUT18), .A2(G131), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n440), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n443), .A2(new_n446), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G131), .B1(new_n441), .B2(new_n442), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n448), .A2(new_n265), .A3(new_n440), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(KEYINPUT17), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT78), .ZN(new_n456));
  INV_X1    g270(.A(G140), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G125), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n456), .B1(new_n458), .B2(KEYINPUT16), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n319), .A2(KEYINPUT16), .A3(G140), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n460), .B1(new_n444), .B2(KEYINPUT16), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n459), .B1(new_n461), .B2(new_n456), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n210), .ZN(new_n463));
  OAI211_X1 g277(.A(G146), .B(new_n459), .C1(new_n461), .C2(new_n456), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT17), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n463), .B(new_n464), .C1(new_n452), .C2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n451), .B1(new_n455), .B2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(G113), .B(G122), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(new_n229), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n469), .B(new_n451), .C1(new_n455), .C2(new_n466), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n191), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G475), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT93), .ZN(new_n476));
  INV_X1    g290(.A(new_n451), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n319), .A2(G140), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n458), .A2(new_n478), .A3(KEYINPUT19), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT19), .B1(new_n458), .B2(new_n478), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n214), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT92), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT92), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n483), .B(new_n214), .C1(new_n479), .C2(new_n480), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n464), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n485), .B1(new_n454), .B2(KEYINPUT91), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT91), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n452), .A2(new_n453), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n477), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n476), .B1(new_n489), .B2(new_n469), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n454), .A2(KEYINPUT91), .ZN(new_n491));
  INV_X1    g305(.A(new_n485), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n451), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(KEYINPUT93), .A3(new_n470), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n490), .A2(new_n495), .A3(new_n472), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT20), .ZN(new_n497));
  NOR2_X1   g311(.A1(G475), .A2(G902), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n497), .B1(new_n496), .B2(new_n498), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n475), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(G234), .A2(G237), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(G952), .A3(new_n288), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n194), .A2(G953), .A3(new_n503), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT21), .B(G898), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n434), .A2(new_n502), .A3(new_n509), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n389), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n463), .A2(new_n464), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT24), .B(G110), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT73), .B(G119), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(G128), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n337), .A2(G128), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n516), .A2(KEYINPUT77), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n514), .A2(KEYINPUT77), .A3(G128), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n513), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G110), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n514), .A2(G128), .B1(KEYINPUT23), .B2(new_n516), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT23), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n514), .B2(G128), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n521), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n512), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n518), .A2(new_n513), .A3(new_n519), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n522), .A2(new_n524), .A3(new_n521), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(new_n464), .A3(new_n445), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT79), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n527), .A2(KEYINPUT79), .A3(new_n531), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT22), .B(G137), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n288), .A2(G221), .A3(G234), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n534), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n532), .A2(new_n533), .A3(new_n538), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n418), .B1(new_n193), .B2(G234), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n543), .A2(G902), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT81), .ZN(new_n546));
  NAND2_X1  g360(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n194), .B1(new_n540), .B2(new_n541), .ZN(new_n548));
  NOR2_X1   g362(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n547), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  AOI211_X1 g365(.A(new_n194), .B(new_n549), .C1(new_n540), .C2(new_n541), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n543), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n546), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n349), .B1(new_n277), .B2(new_n228), .ZN(new_n555));
  OR3_X1    g369(.A1(new_n262), .A2(KEYINPUT69), .A3(G134), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT69), .B1(new_n262), .B2(G134), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n556), .B(new_n557), .C1(new_n259), .C2(G137), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n271), .A2(new_n273), .B1(G131), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n254), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT28), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT74), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n254), .A2(new_n559), .A3(KEYINPUT74), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n565), .A2(new_n566), .A3(new_n555), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT72), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT70), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n254), .B1(new_n559), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n558), .A2(G131), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n274), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n568), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n274), .A2(new_n571), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT70), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n559), .A2(new_n569), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n575), .A2(KEYINPUT72), .A3(new_n576), .A4(new_n254), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT68), .B1(new_n332), .B2(new_n280), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT68), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n277), .A2(new_n579), .A3(new_n228), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n573), .A2(new_n577), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n567), .B1(new_n582), .B2(new_n349), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n563), .B1(new_n583), .B2(new_n562), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n439), .A2(G210), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(KEYINPUT27), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT26), .B(G101), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n277), .A2(new_n228), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n565), .A2(KEYINPUT30), .A3(new_n591), .A4(new_n566), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n349), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT30), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n593), .B1(new_n594), .B2(new_n582), .ZN(new_n595));
  INV_X1    g409(.A(new_n567), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n588), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT31), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n582), .A2(new_n594), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n599), .A2(new_n349), .A3(new_n592), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT31), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n600), .A2(new_n601), .A3(new_n596), .A4(new_n588), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n590), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(G472), .A2(G902), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT32), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT32), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n603), .A2(new_n607), .A3(new_n604), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n584), .A2(new_n588), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n600), .A2(new_n596), .A3(new_n589), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT29), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n565), .A2(new_n566), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n591), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n567), .B1(new_n614), .B2(new_n349), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n563), .B1(new_n615), .B2(new_n562), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n588), .A2(KEYINPUT29), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n193), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(G472), .B1(new_n612), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n554), .B1(new_n609), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n511), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  NAND2_X1  g436(.A1(new_n603), .A2(new_n193), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(G472), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n605), .ZN(new_n625));
  INV_X1    g439(.A(new_n308), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n303), .B1(new_n307), .B2(new_n278), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n190), .B(new_n193), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n192), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(new_n313), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n188), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n625), .A2(new_n554), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n496), .A2(new_n498), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT20), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n634), .A2(new_n499), .B1(G475), .B2(new_n474), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n425), .A2(new_n427), .A3(KEYINPUT33), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT33), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n637), .B1(new_n428), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n194), .A2(new_n430), .ZN(new_n640));
  AOI22_X1  g454(.A1(new_n639), .A2(new_n640), .B1(new_n429), .B2(new_n430), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n509), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n642), .A2(new_n387), .A3(new_n388), .A4(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT98), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n388), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n380), .B2(new_n386), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n648), .A2(KEYINPUT98), .A3(new_n643), .A4(new_n642), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n632), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  NOR2_X1   g466(.A1(new_n502), .A2(new_n433), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n648), .A2(new_n643), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n632), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G107), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT99), .B(KEYINPUT35), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G9));
  INV_X1    g472(.A(new_n625), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n539), .A2(KEYINPUT36), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n532), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n544), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n553), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT100), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT101), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n659), .A2(new_n668), .A3(new_n665), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n667), .A2(new_n511), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  AND3_X1   g486(.A1(new_n603), .A2(new_n607), .A3(new_n604), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n607), .B1(new_n603), .B2(new_n604), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n619), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n434), .A2(new_n635), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n504), .B(KEYINPUT102), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(G900), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n678), .B1(new_n507), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n389), .A2(new_n675), .A3(new_n665), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  XNOR2_X1  g497(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n680), .B(new_n684), .Z(new_n685));
  NOR2_X1   g499(.A1(new_n631), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT40), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n387), .B(KEYINPUT38), .ZN(new_n689));
  INV_X1    g503(.A(new_n663), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n635), .A2(new_n433), .ZN(new_n691));
  AND4_X1   g505(.A1(new_n388), .A2(new_n689), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n615), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n191), .B1(new_n693), .B2(new_n588), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n589), .B1(new_n600), .B2(new_n596), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n696), .B1(new_n673), .B2(new_n674), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT103), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n699), .B(new_n696), .C1(new_n673), .C2(new_n674), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n692), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n688), .B1(new_n702), .B2(KEYINPUT104), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n692), .A2(new_n701), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT104), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G143), .ZN(G45));
  NOR3_X1   g522(.A1(new_n635), .A2(new_n641), .A3(new_n680), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n389), .A2(new_n675), .A3(new_n665), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G146), .ZN(G48));
  OAI21_X1  g525(.A(new_n193), .B1(new_n626), .B2(new_n627), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(G469), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n713), .A2(new_n188), .A3(new_n628), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n620), .A2(new_n646), .A3(new_n649), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT41), .B(G113), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G15));
  INV_X1    g531(.A(KEYINPUT106), .ZN(new_n718));
  INV_X1    g532(.A(new_n554), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n675), .A2(new_n719), .A3(new_n714), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n648), .A2(new_n643), .A3(new_n653), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n718), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n620), .A2(KEYINPUT106), .A3(new_n654), .A4(new_n714), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  AND2_X1   g539(.A1(new_n675), .A2(new_n665), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n510), .A2(new_n648), .A3(new_n714), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G119), .ZN(G21));
  INV_X1    g543(.A(new_n604), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n602), .A2(new_n598), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n616), .A2(new_n589), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n713), .A2(new_n188), .A3(new_n628), .A4(new_n643), .ZN(new_n734));
  XOR2_X1   g548(.A(KEYINPUT107), .B(G472), .Z(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n736), .B1(new_n603), .B2(new_n193), .ZN(new_n737));
  NOR4_X1   g551(.A1(new_n733), .A2(new_n734), .A3(new_n737), .A4(new_n554), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n648), .A2(new_n691), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G122), .ZN(G24));
  AND2_X1   g555(.A1(new_n648), .A2(new_n714), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n733), .A2(new_n737), .A3(new_n690), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n709), .A3(new_n743), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT108), .B(G125), .Z(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G27));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n380), .A2(new_n388), .A3(new_n386), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n631), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n675), .A2(new_n749), .A3(new_n709), .A4(new_n719), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(KEYINPUT109), .A3(KEYINPUT42), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT42), .B1(new_n750), .B2(KEYINPUT109), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n747), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n753), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(KEYINPUT110), .A3(new_n751), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G131), .ZN(G33));
  NAND2_X1  g572(.A1(new_n675), .A2(new_n719), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n759), .A2(new_n631), .A3(new_n748), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n681), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G134), .ZN(G36));
  NOR2_X1   g576(.A1(new_n502), .A2(new_n641), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(KEYINPUT43), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n625), .A3(new_n663), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n748), .B1(new_n765), .B2(new_n766), .ZN(new_n768));
  INV_X1    g582(.A(new_n685), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n311), .B1(new_n312), .B2(new_n303), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n190), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n772), .B1(new_n771), .B2(new_n770), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT46), .B1(new_n773), .B2(new_n629), .ZN(new_n774));
  INV_X1    g588(.A(new_n628), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(KEYINPUT46), .A3(new_n629), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n189), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n767), .A2(new_n768), .A3(new_n769), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  XNOR2_X1  g594(.A(new_n778), .B(KEYINPUT47), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n709), .A2(new_n554), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n675), .A2(new_n782), .A3(new_n748), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  AND3_X1   g599(.A1(new_n682), .A2(new_n710), .A3(new_n744), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n663), .A2(new_n680), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n648), .A2(new_n314), .A3(new_n691), .A4(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT113), .B1(new_n701), .B2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n791));
  AOI211_X1 g605(.A(new_n791), .B(new_n788), .C1(new_n698), .C2(new_n700), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n786), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n786), .B(KEYINPUT52), .C1(new_n790), .C2(new_n792), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(KEYINPUT114), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n632), .A2(new_n648), .A3(new_n643), .A4(new_n642), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n670), .A2(new_n621), .A3(new_n655), .A4(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT111), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n722), .A2(new_n723), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n715), .A2(new_n728), .A3(new_n740), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n726), .A2(new_n727), .B1(new_n738), .B2(new_n739), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n724), .A2(KEYINPUT111), .A3(new_n715), .A4(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n799), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n743), .A2(new_n709), .ZN(new_n807));
  INV_X1    g621(.A(new_n680), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n635), .A2(new_n433), .A3(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT112), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n675), .A2(new_n665), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n807), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n749), .A2(new_n812), .B1(new_n760), .B2(new_n681), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n754), .A2(new_n756), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n793), .A2(new_n815), .A3(new_n794), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n797), .A2(new_n806), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(KEYINPUT115), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n795), .A2(new_n796), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n806), .A2(new_n820), .A3(new_n814), .A4(KEYINPUT53), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT115), .B1(new_n817), .B2(new_n818), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT54), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n806), .A2(new_n820), .A3(new_n814), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n818), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n801), .A2(new_n802), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n752), .A2(new_n753), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n827), .A2(KEYINPUT116), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n724), .A2(new_n715), .A3(new_n804), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n755), .A2(new_n751), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n813), .A2(KEYINPUT53), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n799), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n834), .A2(new_n816), .A3(new_n797), .A4(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n826), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n824), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n713), .A2(new_n628), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NOR4_X1   g657(.A1(new_n689), .A2(new_n388), .A3(new_n189), .A4(new_n843), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n733), .A2(new_n737), .A3(new_n554), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n764), .A2(new_n678), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT50), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n843), .A2(new_n748), .A3(new_n189), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n849), .A2(new_n719), .A3(new_n505), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n850), .A2(new_n701), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(new_n635), .A3(new_n641), .ZN(new_n852));
  INV_X1    g666(.A(new_n743), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n764), .A2(new_n849), .A3(new_n678), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n848), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n748), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n846), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n781), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n843), .A2(new_n188), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n781), .B2(new_n859), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n858), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n841), .B1(new_n856), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n851), .A2(new_n642), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n288), .A2(G952), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n866), .B1(new_n846), .B2(new_n742), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n854), .A2(new_n759), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n868), .A2(KEYINPUT48), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(KEYINPUT48), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n865), .B(new_n867), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n848), .A2(new_n855), .A3(new_n841), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n857), .B(new_n846), .C1(new_n781), .C2(new_n861), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n864), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT118), .ZN(new_n876));
  OAI22_X1  g690(.A1(new_n840), .A2(new_n876), .B1(G952), .B2(G953), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n554), .A2(new_n647), .A3(new_n189), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT49), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n878), .B(new_n763), .C1(new_n879), .C2(new_n842), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n843), .A2(KEYINPUT49), .ZN(new_n881));
  OR3_X1    g695(.A1(new_n689), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n877), .B1(new_n701), .B2(new_n882), .ZN(G75));
  NOR2_X1   g697(.A1(new_n288), .A2(G952), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n193), .B1(new_n826), .B2(new_n837), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n316), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n368), .B(new_n374), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT55), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n890), .A2(KEYINPUT56), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n885), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT56), .B1(new_n887), .B2(KEYINPUT119), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(KEYINPUT119), .B2(new_n887), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n892), .B1(new_n894), .B2(new_n890), .ZN(G51));
  NOR2_X1   g709(.A1(new_n626), .A2(new_n627), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT121), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n826), .A2(new_n837), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT54), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n839), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  XNOR2_X1  g715(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n629), .B(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n897), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n886), .B(new_n772), .C1(new_n771), .C2(new_n770), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n884), .B1(new_n904), .B2(new_n905), .ZN(G54));
  AND2_X1   g720(.A1(KEYINPUT58), .A2(G475), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n886), .A2(new_n496), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n496), .B1(new_n886), .B2(new_n907), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n908), .A2(new_n909), .A3(new_n884), .ZN(G60));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n639), .B(KEYINPUT122), .ZN(new_n912));
  NAND2_X1  g726(.A1(G478), .A2(G902), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT59), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n911), .B1(new_n900), .B2(new_n915), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n826), .A2(new_n838), .A3(new_n837), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n838), .B1(new_n826), .B2(new_n837), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n911), .B(new_n915), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n885), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n912), .B1(new_n840), .B2(new_n914), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n921), .A2(new_n922), .ZN(G63));
  NAND2_X1  g737(.A1(G217), .A2(G902), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT60), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n826), .B2(new_n837), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n926), .A2(new_n542), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n884), .B1(new_n926), .B2(new_n661), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT124), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n929), .A2(KEYINPUT61), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n931));
  AOI211_X1 g745(.A(KEYINPUT124), .B(new_n931), .C1(new_n927), .C2(new_n928), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n930), .A2(new_n932), .ZN(G66));
  OAI21_X1  g747(.A(G953), .B1(new_n508), .B2(new_n325), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(new_n806), .B2(G953), .ZN(new_n935));
  OAI22_X1  g749(.A1(new_n372), .A2(new_n373), .B1(G898), .B2(new_n288), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n935), .B(new_n936), .ZN(G69));
  AOI21_X1  g751(.A(new_n288), .B1(G227), .B2(G900), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT127), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n778), .A2(new_n620), .A3(new_n769), .A4(new_n739), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n940), .A2(new_n761), .A3(new_n786), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n757), .A2(new_n779), .A3(new_n784), .A4(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(G953), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n599), .A2(new_n592), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n479), .A2(new_n480), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n679), .A2(new_n288), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n943), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n676), .B1(new_n635), .B2(new_n641), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n620), .A2(new_n686), .A3(new_n857), .A4(new_n949), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n784), .A2(new_n779), .A3(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n786), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n703), .B2(new_n706), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT62), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n706), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n687), .B1(new_n704), .B2(new_n705), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n954), .B(new_n786), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(KEYINPUT125), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT125), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n953), .A2(new_n960), .A3(new_n954), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n955), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n946), .B1(new_n962), .B2(G953), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n948), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI211_X1 g779(.A(KEYINPUT126), .B(new_n946), .C1(new_n962), .C2(G953), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n939), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n961), .A2(new_n959), .ZN(new_n968));
  INV_X1    g782(.A(new_n955), .ZN(new_n969));
  AOI21_X1  g783(.A(G953), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n946), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n964), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n948), .ZN(new_n973));
  AND4_X1   g787(.A1(new_n939), .A2(new_n972), .A3(new_n966), .A4(new_n973), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n967), .A2(new_n974), .ZN(G72));
  NAND2_X1  g789(.A1(G472), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT63), .Z(new_n977));
  INV_X1    g791(.A(new_n806), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n977), .B1(new_n942), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n611), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n884), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n977), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n982), .B1(new_n962), .B2(new_n806), .ZN(new_n983));
  INV_X1    g797(.A(new_n695), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n981), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n822), .A2(new_n823), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n980), .A2(new_n695), .A3(new_n982), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(G57));
endmodule


