//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT65), .A3(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(G143), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G143), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n191), .B(new_n194), .C1(new_n195), .C2(new_n190), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n190), .A2(G143), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n200), .B1(new_n195), .B2(new_n190), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n197), .B1(new_n192), .B2(KEYINPUT1), .ZN(new_n202));
  OAI22_X1  g016(.A1(new_n196), .A2(new_n199), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  OR2_X1    g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n206), .B(new_n207), .C1(new_n213), .C2(new_n200), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(G146), .ZN(new_n215));
  INV_X1    g029(.A(new_n206), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n215), .A2(new_n191), .A3(new_n194), .A4(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n205), .B1(new_n218), .B2(new_n204), .ZN(new_n219));
  INV_X1    g033(.A(G953), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G224), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n219), .B1(KEYINPUT7), .B2(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT71), .A2(G116), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT71), .A2(G116), .ZN(new_n224));
  OAI21_X1  g038(.A(G119), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G119), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G116), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(KEYINPUT5), .A3(new_n227), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n228), .B(G113), .C1(KEYINPUT5), .C2(new_n227), .ZN(new_n229));
  INV_X1    g043(.A(G113), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT2), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT2), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G113), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n225), .A2(new_n234), .A3(new_n227), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n229), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G104), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G107), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n237), .A2(G107), .ZN(new_n240));
  OAI21_X1  g054(.A(G101), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT3), .B1(new_n237), .B2(G107), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n243));
  INV_X1    g057(.A(G107), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(new_n244), .A3(G104), .ZN(new_n245));
  INV_X1    g059(.A(G101), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n242), .A2(new_n245), .A3(new_n246), .A4(new_n238), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n241), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n236), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n248), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n229), .A2(new_n235), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  XOR2_X1   g066(.A(G110), .B(G122), .Z(new_n253));
  XOR2_X1   g067(.A(new_n253), .B(KEYINPUT8), .Z(new_n254));
  AND2_X1   g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n219), .A2(KEYINPUT7), .A3(new_n221), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n242), .A2(new_n245), .A3(new_n238), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(G101), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(G101), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(KEYINPUT4), .A3(new_n247), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n262));
  AOI211_X1 g076(.A(new_n262), .B(new_n234), .C1(new_n227), .C2(new_n225), .ZN(new_n263));
  INV_X1    g077(.A(new_n234), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n225), .A2(new_n227), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n264), .B1(new_n265), .B2(KEYINPUT70), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n259), .B(new_n261), .C1(new_n263), .C2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n253), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n267), .A2(new_n251), .A3(new_n268), .ZN(new_n269));
  OR4_X1    g083(.A1(new_n222), .A2(new_n255), .A3(new_n256), .A4(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n267), .A2(new_n251), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n253), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n267), .A2(new_n251), .A3(new_n268), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n272), .A2(KEYINPUT86), .A3(KEYINPUT6), .A4(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n268), .B1(new_n267), .B2(new_n251), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n269), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n271), .A2(new_n276), .A3(new_n253), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT86), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n274), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT87), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n219), .B(new_n221), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n282), .B1(new_n281), .B2(new_n283), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n189), .B(new_n270), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(G210), .B1(G237), .B2(G902), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n281), .A2(new_n283), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT87), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n293), .A2(new_n189), .A3(new_n287), .A4(new_n270), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n188), .B1(new_n289), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT15), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n296), .A2(KEYINPUT96), .A3(G478), .ZN(new_n297));
  AOI21_X1  g111(.A(KEYINPUT96), .B1(new_n296), .B2(G478), .ZN(new_n298));
  OR2_X1    g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XOR2_X1   g113(.A(KEYINPUT9), .B(G234), .Z(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(G217), .A3(new_n220), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G122), .ZN(new_n303));
  INV_X1    g117(.A(new_n224), .ZN(new_n304));
  NAND2_X1  g118(.A1(KEYINPUT71), .A2(G116), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G116), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n303), .A2(KEYINPUT93), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT93), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G122), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n307), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(G107), .B1(new_n306), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(G122), .B1(new_n223), .B2(new_n224), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT93), .B(G122), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n313), .B(new_n244), .C1(new_n307), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G134), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT66), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT66), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G134), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n197), .A2(G143), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n321), .B(new_n322), .C1(new_n195), .C2(new_n197), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(KEYINPUT13), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n324), .B1(new_n195), .B2(new_n197), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n212), .A2(KEYINPUT13), .A3(G128), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n325), .A2(new_n326), .A3(KEYINPUT94), .ZN(new_n327));
  OAI21_X1  g141(.A(G134), .B1(new_n325), .B2(KEYINPUT94), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n316), .B(new_n323), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT95), .ZN(new_n330));
  INV_X1    g144(.A(new_n323), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n212), .A2(G128), .B1(KEYINPUT13), .B2(new_n322), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT94), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n317), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n325), .A2(new_n326), .A3(KEYINPUT94), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n331), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT95), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(new_n316), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n330), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n322), .B1(new_n195), .B2(new_n197), .ZN(new_n340));
  INV_X1    g154(.A(new_n321), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n323), .ZN(new_n343));
  OAI221_X1 g157(.A(new_n313), .B1(KEYINPUT14), .B2(new_n244), .C1(new_n307), .C2(new_n314), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT14), .B1(new_n314), .B2(new_n307), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n345), .B(G107), .C1(new_n306), .C2(new_n311), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n302), .B1(new_n339), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n347), .ZN(new_n349));
  AOI211_X1 g163(.A(new_n301), .B(new_n349), .C1(new_n330), .C2(new_n338), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n189), .B(new_n299), .C1(new_n348), .C2(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n329), .A2(KEYINPUT95), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n337), .B1(new_n336), .B2(new_n316), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n347), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n301), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n339), .A2(new_n347), .A3(new_n302), .ZN(new_n356));
  AOI21_X1  g170(.A(G902), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n351), .B1(new_n357), .B2(new_n298), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n220), .A2(G952), .ZN(new_n360));
  NAND2_X1  g174(.A1(G234), .A2(G237), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XOR2_X1   g176(.A(KEYINPUT21), .B(G898), .Z(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(G902), .A3(G953), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT17), .ZN(new_n366));
  NOR2_X1   g180(.A1(G237), .A2(G953), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(G143), .A3(G214), .ZN(new_n368));
  INV_X1    g182(.A(G214), .ZN(new_n369));
  NOR3_X1   g183(.A1(new_n369), .A2(G237), .A3(G953), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n368), .B1(new_n195), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G131), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n209), .A2(new_n211), .B1(new_n367), .B2(G214), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n367), .A2(G143), .A3(G214), .ZN(new_n376));
  OAI211_X1 g190(.A(KEYINPUT90), .B(G131), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT90), .B1(new_n371), .B2(G131), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n366), .B(new_n374), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT16), .ZN(new_n381));
  INV_X1    g195(.A(G140), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(G125), .ZN(new_n383));
  AND2_X1   g197(.A1(G125), .A2(G140), .ZN(new_n384));
  NOR2_X1   g198(.A1(G125), .A2(G140), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n383), .B1(new_n386), .B2(new_n381), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n387), .B(G146), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n371), .A2(G131), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT90), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(KEYINPUT17), .A3(new_n377), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n380), .A2(new_n388), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n371), .A2(KEYINPUT18), .A3(G131), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT18), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n372), .B1(new_n395), .B2(new_n373), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT80), .B1(new_n386), .B2(G146), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n204), .A2(new_n382), .ZN(new_n398));
  NAND2_X1  g212(.A1(G125), .A2(G140), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT80), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(new_n401), .A3(new_n190), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT88), .ZN(new_n404));
  NOR3_X1   g218(.A1(new_n384), .A2(new_n385), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT88), .B1(new_n398), .B2(new_n399), .ZN(new_n406));
  OAI21_X1  g220(.A(G146), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n403), .A2(KEYINPUT89), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(KEYINPUT89), .B1(new_n403), .B2(new_n407), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n394), .B(new_n396), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G113), .B(G122), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(new_n237), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n393), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n412), .B1(new_n393), .B2(new_n410), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n189), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G475), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT20), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n374), .B1(new_n378), .B2(new_n379), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n386), .A2(KEYINPUT19), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n400), .A2(new_n404), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n386), .A2(KEYINPUT88), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n420), .B1(new_n423), .B2(KEYINPUT19), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n190), .ZN(new_n425));
  OR2_X1    g239(.A1(new_n387), .A2(new_n190), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n419), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n412), .B1(new_n410), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT91), .B1(new_n413), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n410), .A2(new_n427), .ZN(new_n430));
  INV_X1    g244(.A(new_n412), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT91), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n393), .A2(new_n410), .A3(new_n412), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n429), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(G475), .A2(G902), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n418), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n437), .B1(KEYINPUT92), .B2(KEYINPUT20), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n437), .A2(KEYINPUT92), .ZN(new_n441));
  AOI211_X1 g255(.A(new_n440), .B(new_n441), .C1(new_n432), .C2(new_n434), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n417), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AND4_X1   g258(.A1(new_n295), .A2(new_n359), .A3(new_n365), .A4(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G221), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(new_n300), .B2(new_n189), .ZN(new_n447));
  INV_X1    g261(.A(G469), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(new_n189), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT85), .ZN(new_n450));
  INV_X1    g264(.A(G137), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT11), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n319), .A2(G134), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n317), .A2(KEYINPUT66), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n451), .A2(KEYINPUT11), .A3(G134), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT11), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G137), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n373), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n455), .A2(new_n459), .A3(new_n373), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT67), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n455), .A2(new_n459), .A3(KEYINPUT67), .A4(new_n373), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(KEYINPUT83), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n203), .A2(KEYINPUT10), .A3(new_n250), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n261), .A2(new_n259), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n467), .B1(new_n218), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT1), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n470), .B1(new_n195), .B2(new_n190), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n196), .B1(new_n471), .B2(new_n197), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n215), .A2(new_n191), .A3(new_n194), .A4(new_n198), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n248), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(KEYINPUT10), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n466), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(G110), .B(G140), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n220), .A2(G227), .ZN(new_n479));
  XOR2_X1   g293(.A(new_n478), .B(new_n479), .Z(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n450), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n456), .A2(new_n458), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n483), .B1(new_n321), .B2(new_n452), .ZN(new_n484));
  AOI21_X1  g298(.A(KEYINPUT67), .B1(new_n484), .B2(new_n373), .ZN(new_n485));
  INV_X1    g299(.A(new_n464), .ZN(new_n486));
  OAI22_X1  g300(.A1(new_n485), .A2(new_n486), .B1(new_n373), .B2(new_n484), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n203), .A2(new_n250), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n487), .B1(new_n488), .B2(new_n474), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT12), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n487), .B(KEYINPUT12), .C1(new_n488), .C2(new_n474), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n466), .A2(new_n476), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(KEYINPUT85), .A3(new_n480), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n482), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  OAI221_X1 g310(.A(new_n467), .B1(new_n218), .B2(new_n468), .C1(new_n474), .C2(KEYINPUT10), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n487), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n481), .ZN(new_n500));
  AOI21_X1  g314(.A(G902), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n449), .B1(new_n501), .B2(new_n448), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT84), .ZN(new_n503));
  AOI22_X1  g317(.A1(new_n492), .A2(new_n491), .B1(new_n466), .B2(new_n476), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(new_n480), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n494), .A2(new_n498), .A3(new_n480), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n503), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n506), .B(KEYINPUT84), .C1(new_n504), .C2(new_n480), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G469), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n447), .B1(new_n502), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n197), .A2(G119), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT76), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n514), .B1(G119), .B2(new_n197), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT24), .B(G110), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OR2_X1    g331(.A1(new_n513), .A2(KEYINPUT79), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n513), .A2(KEYINPUT79), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT23), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n197), .A2(G119), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n518), .B(new_n519), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT78), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n513), .B2(new_n520), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n197), .A2(KEYINPUT78), .A3(KEYINPUT23), .A4(G119), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n517), .B1(new_n526), .B2(G110), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(new_n426), .A3(new_n403), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT81), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n388), .B1(G110), .B2(new_n526), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n515), .A2(new_n516), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n531), .A2(KEYINPUT77), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(KEYINPUT77), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT81), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n527), .A2(new_n535), .A3(new_n426), .A4(new_n403), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n529), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n220), .A2(G221), .A3(G234), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(KEYINPUT22), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(G137), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n537), .A2(new_n541), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT25), .B1(new_n544), .B2(G902), .ZN(new_n545));
  INV_X1    g359(.A(G234), .ZN(new_n546));
  OAI21_X1  g360(.A(G217), .B1(new_n546), .B2(G902), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT25), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n542), .A2(new_n549), .A3(new_n189), .A4(new_n543), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n545), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n547), .A2(new_n189), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(KEYINPUT82), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n542), .A2(new_n553), .A3(new_n543), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT32), .ZN(new_n556));
  XOR2_X1   g370(.A(KEYINPUT73), .B(KEYINPUT27), .Z(new_n557));
  NAND2_X1  g371(.A1(new_n367), .A2(G210), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT26), .B(G101), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n263), .A2(new_n266), .ZN(new_n562));
  INV_X1    g376(.A(new_n218), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n487), .A2(new_n563), .A3(KEYINPUT68), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT68), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n565), .B1(new_n465), .B2(new_n218), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(G134), .A2(G137), .ZN(new_n568));
  OAI211_X1 g382(.A(G131), .B(new_n568), .C1(new_n341), .C2(G137), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n485), .B2(new_n486), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT69), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n463), .A2(new_n464), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(KEYINPUT69), .A3(new_n569), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(new_n203), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n562), .B1(new_n567), .B2(new_n575), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n203), .B(new_n569), .C1(new_n485), .C2(new_n486), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT72), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n487), .A2(new_n563), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n573), .A2(KEYINPUT72), .A3(new_n203), .A4(new_n569), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n579), .A2(new_n580), .A3(new_n562), .A4(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT28), .B1(new_n576), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n562), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n585), .B1(new_n487), .B2(new_n563), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT28), .B1(new_n586), .B2(new_n577), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n561), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT30), .A4(new_n581), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n567), .A2(new_n575), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n585), .B(new_n590), .C1(new_n591), .C2(KEYINPUT30), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n592), .A2(new_n582), .A3(new_n561), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT31), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n592), .A2(KEYINPUT31), .A3(new_n582), .A4(new_n561), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n589), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(G472), .A2(G902), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(KEYINPUT74), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n556), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT30), .B1(new_n567), .B2(new_n575), .ZN(new_n601));
  INV_X1    g415(.A(new_n590), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n583), .B1(new_n603), .B2(new_n585), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT31), .B1(new_n604), .B2(new_n561), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n601), .A2(new_n602), .A3(new_n562), .ZN(new_n606));
  INV_X1    g420(.A(new_n561), .ZN(new_n607));
  NOR4_X1   g421(.A1(new_n606), .A2(new_n594), .A3(new_n583), .A4(new_n607), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n584), .A2(new_n588), .ZN(new_n609));
  OAI22_X1  g423(.A1(new_n605), .A2(new_n608), .B1(new_n561), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n599), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(KEYINPUT32), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT75), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n607), .B1(new_n606), .B2(new_n583), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT29), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n584), .A2(new_n588), .A3(new_n561), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n585), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n582), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n587), .B1(new_n620), .B2(KEYINPUT28), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n607), .A2(new_n615), .ZN(new_n622));
  AOI21_X1  g436(.A(G902), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n613), .B1(new_n624), .B2(G472), .ZN(new_n625));
  INV_X1    g439(.A(G472), .ZN(new_n626));
  AOI211_X1 g440(.A(KEYINPUT75), .B(new_n626), .C1(new_n617), .C2(new_n623), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n600), .B(new_n612), .C1(new_n625), .C2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n445), .A2(new_n512), .A3(new_n555), .A4(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G101), .ZN(G3));
  OAI21_X1  g444(.A(G472), .B1(new_n597), .B2(G902), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n610), .A2(new_n611), .ZN(new_n632));
  AND4_X1   g446(.A1(new_n512), .A2(new_n631), .A3(new_n555), .A4(new_n632), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n348), .A2(new_n350), .A3(KEYINPUT33), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT33), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n355), .B2(new_n356), .ZN(new_n636));
  OAI211_X1 g450(.A(G478), .B(new_n189), .C1(new_n634), .C2(new_n636), .ZN(new_n637));
  OR2_X1    g451(.A1(new_n357), .A2(G478), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n444), .A2(new_n640), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n295), .A2(new_n365), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n633), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT34), .B(G104), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  INV_X1    g459(.A(new_n437), .ZN(new_n646));
  AOI211_X1 g460(.A(KEYINPUT20), .B(new_n646), .C1(new_n429), .C2(new_n435), .ZN(new_n647));
  OAI21_X1  g461(.A(KEYINPUT97), .B1(new_n438), .B2(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n413), .A2(new_n428), .A3(KEYINPUT91), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n433), .B1(new_n432), .B2(new_n434), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n437), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(KEYINPUT20), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT97), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n436), .A2(new_n418), .A3(new_n437), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n648), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n656), .A2(new_n358), .A3(new_n365), .A4(new_n417), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(KEYINPUT98), .ZN(new_n658));
  AOI22_X1  g472(.A1(new_n648), .A2(new_n655), .B1(G475), .B2(new_n416), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT98), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n659), .A2(new_n660), .A3(new_n358), .A4(new_n365), .ZN(new_n661));
  AND3_X1   g475(.A1(new_n658), .A2(new_n295), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n633), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT35), .B(G107), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G9));
  NOR2_X1   g479(.A1(new_n541), .A2(KEYINPUT36), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n537), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n553), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n551), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n512), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n445), .A2(new_n632), .A3(new_n631), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT37), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n672), .B(G110), .Z(G12));
  NAND2_X1  g487(.A1(new_n512), .A2(new_n669), .ZN(new_n674));
  AOI21_X1  g488(.A(KEYINPUT32), .B1(new_n610), .B2(new_n611), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n597), .A2(new_n556), .A3(new_n599), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n621), .A2(new_n622), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n189), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n592), .A2(new_n582), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT29), .B1(new_n680), .B2(new_n607), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n679), .B1(new_n681), .B2(new_n616), .ZN(new_n682));
  OAI21_X1  g496(.A(KEYINPUT75), .B1(new_n682), .B2(new_n626), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n624), .A2(new_n613), .A3(G472), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n674), .B1(new_n677), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n362), .B1(G900), .B2(new_n364), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n659), .A2(new_n687), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n688), .A2(new_n295), .A3(new_n358), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  XOR2_X1   g505(.A(new_n687), .B(KEYINPUT39), .Z(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n512), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT99), .B(KEYINPUT40), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n289), .A2(new_n294), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT38), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n444), .A2(new_n188), .A3(new_n359), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n604), .A2(new_n607), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n189), .B1(new_n620), .B2(new_n561), .ZN(new_n701));
  OAI21_X1  g515(.A(G472), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n612), .A2(new_n600), .A3(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n669), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n696), .A2(new_n698), .A3(new_n699), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n195), .ZN(G45));
  NAND3_X1  g521(.A1(new_n443), .A2(new_n639), .A3(new_n687), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT100), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n443), .A2(new_n639), .A3(KEYINPUT100), .A4(new_n687), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n295), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT101), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n295), .A2(new_n710), .A3(KEYINPUT101), .A4(new_n711), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n714), .A2(new_n628), .A3(new_n670), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT102), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT102), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n686), .A2(new_n718), .A3(new_n715), .A4(new_n714), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G146), .ZN(G48));
  NOR2_X1   g535(.A1(new_n448), .A2(KEYINPUT103), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n501), .B(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n447), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n642), .A2(new_n628), .A3(new_n555), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT41), .B(G113), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  INV_X1    g542(.A(new_n555), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n677), .B2(new_n685), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT104), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n662), .A2(new_n730), .A3(new_n731), .A4(new_n725), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n628), .A2(new_n555), .A3(new_n725), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n658), .A2(new_n295), .A3(new_n661), .ZN(new_n734));
  OAI21_X1  g548(.A(KEYINPUT104), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G116), .ZN(G18));
  AND3_X1   g551(.A1(new_n723), .A2(new_n724), .A3(new_n669), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n445), .A2(new_n628), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G119), .ZN(G21));
  OAI22_X1  g554(.A1(new_n605), .A2(new_n608), .B1(new_n621), .B2(new_n561), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n611), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n631), .A2(new_n555), .A3(new_n742), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n699), .A2(new_n697), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n743), .A2(new_n744), .A3(new_n365), .A4(new_n725), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G122), .ZN(G24));
  NAND3_X1  g560(.A1(new_n631), .A2(new_n742), .A3(new_n669), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT105), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n631), .A2(new_n742), .A3(KEYINPUT105), .A4(new_n669), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n712), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n725), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G125), .ZN(G27));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n754), .B1(new_n697), .B2(new_n188), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n289), .A2(new_n294), .A3(KEYINPUT108), .A4(new_n187), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n628), .A2(new_n555), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT106), .B1(new_n504), .B2(new_n480), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n493), .A2(new_n494), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT106), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n760), .A3(new_n481), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n758), .A2(new_n761), .A3(G469), .A4(new_n506), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT107), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n447), .B1(new_n763), .B2(new_n502), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n710), .A3(new_n711), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT109), .B1(new_n757), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n755), .A2(new_n756), .ZN(new_n768));
  INV_X1    g582(.A(new_n765), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n730), .A2(new_n767), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  XOR2_X1   g584(.A(KEYINPUT110), .B(KEYINPUT42), .Z(new_n771));
  NAND3_X1  g585(.A1(new_n766), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n600), .A2(KEYINPUT111), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n774), .B(new_n556), .C1(new_n597), .C2(new_n599), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n685), .A2(new_n612), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n776), .A2(new_n555), .ZN(new_n777));
  AND4_X1   g591(.A1(new_n710), .A2(new_n755), .A3(new_n711), .A4(new_n756), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n777), .A2(KEYINPUT42), .A3(new_n764), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n772), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G131), .ZN(G33));
  INV_X1    g595(.A(new_n757), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n782), .A2(new_n358), .A3(new_n688), .A4(new_n764), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  OR2_X1    g598(.A1(new_n510), .A2(KEYINPUT45), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n758), .A2(new_n761), .A3(KEYINPUT45), .A4(new_n506), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(G469), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n449), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT46), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n501), .A2(new_n448), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n787), .A2(KEYINPUT46), .A3(new_n788), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n724), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n692), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n640), .A2(new_n443), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n797), .A2(KEYINPUT43), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(KEYINPUT43), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n631), .A2(new_n632), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(new_n801), .A3(new_n669), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT44), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n796), .A2(new_n768), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G137), .ZN(G39));
  INV_X1    g621(.A(KEYINPUT47), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n795), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n794), .A2(KEYINPUT47), .A3(new_n724), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n628), .A2(new_n555), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n778), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G140), .ZN(G42));
  INV_X1    g628(.A(new_n698), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n723), .B(KEYINPUT49), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n815), .A2(new_n555), .A3(new_n797), .A4(new_n816), .ZN(new_n817));
  OR4_X1    g631(.A1(new_n188), .A2(new_n817), .A3(new_n447), .A4(new_n703), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n723), .A2(new_n447), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n809), .A2(new_n810), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n362), .B1(new_n798), .B2(new_n799), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n821), .A2(new_n743), .A3(new_n768), .A4(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(new_n725), .A3(new_n743), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n815), .A2(new_n188), .ZN(new_n825));
  OR4_X1    g639(.A1(KEYINPUT118), .A2(new_n824), .A3(new_n825), .A4(KEYINPUT50), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n822), .A2(new_n768), .A3(new_n725), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n749), .A2(new_n750), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n768), .A2(new_n555), .A3(new_n725), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n703), .A2(new_n362), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n443), .A2(new_n639), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n829), .A2(new_n830), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  XOR2_X1   g649(.A(KEYINPUT118), .B(KEYINPUT50), .Z(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(new_n824), .B2(new_n825), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n823), .A2(new_n826), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n829), .A2(new_n830), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n819), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n360), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n838), .A2(new_n819), .A3(new_n839), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n751), .A2(new_n725), .B1(new_n689), .B2(new_n686), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n687), .A2(KEYINPUT114), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n687), .A2(KEYINPUT114), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n764), .A2(new_n704), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n850), .A2(KEYINPUT115), .A3(new_n703), .A4(new_n744), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n744), .A2(new_n703), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n852), .B1(new_n853), .B2(new_n849), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n720), .A2(new_n846), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n720), .A2(KEYINPUT52), .A3(new_n846), .A4(new_n855), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n726), .A2(new_n745), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n736), .A2(new_n739), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT112), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n359), .A2(new_n863), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n351), .B(new_n863), .C1(new_n357), .C2(new_n298), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n864), .A2(new_n443), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n295), .A2(new_n365), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT113), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT113), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n295), .A2(new_n870), .A3(new_n365), .A4(new_n867), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n869), .A2(new_n633), .A3(new_n871), .ZN(new_n872));
  AND4_X1   g686(.A1(new_n629), .A2(new_n872), .A3(new_n671), .A4(new_n643), .ZN(new_n873));
  OR2_X1    g687(.A1(new_n864), .A2(new_n866), .ZN(new_n874));
  AND4_X1   g688(.A1(new_n628), .A2(new_n670), .A3(new_n688), .A4(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n765), .B1(new_n749), .B2(new_n750), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n768), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n862), .A2(new_n878), .A3(new_n780), .A4(new_n783), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n845), .B1(new_n860), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n780), .A2(new_n783), .ZN(new_n882));
  INV_X1    g696(.A(new_n739), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n732), .B2(new_n735), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n884), .A2(new_n873), .A3(new_n877), .A4(new_n861), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  XOR2_X1   g700(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n887));
  NAND2_X1  g701(.A1(new_n856), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n859), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n886), .A2(new_n889), .A3(KEYINPUT53), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n880), .A2(new_n881), .A3(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n822), .A2(new_n295), .A3(new_n725), .A4(new_n743), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n860), .A2(new_n879), .A3(new_n845), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT53), .B1(new_n886), .B2(new_n889), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT54), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n843), .A2(new_n891), .A3(new_n892), .A4(new_n895), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n833), .A2(new_n641), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n827), .A2(new_n777), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT48), .Z(new_n899));
  NOR3_X1   g713(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(G952), .A2(G953), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n818), .B1(new_n900), .B2(new_n901), .ZN(G75));
  AOI21_X1  g716(.A(new_n189), .B1(new_n880), .B2(new_n890), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(G210), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n281), .B(new_n283), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT55), .Z(new_n907));
  AND3_X1   g721(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n907), .B1(new_n904), .B2(new_n905), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n220), .A2(G952), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(G51));
  NAND2_X1  g725(.A1(new_n496), .A2(new_n500), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n880), .A2(new_n890), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT54), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n891), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n788), .A2(KEYINPUT57), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n788), .A2(KEYINPUT57), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n912), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n787), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n903), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT120), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n910), .B1(new_n919), .B2(new_n923), .ZN(G54));
  NAND2_X1  g738(.A1(KEYINPUT58), .A2(G475), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n886), .A2(new_n889), .A3(KEYINPUT53), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n858), .A2(new_n859), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n844), .B1(new_n886), .B2(new_n928), .ZN(new_n929));
  OAI211_X1 g743(.A(G902), .B(new_n926), .C1(new_n927), .C2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n436), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT121), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT121), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n903), .A2(new_n933), .A3(new_n436), .A4(new_n926), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n910), .B1(new_n930), .B2(new_n931), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n935), .A2(KEYINPUT122), .A3(new_n936), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(G60));
  NOR2_X1   g755(.A1(new_n634), .A2(new_n636), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(G478), .A2(G902), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT59), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n915), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n895), .A2(new_n891), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n943), .B1(new_n947), .B2(new_n945), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n946), .A2(new_n948), .A3(new_n910), .ZN(G63));
  NAND2_X1  g763(.A1(G217), .A2(G902), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT60), .Z(new_n951));
  NAND2_X1  g765(.A1(new_n913), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n544), .ZN(new_n953));
  INV_X1    g767(.A(new_n910), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n913), .A2(new_n667), .A3(new_n951), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT61), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(G66));
  NAND2_X1  g772(.A1(new_n862), .A2(new_n873), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n220), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n363), .A2(G224), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n960), .B(KEYINPUT123), .C1(new_n220), .C2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(KEYINPUT123), .B2(new_n960), .ZN(new_n963));
  INV_X1    g777(.A(G898), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n281), .B1(new_n964), .B2(G953), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT124), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n963), .B(new_n966), .ZN(G69));
  XNOR2_X1  g781(.A(new_n603), .B(new_n424), .ZN(new_n968));
  NAND2_X1  g782(.A1(G900), .A2(G953), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n813), .A2(new_n806), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n720), .A2(new_n846), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n796), .A2(new_n744), .A3(new_n777), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n970), .A2(new_n780), .A3(new_n783), .A4(new_n973), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n968), .B(new_n969), .C1(new_n974), .C2(G953), .ZN(new_n975));
  INV_X1    g789(.A(new_n694), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n782), .B(new_n976), .C1(new_n641), .C2(new_n867), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n971), .A2(KEYINPUT62), .A3(new_n706), .ZN(new_n978));
  AOI21_X1  g792(.A(KEYINPUT62), .B1(new_n971), .B2(new_n706), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n970), .B(new_n977), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT125), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n981), .ZN(new_n983));
  AOI21_X1  g797(.A(G953), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n975), .B1(new_n984), .B2(new_n968), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n220), .B1(G227), .B2(G900), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n986), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n988), .B(new_n975), .C1(new_n984), .C2(new_n968), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n987), .A2(new_n989), .ZN(G72));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT63), .Z(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT126), .Z(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(new_n974), .B2(new_n959), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n680), .B1(new_n994), .B2(KEYINPUT127), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n995), .B(new_n607), .C1(KEYINPUT127), .C2(new_n994), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n614), .A2(new_n593), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n992), .B(new_n997), .C1(new_n893), .C2(new_n894), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n996), .A2(new_n954), .A3(new_n998), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n982), .A2(new_n873), .A3(new_n862), .A4(new_n983), .ZN(new_n1000));
  AOI211_X1 g814(.A(new_n607), .B(new_n604), .C1(new_n1000), .C2(new_n993), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n999), .A2(new_n1001), .ZN(G57));
endmodule


