//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n802, new_n804, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983, new_n984, new_n985;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202));
  INV_X1    g001(.A(G227gat), .ZN(new_n203));
  INV_X1    g002(.A(G233gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206));
  INV_X1    g005(.A(G169gat), .ZN(new_n207));
  INV_X1    g006(.A(G176gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n210));
  AOI22_X1  g009(.A1(new_n209), .A2(new_n210), .B1(G169gat), .B2(G176gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT24), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n215));
  INV_X1    g014(.A(G183gat), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n214), .A2(new_n215), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n211), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT25), .B1(new_n220), .B2(KEYINPUT64), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT25), .ZN(new_n223));
  AOI211_X1 g022(.A(new_n222), .B(new_n223), .C1(new_n211), .C2(new_n219), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT65), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n210), .ZN(new_n226));
  NOR3_X1   g025(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n227));
  OAI22_X1  g026(.A1(new_n226), .A2(new_n227), .B1(new_n207), .B2(new_n208), .ZN(new_n228));
  AND3_X1   g027(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231));
  NOR3_X1   g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT64), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n223), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n220), .A2(KEYINPUT64), .A3(KEYINPUT25), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n225), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n239), .B1(new_n207), .B2(new_n208), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT26), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(new_n207), .A3(new_n208), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n212), .B1(new_n240), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(new_n216), .B2(KEYINPUT27), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT27), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n247), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n216), .A2(KEYINPUT27), .ZN(new_n249));
  NOR2_X1   g048(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n246), .A2(new_n248), .A3(new_n249), .A4(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n247), .A2(G183gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n216), .A2(KEYINPUT27), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n247), .A2(G183gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n249), .A2(new_n256), .A3(KEYINPUT67), .ZN(new_n257));
  AOI21_X1  g056(.A(G190gat), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT28), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n251), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n249), .A2(new_n256), .A3(KEYINPUT67), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT67), .B1(new_n249), .B2(new_n256), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n217), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT28), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(KEYINPUT68), .A3(new_n251), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n244), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(G113gat), .B(G120gat), .Z(new_n269));
  XNOR2_X1  g068(.A(G127gat), .B(G134gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT1), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G113gat), .B(G120gat), .ZN(new_n273));
  INV_X1    g072(.A(G127gat), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n274), .A2(G134gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(G134gat), .ZN(new_n276));
  OAI22_X1  g075(.A1(new_n273), .A2(KEYINPUT1), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n272), .A2(new_n277), .A3(KEYINPUT69), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT69), .B1(new_n272), .B2(new_n277), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NOR3_X1   g079(.A1(new_n238), .A2(new_n268), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n280), .ZN(new_n282));
  INV_X1    g081(.A(new_n244), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT68), .B1(new_n266), .B2(new_n251), .ZN(new_n284));
  INV_X1    g083(.A(new_n251), .ZN(new_n285));
  AOI211_X1 g084(.A(new_n261), .B(new_n285), .C1(new_n265), .C2(KEYINPUT28), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n283), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n225), .A2(new_n237), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n282), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n205), .B1(new_n281), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT32), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT33), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G15gat), .B(G43gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(G71gat), .B(G99gat), .ZN(new_n295));
  XOR2_X1   g094(.A(new_n294), .B(new_n295), .Z(new_n296));
  NAND3_X1  g095(.A1(new_n291), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT32), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n280), .B1(new_n238), .B2(new_n268), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n287), .A2(new_n282), .A3(new_n288), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n298), .B1(new_n301), .B2(new_n205), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n296), .A2(KEYINPUT33), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT70), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n205), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n305), .B1(new_n299), .B2(new_n300), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT70), .ZN(new_n307));
  INV_X1    g106(.A(new_n303), .ZN(new_n308));
  NOR4_X1   g107(.A1(new_n306), .A2(new_n307), .A3(new_n298), .A4(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n297), .B1(new_n304), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n281), .A2(new_n289), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT71), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT34), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n311), .A2(new_n312), .A3(new_n313), .A4(new_n305), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n299), .A2(new_n305), .A3(new_n300), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT71), .B1(new_n315), .B2(KEYINPUT34), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(KEYINPUT34), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n314), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n310), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n290), .A2(KEYINPUT32), .A3(new_n303), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(new_n307), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n302), .A2(KEYINPUT70), .A3(new_n303), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n314), .A2(new_n316), .A3(new_n317), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(new_n324), .A3(new_n297), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n202), .B1(new_n319), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT72), .B1(new_n310), .B2(new_n318), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(G106gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(G50gat), .B(G78gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G141gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(G148gat), .ZN(new_n335));
  INV_X1    g134(.A(G148gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G141gat), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT2), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G155gat), .B(G162gat), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT76), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AND2_X1   g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n344));
  XNOR2_X1  g143(.A(G141gat), .B(G148gat), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n343), .B(new_n344), .C1(new_n345), .C2(KEYINPUT2), .ZN(new_n346));
  AND2_X1   g145(.A1(KEYINPUT77), .A2(G148gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(KEYINPUT77), .A2(G148gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n335), .B1(new_n349), .B2(new_n334), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT2), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n342), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G155gat), .ZN(new_n353));
  INV_X1    g152(.A(G162gat), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n340), .A2(new_n346), .B1(new_n350), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT29), .ZN(new_n357));
  XNOR2_X1  g156(.A(G211gat), .B(G218gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(G197gat), .B(G204gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT22), .ZN(new_n360));
  INV_X1    g159(.A(G211gat), .ZN(new_n361));
  INV_X1    g160(.A(G218gat), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n358), .A2(new_n359), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n358), .B1(new_n363), .B2(new_n359), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n357), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n366), .A2(KEYINPUT80), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT3), .B1(new_n366), .B2(KEYINPUT80), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n356), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n364), .A2(new_n365), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n350), .A2(new_n355), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n335), .A2(new_n337), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(new_n351), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n344), .B1(new_n375), .B2(new_n343), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n338), .A2(KEYINPUT76), .A3(new_n339), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n372), .B(new_n373), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n371), .B1(new_n378), .B2(new_n357), .ZN(new_n379));
  INV_X1    g178(.A(G228gat), .ZN(new_n380));
  OAI22_X1  g179(.A1(new_n369), .A2(new_n379), .B1(new_n380), .B2(new_n204), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n373), .B1(new_n376), .B2(new_n377), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT3), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n380), .A2(new_n204), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n379), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT81), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n382), .A2(new_n371), .A3(new_n357), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n385), .A2(new_n386), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(new_n383), .A3(new_n384), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT81), .B1(new_n390), .B2(new_n379), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n381), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(G22gat), .ZN(new_n393));
  INV_X1    g192(.A(G22gat), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n381), .A2(new_n389), .A3(new_n391), .A4(new_n394), .ZN(new_n395));
  AOI211_X1 g194(.A(KEYINPUT82), .B(new_n333), .C1(new_n393), .C2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n393), .A2(new_n395), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n332), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n393), .A2(KEYINPUT82), .A3(new_n395), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n396), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G8gat), .B(G36gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(G64gat), .B(G92gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT74), .ZN(new_n406));
  AND2_X1   g205(.A1(G226gat), .A2(G233gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(KEYINPUT29), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n408), .B1(new_n238), .B2(new_n268), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n221), .A2(new_n224), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n287), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n409), .A2(new_n370), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n410), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n408), .B1(new_n268), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n287), .A2(new_n407), .A3(new_n288), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n370), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n412), .B1(new_n416), .B2(KEYINPUT73), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT73), .ZN(new_n418));
  AOI211_X1 g217(.A(new_n418), .B(new_n370), .C1(new_n414), .C2(new_n415), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n406), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n287), .A2(new_n407), .A3(new_n288), .ZN(new_n421));
  INV_X1    g220(.A(new_n408), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n422), .B1(new_n287), .B2(new_n410), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n371), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n418), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n416), .A2(KEYINPUT73), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n425), .A2(KEYINPUT74), .A3(new_n426), .A4(new_n412), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n405), .B1(new_n420), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n417), .A2(new_n419), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT30), .B1(new_n429), .B2(new_n405), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT30), .ZN(new_n431));
  NOR4_X1   g230(.A1(new_n417), .A2(new_n419), .A3(new_n431), .A4(new_n404), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n428), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  XOR2_X1   g232(.A(KEYINPUT88), .B(KEYINPUT35), .Z(new_n434));
  NAND2_X1  g233(.A1(new_n272), .A2(new_n277), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n383), .A2(new_n435), .A3(new_n378), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n437), .B1(new_n280), .B2(new_n382), .ZN(new_n438));
  INV_X1    g237(.A(new_n435), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n356), .A2(KEYINPUT4), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(G225gat), .A2(G233gat), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n442), .A2(KEYINPUT5), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n436), .A2(new_n438), .A3(new_n440), .A4(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT78), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n445), .B1(new_n356), .B2(new_n439), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n382), .A2(new_n435), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n382), .A2(new_n445), .A3(new_n435), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n442), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT5), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n356), .B(KEYINPUT4), .C1(new_n278), .C2(new_n279), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n441), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n378), .A2(new_n435), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n356), .A2(new_n372), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT4), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n356), .A2(new_n439), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n453), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n444), .B1(new_n451), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G1gat), .B(G29gat), .ZN(new_n460));
  INV_X1    g259(.A(G85gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(KEYINPUT0), .B(G57gat), .ZN(new_n463));
  XOR2_X1   g262(.A(new_n462), .B(new_n463), .Z(new_n464));
  NAND3_X1  g263(.A1(new_n459), .A2(KEYINPUT6), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT86), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT84), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n459), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g268(.A(KEYINPUT84), .B(new_n444), .C1(new_n451), .C2(new_n458), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(new_n464), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n464), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n472), .B(new_n444), .C1(new_n451), .C2(new_n458), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT6), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n434), .B1(new_n467), .B2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n328), .A2(new_n401), .A3(new_n433), .A4(new_n478), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n401), .A2(new_n319), .A3(new_n325), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n459), .A2(new_n464), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n465), .B1(new_n481), .B2(new_n475), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n417), .A2(new_n404), .A3(new_n419), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n482), .B1(KEYINPUT30), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n420), .A2(new_n427), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n432), .B1(new_n485), .B2(new_n404), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n484), .B1(new_n486), .B2(KEYINPUT75), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT75), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(new_n428), .B2(new_n432), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n480), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT35), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n479), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n465), .A2(KEYINPUT86), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n481), .A2(new_n466), .A3(KEYINPUT6), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT37), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n425), .A2(new_n496), .A3(new_n426), .A4(new_n412), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n405), .A2(KEYINPUT38), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n414), .A2(new_n415), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n496), .B1(new_n499), .B2(new_n370), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n409), .A2(new_n371), .A3(new_n411), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n429), .A2(new_n405), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT87), .B1(new_n495), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n483), .B1(new_n497), .B2(new_n502), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT87), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n507), .A2(new_n508), .A3(new_n467), .A4(new_n477), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n496), .B1(new_n420), .B2(new_n427), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n497), .A2(new_n404), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT38), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n506), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n436), .A2(new_n438), .A3(new_n440), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n442), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n448), .A2(new_n449), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n441), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(KEYINPUT39), .A3(new_n517), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n518), .B(new_n472), .C1(KEYINPUT39), .C2(new_n515), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT40), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT83), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n519), .A2(new_n520), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n515), .A2(KEYINPUT39), .A3(new_n517), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n472), .B1(new_n515), .B2(KEYINPUT39), .ZN(new_n525));
  OAI211_X1 g324(.A(KEYINPUT83), .B(new_n520), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n522), .A2(new_n523), .A3(new_n471), .A4(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT85), .B1(new_n433), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n485), .A2(new_n404), .ZN(new_n529));
  INV_X1    g328(.A(new_n432), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n504), .A2(new_n431), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT85), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n526), .B1(new_n519), .B2(new_n520), .ZN(new_n534));
  INV_X1    g333(.A(new_n471), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n534), .A2(new_n521), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n532), .A2(new_n533), .A3(new_n536), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n513), .A2(new_n528), .A3(new_n401), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n487), .A2(new_n489), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n397), .A2(new_n398), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(new_n333), .A3(new_n400), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(new_n540), .B2(new_n333), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n310), .A2(new_n318), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n324), .B1(new_n323), .B2(new_n297), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT72), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n327), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT36), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT36), .ZN(new_n550));
  NOR3_X1   g349(.A1(new_n545), .A2(new_n546), .A3(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n492), .B1(new_n544), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G43gat), .B(G50gat), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n554), .A2(KEYINPUT15), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n555), .B(KEYINPUT90), .Z(new_n556));
  INV_X1    g355(.A(KEYINPUT89), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT15), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n558), .B1(new_n557), .B2(new_n554), .ZN(new_n559));
  NOR2_X1   g358(.A1(G29gat), .A2(G36gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT14), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT91), .ZN(new_n562));
  OR4_X1    g361(.A1(KEYINPUT91), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(G29gat), .A2(G36gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT92), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  OR3_X1    g365(.A1(new_n556), .A2(new_n559), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n564), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n559), .B1(new_n568), .B2(new_n561), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(KEYINPUT17), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G15gat), .B(G22gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT16), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n571), .B1(new_n572), .B2(G1gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(G1gat), .B2(new_n571), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n574), .B(G8gat), .Z(new_n575));
  AND2_X1   g374(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n567), .A2(new_n569), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT17), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n575), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n576), .A2(new_n579), .B1(new_n580), .B2(new_n577), .ZN(new_n581));
  NAND2_X1  g380(.A1(G229gat), .A2(G233gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(KEYINPUT18), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n577), .B(new_n580), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n582), .B(KEYINPUT13), .Z(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n583), .A2(KEYINPUT93), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G113gat), .B(G141gat), .ZN(new_n588));
  INV_X1    g387(.A(G197gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT11), .B(G169gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT12), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n587), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT18), .B1(new_n581), .B2(new_n582), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n595), .A2(new_n597), .A3(new_n586), .A4(new_n583), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(new_n586), .A3(new_n583), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n599), .A2(new_n587), .A3(new_n594), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n553), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT95), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(G57gat), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n606), .A2(G64gat), .ZN(new_n607));
  INV_X1    g406(.A(G64gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n608), .A2(G57gat), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n605), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G71gat), .A2(G78gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(G71gat), .A2(G78gat), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT94), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n614), .B1(new_n613), .B2(new_n612), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT96), .B1(new_n606), .B2(G64gat), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n617), .B1(G57gat), .B2(new_n608), .ZN(new_n618));
  NOR3_X1   g417(.A1(new_n606), .A2(KEYINPUT96), .A3(G64gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n611), .ZN(new_n620));
  OAI221_X1 g419(.A(new_n605), .B1(new_n618), .B2(new_n619), .C1(new_n620), .C2(new_n612), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n623), .A2(KEYINPUT21), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n622), .B(KEYINPUT98), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n624), .B1(new_n625), .B2(KEYINPUT21), .ZN(new_n626));
  MUX2_X1   g425(.A(new_n624), .B(new_n626), .S(new_n575), .Z(new_n627));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT97), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n216), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(new_n361), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n627), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G127gat), .B(G155gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(KEYINPUT103), .B(G85gat), .Z(new_n639));
  INV_X1    g438(.A(G92gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(G99gat), .A2(G106gat), .ZN(new_n641));
  AOI22_X1  g440(.A1(new_n639), .A2(new_n640), .B1(KEYINPUT8), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n643));
  AOI21_X1  g442(.A(KEYINPUT101), .B1(new_n643), .B2(KEYINPUT7), .ZN(new_n644));
  AND2_X1   g443(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n645));
  OAI211_X1 g444(.A(G85gat), .B(G92gat), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n643), .B(KEYINPUT7), .C1(new_n461), .C2(new_n640), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n647), .B1(new_n646), .B2(new_n648), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n642), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(G99gat), .B(G106gat), .Z(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n652), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n654), .B(new_n642), .C1(new_n649), .C2(new_n650), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n578), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n577), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(G232gat), .A2(G233gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n659), .B(KEYINPUT99), .Z(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n658), .B1(KEYINPUT41), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n660), .B(KEYINPUT41), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n662), .B1(new_n658), .B2(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(G134gat), .B(G162gat), .Z(new_n665));
  XNOR2_X1  g464(.A(G190gat), .B(G218gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n664), .A2(new_n668), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n638), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(G230gat), .A2(G233gat), .ZN(new_n674));
  AND4_X1   g473(.A1(KEYINPUT10), .A2(new_n625), .A3(new_n655), .A4(new_n653), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n622), .B1(new_n655), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n656), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n653), .B(new_n655), .C1(new_n676), .C2(new_n622), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT10), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n674), .B1(new_n675), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n674), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n678), .A2(new_n682), .A3(new_n679), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(G120gat), .B(G148gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(G176gat), .B(G204gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n684), .A2(new_n687), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n673), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n602), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n482), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT105), .B(G1gat), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1324gat));
  NAND3_X1  g497(.A1(new_n602), .A2(new_n532), .A3(new_n693), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT16), .B(G8gat), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n699), .A2(KEYINPUT106), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n699), .A2(KEYINPUT106), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n702), .B1(new_n705), .B2(G8gat), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n701), .B(KEYINPUT107), .Z(new_n707));
  NAND3_X1  g506(.A1(new_n703), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n708), .A2(KEYINPUT108), .A3(new_n700), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT108), .B1(new_n708), .B2(new_n700), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n706), .B1(new_n709), .B2(new_n710), .ZN(G1325gat));
  AOI21_X1  g510(.A(G15gat), .B1(new_n694), .B2(new_n328), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT109), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(new_n549), .B2(new_n551), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n550), .B1(new_n326), .B2(new_n327), .ZN(new_n715));
  INV_X1    g514(.A(new_n551), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n715), .A2(new_n716), .A3(KEYINPUT109), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n719), .A2(G15gat), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n712), .B1(new_n694), .B2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT110), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1326gat));
  NAND2_X1  g522(.A1(new_n694), .A2(new_n542), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT43), .B(G22gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1327gat));
  NOR3_X1   g525(.A1(new_n638), .A2(new_n672), .A3(new_n692), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n602), .A2(new_n727), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n728), .A2(G29gat), .A3(new_n482), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT111), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(KEYINPUT45), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT111), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n729), .B(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n638), .B(KEYINPUT112), .Z(new_n736));
  NAND3_X1  g535(.A1(new_n736), .A2(new_n601), .A3(new_n691), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n672), .A2(KEYINPUT44), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT113), .ZN(new_n739));
  NOR4_X1   g538(.A1(new_n326), .A2(new_n532), .A3(new_n542), .A4(new_n327), .ZN(new_n740));
  AOI22_X1  g539(.A1(new_n740), .A2(new_n478), .B1(new_n490), .B2(KEYINPUT35), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n538), .A2(new_n543), .ZN(new_n742));
  AOI211_X1 g541(.A(new_n739), .B(new_n741), .C1(new_n718), .C2(new_n742), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n715), .A2(KEYINPUT109), .A3(new_n716), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT109), .B1(new_n715), .B2(new_n716), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n543), .B(new_n538), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT113), .B1(new_n746), .B2(new_n492), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n738), .B1(new_n743), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n553), .A2(new_n671), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT44), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n737), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G29gat), .B1(new_n752), .B2(new_n482), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n731), .A2(new_n735), .A3(new_n753), .ZN(G1328gat));
  OAI21_X1  g553(.A(G36gat), .B1(new_n752), .B2(new_n433), .ZN(new_n755));
  OR3_X1    g554(.A1(new_n728), .A2(G36gat), .A3(new_n433), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n756), .A2(KEYINPUT114), .A3(KEYINPUT46), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT114), .B1(new_n756), .B2(KEYINPUT46), .ZN(new_n758));
  OAI221_X1 g557(.A(new_n755), .B1(KEYINPUT46), .B2(new_n756), .C1(new_n757), .C2(new_n758), .ZN(G1329gat));
  INV_X1    g558(.A(KEYINPUT47), .ZN(new_n760));
  INV_X1    g559(.A(new_n328), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n728), .A2(G43gat), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n737), .ZN(new_n763));
  INV_X1    g562(.A(new_n738), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n544), .B1(new_n717), .B2(new_n714), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n739), .B1(new_n765), .B2(new_n741), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n746), .A2(KEYINPUT113), .A3(new_n492), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n764), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n750), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n719), .B(new_n763), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n762), .B1(new_n770), .B2(G43gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n760), .B1(new_n771), .B2(KEYINPUT115), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773));
  INV_X1    g572(.A(G43gat), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n751), .B2(new_n719), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n773), .B(KEYINPUT47), .C1(new_n775), .C2(new_n762), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n772), .A2(new_n776), .ZN(G1330gat));
  INV_X1    g576(.A(G50gat), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n778), .B1(new_n751), .B2(new_n542), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT48), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n728), .A2(G50gat), .A3(new_n401), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n780), .B1(new_n779), .B2(new_n781), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(G1331gat));
  NAND2_X1  g583(.A1(new_n766), .A2(new_n767), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n673), .A2(new_n601), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n692), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT116), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n482), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(new_n606), .ZN(G1332gat));
  NOR2_X1   g590(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n792));
  INV_X1    g591(.A(new_n789), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(new_n793), .B2(new_n532), .ZN(new_n794));
  XOR2_X1   g593(.A(KEYINPUT49), .B(G64gat), .Z(new_n795));
  NOR3_X1   g594(.A1(new_n789), .A2(new_n433), .A3(new_n795), .ZN(new_n796));
  OR3_X1    g595(.A1(new_n794), .A2(KEYINPUT117), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT117), .B1(new_n794), .B2(new_n796), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(G1333gat));
  NOR2_X1   g598(.A1(new_n789), .A2(new_n761), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n719), .A2(G71gat), .ZN(new_n801));
  OAI22_X1  g600(.A1(new_n800), .A2(G71gat), .B1(new_n789), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g602(.A1(new_n793), .A2(new_n542), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(G78gat), .ZN(G1335gat));
  INV_X1    g604(.A(new_n601), .ZN(new_n806));
  INV_X1    g605(.A(new_n638), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(KEYINPUT118), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n692), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n748), .B2(new_n750), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT119), .B1(new_n812), .B2(new_n482), .ZN(new_n813));
  INV_X1    g612(.A(new_n639), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n812), .A2(KEYINPUT119), .A3(new_n482), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n671), .B(new_n809), .C1(new_n765), .C2(new_n741), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n817), .A2(KEYINPUT51), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(KEYINPUT51), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n818), .A2(new_n692), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n695), .A2(new_n639), .ZN(new_n821));
  OAI22_X1  g620(.A1(new_n815), .A2(new_n816), .B1(new_n820), .B2(new_n821), .ZN(G1336gat));
  NOR3_X1   g621(.A1(new_n820), .A2(G92gat), .A3(new_n433), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n640), .B1(new_n811), .B2(new_n532), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT52), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n824), .ZN(new_n826));
  INV_X1    g625(.A(new_n820), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n433), .A2(G92gat), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n826), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n825), .A2(new_n831), .ZN(G1337gat));
  AOI21_X1  g631(.A(G99gat), .B1(new_n827), .B2(new_n328), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n811), .A2(G99gat), .A3(new_n719), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(G1338gat));
  NOR3_X1   g634(.A1(new_n820), .A2(G106gat), .A3(new_n401), .ZN(new_n836));
  INV_X1    g635(.A(G106gat), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(new_n811), .B2(new_n542), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT53), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n838), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n401), .A2(G106gat), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n827), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n839), .A2(new_n844), .ZN(G1339gat));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n687), .B1(new_n681), .B2(KEYINPUT54), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n681), .A2(KEYINPUT54), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n675), .A2(new_n680), .A3(new_n674), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OR3_X1    g650(.A1(new_n675), .A2(new_n674), .A3(new_n680), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n852), .A2(KEYINPUT120), .A3(KEYINPUT54), .A4(new_n681), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n847), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n854), .A2(KEYINPUT55), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n688), .B1(new_n854), .B2(KEYINPUT55), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n597), .A2(new_n586), .A3(new_n583), .A4(new_n593), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n581), .A2(new_n582), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n584), .A2(new_n585), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n592), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n855), .A2(new_n856), .A3(new_n671), .A4(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n601), .A2(new_n855), .A3(new_n856), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n692), .A2(new_n861), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n846), .B(new_n862), .C1(new_n865), .C2(new_n671), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n671), .B1(new_n863), .B2(new_n864), .ZN(new_n867));
  INV_X1    g666(.A(new_n862), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT121), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n866), .A2(new_n869), .A3(new_n736), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n786), .A2(new_n691), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n482), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n872), .A2(new_n433), .A3(new_n480), .ZN(new_n873));
  INV_X1    g672(.A(G113gat), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(new_n874), .A3(new_n601), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n872), .A2(new_n740), .ZN(new_n876));
  OAI21_X1  g675(.A(G113gat), .B1(new_n876), .B2(new_n806), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(G1340gat));
  INV_X1    g677(.A(G120gat), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n873), .A2(new_n879), .A3(new_n692), .ZN(new_n880));
  OAI21_X1  g679(.A(G120gat), .B1(new_n876), .B2(new_n691), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(G1341gat));
  NOR3_X1   g681(.A1(new_n876), .A2(new_n274), .A3(new_n736), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n873), .A2(new_n638), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n883), .B1(new_n884), .B2(new_n274), .ZN(G1342gat));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n672), .A2(G134gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n873), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n873), .A2(new_n887), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(KEYINPUT56), .ZN(new_n893));
  OAI21_X1  g692(.A(G134gat), .B1(new_n876), .B2(new_n672), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n890), .A2(new_n891), .A3(new_n893), .A4(new_n894), .ZN(G1343gat));
  AOI21_X1  g694(.A(new_n401), .B1(new_n870), .B2(new_n871), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n807), .B1(new_n867), .B2(new_n868), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n401), .B1(new_n899), .B2(new_n871), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(new_n897), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n719), .A2(new_n482), .A3(new_n532), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n898), .A2(new_n904), .A3(new_n601), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(G141gat), .ZN(new_n906));
  XNOR2_X1  g705(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n896), .A2(new_n902), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n334), .A3(new_n601), .ZN(new_n910));
  AND3_X1   g709(.A1(new_n906), .A2(new_n907), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n907), .B1(new_n906), .B2(new_n910), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n911), .A2(new_n912), .ZN(G1344gat));
  OR3_X1    g712(.A1(new_n908), .A2(new_n349), .A3(new_n691), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT59), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n899), .A2(new_n871), .ZN(new_n916));
  OAI211_X1 g715(.A(KEYINPUT124), .B(new_n897), .C1(new_n916), .C2(new_n401), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n918), .B1(new_n900), .B2(KEYINPUT57), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  AOI211_X1 g719(.A(new_n897), .B(new_n401), .C1(new_n870), .C2(new_n871), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n692), .B(new_n902), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n915), .B1(new_n922), .B2(G148gat), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n349), .A2(new_n915), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n898), .A2(new_n904), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n925), .B2(new_n692), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n914), .B1(new_n923), .B2(new_n926), .ZN(G1345gat));
  NAND2_X1  g726(.A1(new_n909), .A2(new_n638), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n928), .A2(KEYINPUT125), .ZN(new_n929));
  AOI21_X1  g728(.A(G155gat), .B1(new_n928), .B2(KEYINPUT125), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n736), .A2(new_n353), .ZN(new_n931));
  AOI22_X1  g730(.A1(new_n929), .A2(new_n930), .B1(new_n925), .B2(new_n931), .ZN(G1346gat));
  AOI21_X1  g731(.A(G162gat), .B1(new_n909), .B2(new_n671), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n672), .A2(new_n354), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n933), .B1(new_n925), .B2(new_n934), .ZN(G1347gat));
  NAND2_X1  g734(.A1(new_n870), .A2(new_n871), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n433), .A2(new_n695), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n936), .A2(new_n480), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n938), .A2(new_n207), .A3(new_n601), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n761), .A2(new_n542), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n936), .A2(new_n940), .A3(new_n937), .ZN(new_n941));
  OAI21_X1  g740(.A(G169gat), .B1(new_n941), .B2(new_n806), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n939), .A2(new_n942), .ZN(G1348gat));
  AOI21_X1  g742(.A(G176gat), .B1(new_n938), .B2(new_n692), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n941), .A2(new_n208), .A3(new_n691), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n944), .A2(new_n945), .ZN(G1349gat));
  AOI21_X1  g745(.A(new_n807), .B1(new_n257), .B2(new_n255), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n938), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(G183gat), .B1(new_n941), .B2(new_n736), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g750(.A1(new_n936), .A2(new_n940), .A3(new_n671), .A4(new_n937), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G190gat), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT126), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n952), .A2(new_n955), .A3(G190gat), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n938), .A2(new_n217), .A3(new_n671), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n954), .A2(KEYINPUT61), .A3(new_n956), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(G1351gat));
  AND2_X1   g761(.A1(new_n718), .A2(new_n937), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n896), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n964), .A2(new_n589), .A3(new_n601), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT127), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n963), .B1(new_n920), .B2(new_n921), .ZN(new_n967));
  OAI21_X1  g766(.A(G197gat), .B1(new_n967), .B2(new_n806), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(G1352gat));
  INV_X1    g768(.A(G204gat), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n964), .A2(new_n970), .A3(new_n692), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n972));
  OAI211_X1 g771(.A(new_n692), .B(new_n963), .C1(new_n920), .C2(new_n921), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(G204gat), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(G1353gat));
  NAND3_X1  g775(.A1(new_n964), .A2(new_n361), .A3(new_n638), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n638), .B(new_n963), .C1(new_n920), .C2(new_n921), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n978), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n979));
  AOI21_X1  g778(.A(KEYINPUT63), .B1(new_n978), .B2(G211gat), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(G1354gat));
  NAND2_X1  g780(.A1(new_n671), .A2(G218gat), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n967), .A2(new_n982), .ZN(new_n983));
  INV_X1    g782(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(G218gat), .B1(new_n964), .B2(new_n671), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n984), .A2(new_n985), .ZN(G1355gat));
endmodule


