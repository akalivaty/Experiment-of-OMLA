//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1217, new_n1218, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G20), .ZN(new_n216));
  INV_X1    g0016(.A(new_n201), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n211), .A2(new_n213), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n219), .B(new_n230), .C1(new_n211), .C2(new_n213), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G58), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n248), .A2(new_n221), .ZN(new_n249));
  OR2_X1    g0049(.A1(new_n249), .A2(new_n201), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n250), .A2(G20), .B1(G159), .B2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT7), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n253), .B1(new_n258), .B2(G20), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G68), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n265), .A2(KEYINPUT79), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(KEYINPUT79), .ZN(new_n267));
  OAI211_X1 g0067(.A(KEYINPUT16), .B(new_n252), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n214), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n265), .A2(new_n252), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT16), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n268), .A2(new_n270), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT8), .B(G58), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(new_n206), .B2(G20), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(KEYINPUT80), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n270), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n281), .B1(new_n276), .B2(KEYINPUT80), .ZN(new_n282));
  INV_X1    g0082(.A(new_n280), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n278), .A2(new_n282), .B1(new_n283), .B2(new_n275), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n285));
  INV_X1    g0085(.A(G41), .ZN(new_n286));
  INV_X1    g0086(.A(G45), .ZN(new_n287));
  AOI21_X1  g0087(.A(G1), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G232), .ZN(new_n290));
  INV_X1    g0090(.A(new_n285), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G274), .A3(new_n288), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT81), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT66), .B(G1698), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n258), .A2(new_n295), .A3(G223), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n258), .A2(G1698), .ZN(new_n297));
  INV_X1    g0097(.A(G226), .ZN(new_n298));
  OAI221_X1 g0098(.A(new_n296), .B1(new_n255), .B2(new_n223), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n285), .ZN(new_n300));
  INV_X1    g0100(.A(G190), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n293), .B1(new_n299), .B2(new_n285), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n294), .A2(new_n302), .B1(G200), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n274), .A2(new_n284), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT17), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n274), .A2(KEYINPUT17), .A3(new_n284), .A4(new_n304), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n307), .A2(KEYINPUT83), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(KEYINPUT83), .B1(new_n307), .B2(new_n308), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n274), .A2(new_n284), .ZN(new_n311));
  INV_X1    g0111(.A(G179), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n300), .A2(new_n312), .ZN(new_n313));
  OAI22_X1  g0113(.A1(new_n294), .A2(new_n313), .B1(G169), .B2(new_n303), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT18), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n314), .B1(new_n274), .B2(new_n284), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n319), .A2(KEYINPUT82), .A3(KEYINPUT18), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  AOI211_X1 g0121(.A(new_n317), .B(new_n314), .C1(new_n274), .C2(new_n284), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(KEYINPUT82), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n309), .A2(new_n310), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n292), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n325), .B1(G226), .B2(new_n289), .ZN(new_n326));
  INV_X1    g0126(.A(G1698), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n262), .A2(new_n327), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n328), .A2(G223), .B1(G77), .B2(new_n262), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(KEYINPUT66), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT66), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G1698), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n330), .B(new_n332), .C1(new_n260), .C2(new_n261), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G222), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n326), .B1(new_n336), .B2(new_n291), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(G179), .ZN(new_n338));
  INV_X1    g0138(.A(new_n275), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n207), .A2(G33), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n339), .A2(new_n341), .B1(G150), .B2(new_n251), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n203), .A2(G20), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n279), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n283), .A2(new_n270), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n206), .A2(G20), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(G50), .A3(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(G50), .B2(new_n280), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G169), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n349), .B1(new_n337), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n338), .B1(new_n352), .B2(KEYINPUT67), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(KEYINPUT67), .B2(new_n352), .ZN(new_n354));
  INV_X1    g0154(.A(G244), .ZN(new_n355));
  NOR3_X1   g0155(.A1(new_n285), .A2(new_n288), .A3(new_n355), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n334), .A2(G232), .B1(G107), .B2(new_n262), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n222), .B2(new_n297), .ZN(new_n358));
  AOI211_X1 g0158(.A(new_n325), .B(new_n356), .C1(new_n358), .C2(new_n285), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n359), .A2(new_n312), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n339), .A2(new_n251), .B1(G20), .B2(G77), .ZN(new_n361));
  XOR2_X1   g0161(.A(KEYINPUT15), .B(G87), .Z(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n341), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n279), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n345), .A2(G77), .A3(new_n346), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(G77), .B2(new_n280), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n359), .B2(G169), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n360), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n367), .B1(new_n359), .B2(G190), .ZN(new_n371));
  INV_X1    g0171(.A(G200), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n371), .B1(new_n372), .B2(new_n359), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n354), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n337), .A2(new_n301), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(G200), .B2(new_n337), .ZN(new_n376));
  XOR2_X1   g0176(.A(new_n349), .B(KEYINPUT9), .Z(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT10), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n377), .B(KEYINPUT68), .ZN(new_n380));
  XOR2_X1   g0180(.A(KEYINPUT69), .B(KEYINPUT10), .Z(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n379), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n374), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT14), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT13), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n333), .A2(new_n298), .ZN(new_n388));
  AND3_X1   g0188(.A1(KEYINPUT70), .A2(G33), .A3(G97), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT70), .B1(G33), .B2(G97), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AND2_X1   g0191(.A1(G232), .A2(G1698), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n260), .B2(new_n261), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT71), .ZN(new_n395));
  NOR3_X1   g0195(.A1(new_n388), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G232), .A2(G1698), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(new_n256), .B2(new_n257), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G97), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT70), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(KEYINPUT70), .A2(G33), .A3(G97), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n258), .A2(new_n295), .A3(G226), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT71), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n285), .B1(new_n396), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT72), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n395), .B1(new_n388), .B2(new_n394), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n404), .A2(KEYINPUT71), .A3(new_n405), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n412), .A2(KEYINPUT72), .A3(new_n285), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n289), .A2(G238), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT73), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n415), .A2(new_n416), .A3(new_n292), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n416), .B1(new_n415), .B2(new_n292), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n387), .B1(new_n414), .B2(new_n420), .ZN(new_n421));
  AOI211_X1 g0221(.A(KEYINPUT13), .B(new_n419), .C1(new_n409), .C2(new_n413), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n386), .B(G169), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT72), .B1(new_n412), .B2(new_n285), .ZN(new_n424));
  AOI211_X1 g0224(.A(new_n408), .B(new_n291), .C1(new_n410), .C2(new_n411), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n420), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT13), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n420), .B(new_n387), .C1(new_n424), .C2(new_n425), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(G179), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n350), .B1(new_n427), .B2(new_n428), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT76), .B1(new_n431), .B2(new_n386), .ZN(new_n432));
  OAI21_X1  g0232(.A(G169), .B1(new_n421), .B2(new_n422), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT76), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(new_n434), .A3(KEYINPUT14), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n430), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n283), .A2(new_n221), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n437), .B(KEYINPUT12), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n345), .A2(G68), .A3(new_n346), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT11), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n251), .A2(G50), .B1(G20), .B2(new_n221), .ZN(new_n441));
  INV_X1    g0241(.A(G77), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n441), .B1(new_n442), .B2(new_n340), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n270), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n438), .B(new_n439), .C1(new_n440), .C2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n445), .B1(new_n440), .B2(new_n444), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n446), .B(KEYINPUT74), .ZN(new_n447));
  XNOR2_X1  g0247(.A(new_n447), .B(KEYINPUT77), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n436), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT75), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n427), .A2(G190), .A3(new_n428), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n447), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n372), .B1(new_n427), .B2(new_n428), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(G200), .B1(new_n421), .B2(new_n422), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n456), .A2(KEYINPUT75), .A3(new_n452), .A4(new_n447), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n450), .A2(new_n458), .ZN(new_n459));
  AOI211_X1 g0259(.A(new_n324), .B(new_n385), .C1(new_n459), .C2(KEYINPUT78), .ZN(new_n460));
  OR2_X1    g0260(.A1(new_n459), .A2(KEYINPUT78), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n258), .A2(new_n207), .A3(G87), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n463), .B(KEYINPUT22), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT24), .ZN(new_n465));
  INV_X1    g0265(.A(G107), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G20), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n467), .B(KEYINPUT23), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G116), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G20), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(KEYINPUT90), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT90), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n469), .A2(new_n472), .A3(G20), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n468), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n464), .A2(new_n465), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n465), .B1(new_n464), .B2(new_n474), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n270), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n345), .B1(G1), .B2(new_n255), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT25), .B1(new_n283), .B2(new_n466), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n283), .A2(KEYINPUT25), .A3(new_n466), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n480), .A2(G107), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n478), .A2(KEYINPUT91), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT91), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n463), .A2(KEYINPUT22), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n463), .A2(KEYINPUT22), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n474), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT24), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n279), .B1(new_n490), .B2(new_n475), .ZN(new_n491));
  INV_X1    g0291(.A(new_n484), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n486), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n258), .A2(G257), .A3(G1698), .ZN(new_n494));
  INV_X1    g0294(.A(G294), .ZN(new_n495));
  OAI221_X1 g0295(.A(new_n494), .B1(new_n255), .B2(new_n495), .C1(new_n224), .C2(new_n333), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n285), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n287), .A2(G1), .ZN(new_n498));
  XNOR2_X1  g0298(.A(KEYINPUT5), .B(G41), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n285), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G264), .ZN(new_n501));
  INV_X1    g0301(.A(G274), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n285), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(new_n498), .A3(new_n499), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n497), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G169), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n312), .B2(new_n506), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n485), .A2(new_n493), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n466), .A2(KEYINPUT6), .A3(G97), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT84), .ZN(new_n511));
  OR2_X1    g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n511), .ZN(new_n513));
  XOR2_X1   g0313(.A(G97), .B(G107), .Z(new_n514));
  OAI211_X1 g0314(.A(new_n512), .B(new_n513), .C1(new_n514), .C2(KEYINPUT6), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n515), .A2(G20), .B1(G77), .B2(new_n251), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n264), .A2(G107), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n279), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(G97), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n283), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n479), .B2(new_n519), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n328), .A2(G250), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G283), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n258), .A2(new_n295), .A3(KEYINPUT4), .A4(G244), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT4), .B1(new_n334), .B2(G244), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n285), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n500), .A2(G257), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n530), .A2(new_n504), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n350), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n523), .B(new_n533), .C1(G179), .C2(new_n532), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(G200), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n535), .B(new_n522), .C1(new_n301), .C2(new_n532), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n497), .A2(new_n505), .A3(G190), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n506), .A2(G200), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n478), .A2(new_n484), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n509), .A2(new_n534), .A3(new_n536), .A4(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n525), .B(new_n207), .C1(G33), .C2(new_n519), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n541), .B(new_n270), .C1(new_n207), .C2(G116), .ZN(new_n542));
  XNOR2_X1  g0342(.A(new_n542), .B(KEYINPUT20), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n280), .A2(G116), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(G116), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(new_n479), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n551), .A2(new_n312), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n258), .A2(new_n295), .A3(G257), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n258), .A2(G264), .A3(G1698), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n262), .A2(G303), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n285), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT88), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n556), .A2(KEYINPUT88), .A3(new_n285), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n500), .A2(G270), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n562), .A2(new_n504), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(G169), .B1(new_n543), .B2(new_n548), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n566), .B1(new_n561), .B2(new_n563), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n552), .A2(new_n565), .B1(new_n567), .B2(KEYINPUT21), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n550), .B1(new_n564), .B2(G200), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n301), .B2(new_n564), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n564), .A2(G169), .A3(new_n550), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT21), .ZN(new_n572));
  AOI21_X1  g0372(.A(KEYINPUT89), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT89), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n567), .A2(new_n574), .A3(KEYINPUT21), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n568), .B(new_n570), .C1(new_n573), .C2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n540), .A2(new_n576), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n285), .A2(new_n224), .A3(new_n498), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(new_n498), .B2(new_n503), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n469), .B1(new_n333), .B2(new_n222), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT85), .B1(new_n297), .B2(new_n355), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT85), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n328), .A2(new_n582), .A3(G244), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n580), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n579), .B1(new_n584), .B2(new_n291), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G169), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n312), .B2(new_n585), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT86), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n586), .B(KEYINPUT86), .C1(new_n312), .C2(new_n585), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n403), .A2(KEYINPUT19), .ZN(new_n591));
  NOR2_X1   g0391(.A1(G97), .A2(G107), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n591), .A2(new_n207), .B1(new_n223), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n258), .A2(new_n207), .A3(G68), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n340), .A2(new_n519), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n594), .B1(KEYINPUT19), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n270), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n362), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n283), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n597), .B(new_n599), .C1(new_n598), .C2(new_n479), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n589), .A2(new_n590), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT87), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n597), .A2(new_n599), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n603), .B1(G87), .B2(new_n480), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n585), .A2(G200), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n604), .B(new_n605), .C1(new_n301), .C2(new_n585), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n601), .A2(new_n602), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n601), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(KEYINPUT87), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n577), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n462), .A2(new_n610), .ZN(G372));
  XOR2_X1   g0411(.A(new_n384), .B(KEYINPUT94), .Z(new_n612));
  NOR2_X1   g0412(.A1(new_n309), .A2(new_n310), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n458), .A2(new_n369), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n613), .B1(new_n450), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n322), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT93), .B1(new_n616), .B2(new_n318), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n319), .A2(KEYINPUT18), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT93), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n618), .A2(new_n322), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n612), .B1(new_n615), .B2(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n622), .A2(new_n354), .ZN(new_n623));
  INV_X1    g0423(.A(new_n534), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n609), .A2(new_n607), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT26), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n587), .A2(new_n600), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n606), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT92), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT92), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n628), .A2(new_n606), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n534), .A2(new_n536), .A3(new_n539), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n508), .B1(new_n491), .B2(new_n492), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n568), .B(new_n635), .C1(new_n573), .C2(new_n575), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n633), .A2(new_n638), .A3(new_n624), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n637), .A2(new_n639), .A3(new_n628), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n627), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n623), .B1(new_n462), .B2(new_n641), .ZN(G369));
  OAI21_X1  g0442(.A(new_n568), .B1(new_n573), .B2(new_n575), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(G213), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g0447(.A(KEYINPUT95), .B(G343), .Z(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n551), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n643), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n576), .B2(new_n651), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(G330), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n485), .A2(new_n493), .A3(new_n649), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n656), .A2(new_n509), .A3(new_n539), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n509), .B2(new_n650), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n635), .A2(new_n649), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n643), .A2(new_n650), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(new_n657), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n659), .A2(new_n660), .A3(new_n662), .ZN(G399));
  INV_X1    g0463(.A(new_n210), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(G41), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n592), .A2(new_n223), .A3(new_n547), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(G1), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT96), .ZN(new_n670));
  OAI22_X1  g0470(.A1(new_n669), .A2(new_n670), .B1(new_n218), .B2(new_n666), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n670), .B2(new_n669), .ZN(new_n672));
  XOR2_X1   g0472(.A(new_n672), .B(KEYINPUT28), .Z(new_n673));
  INV_X1    g0473(.A(KEYINPUT99), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n637), .A2(new_n639), .A3(new_n628), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n649), .B1(new_n675), .B2(new_n626), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n674), .B1(new_n676), .B2(KEYINPUT29), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n650), .B1(new_n627), .B2(new_n640), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT29), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(KEYINPUT99), .A3(new_n679), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n509), .B(new_n568), .C1(new_n573), .C2(new_n575), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n633), .A2(new_n634), .A3(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(new_n628), .ZN(new_n683));
  INV_X1    g0483(.A(new_n633), .ZN(new_n684));
  OAI21_X1  g0484(.A(KEYINPUT26), .B1(new_n684), .B2(new_n534), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n683), .B(new_n685), .C1(KEYINPUT26), .C2(new_n625), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n650), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n677), .B(new_n680), .C1(new_n679), .C2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n562), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n585), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n532), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n506), .A2(new_n312), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n690), .A2(new_n691), .A3(new_n692), .A4(new_n561), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  AND4_X1   g0494(.A1(new_n312), .A2(new_n532), .A3(new_n585), .A4(new_n506), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n693), .A2(new_n694), .B1(new_n695), .B2(new_n564), .ZN(new_n696));
  AND4_X1   g0496(.A1(new_n561), .A2(new_n690), .A3(new_n691), .A4(new_n692), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT97), .B1(new_n697), .B2(KEYINPUT30), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT97), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n693), .A2(new_n699), .A3(new_n694), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n696), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(KEYINPUT31), .A3(new_n649), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT98), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n701), .A2(new_n649), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n577), .A2(new_n607), .A3(new_n609), .A4(new_n650), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n706), .B1(new_n707), .B2(KEYINPUT31), .ZN(new_n708));
  OAI21_X1  g0508(.A(G330), .B1(new_n704), .B2(new_n708), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n688), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n673), .B1(new_n710), .B2(G1), .ZN(G364));
  AOI21_X1  g0511(.A(new_n214), .B1(G20), .B2(new_n350), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n207), .A2(G179), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(G190), .A3(G200), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n223), .ZN(new_n716));
  NOR2_X1   g0516(.A1(G190), .A2(G200), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G159), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(KEYINPUT32), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n207), .A2(new_n312), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G200), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G190), .ZN(new_n724));
  AOI211_X1 g0524(.A(new_n716), .B(new_n721), .C1(G68), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n722), .A2(new_n717), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n258), .B1(new_n726), .B2(new_n442), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n722), .A2(G190), .A3(new_n372), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n727), .B1(G58), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n714), .A2(new_n301), .A3(G200), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n720), .A2(KEYINPUT32), .B1(G107), .B2(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n301), .A2(G179), .A3(G200), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(new_n207), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n723), .A2(new_n301), .ZN(new_n737));
  AOI22_X1  g0537(.A1(G97), .A2(new_n736), .B1(new_n737), .B2(G50), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n725), .A2(new_n730), .A3(new_n733), .A4(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G322), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n728), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(G311), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n262), .B1(new_n726), .B2(new_n742), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n741), .B(new_n743), .C1(G329), .C2(new_n719), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n737), .A2(G326), .ZN(new_n745));
  XNOR2_X1  g0545(.A(KEYINPUT33), .B(G317), .ZN(new_n746));
  INV_X1    g0546(.A(new_n715), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n724), .A2(new_n746), .B1(new_n747), .B2(G303), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n736), .A2(G294), .B1(new_n732), .B2(G283), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n744), .A2(new_n745), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n713), .B1(new_n739), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G13), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n206), .B1(new_n753), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n665), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n210), .A2(new_n258), .ZN(new_n757));
  INV_X1    g0557(.A(G355), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n757), .A2(new_n758), .B1(G116), .B2(new_n210), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n664), .A2(new_n258), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n218), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n761), .B1(new_n287), .B2(new_n762), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n243), .A2(new_n287), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n759), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT100), .Z(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n712), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n756), .B1(new_n765), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n751), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n768), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n772), .B1(new_n653), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n756), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n654), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n653), .A2(G330), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT101), .Z(G396));
  INV_X1    g0579(.A(new_n367), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n373), .B1(new_n780), .B2(new_n650), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n370), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n369), .A2(new_n650), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n678), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n676), .A2(new_n786), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n756), .B1(new_n790), .B2(new_n709), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n709), .B2(new_n790), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n712), .A2(new_n766), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n775), .B1(new_n442), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G132), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n258), .B1(new_n718), .B2(new_n795), .C1(new_n221), .C2(new_n731), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n735), .A2(new_n248), .B1(new_n715), .B2(new_n202), .ZN(new_n797));
  INV_X1    g0597(.A(new_n726), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n729), .A2(G143), .B1(new_n798), .B2(G159), .ZN(new_n799));
  INV_X1    g0599(.A(new_n724), .ZN(new_n800));
  INV_X1    g0600(.A(G150), .ZN(new_n801));
  INV_X1    g0601(.A(G137), .ZN(new_n802));
  INV_X1    g0602(.A(new_n737), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n799), .B1(new_n800), .B2(new_n801), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT103), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT34), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n796), .B(new_n797), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n735), .A2(new_n519), .B1(new_n728), .B2(new_n495), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT102), .ZN(new_n810));
  INV_X1    g0610(.A(G303), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n803), .A2(new_n811), .B1(new_n731), .B2(new_n223), .ZN(new_n812));
  INV_X1    g0612(.A(G283), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n800), .A2(new_n813), .B1(new_n715), .B2(new_n466), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n262), .B1(new_n718), .B2(new_n742), .C1(new_n547), .C2(new_n726), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n807), .A2(new_n808), .B1(new_n810), .B2(new_n816), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n794), .B1(new_n713), .B2(new_n817), .C1(new_n786), .C2(new_n767), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n792), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G384));
  NOR2_X1   g0620(.A1(new_n753), .A2(new_n206), .ZN(new_n821));
  INV_X1    g0621(.A(G330), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n702), .A2(KEYINPUT112), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT112), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n701), .A2(new_n824), .A3(KEYINPUT31), .A4(new_n649), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n786), .B1(new_n708), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT107), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n448), .A2(new_n650), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n455), .A2(new_n457), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n432), .A2(new_n435), .ZN(new_n831));
  INV_X1    g0631(.A(new_n430), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n828), .B(new_n829), .C1(new_n830), .C2(new_n833), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n447), .B(KEYINPUT77), .Z(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n649), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n836), .B(new_n458), .C1(new_n448), .C2(new_n436), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n458), .A2(new_n436), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n828), .B1(new_n839), .B2(new_n829), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT108), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n839), .A2(new_n829), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(KEYINPUT107), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT108), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n843), .A2(new_n844), .A3(new_n837), .A4(new_n834), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n827), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n284), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n268), .A2(new_n270), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n252), .B1(new_n266), .B2(new_n267), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n272), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n847), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n851), .A2(new_n647), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n324), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n305), .B1(new_n851), .B2(new_n647), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n851), .A2(new_n314), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT37), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n305), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n857), .A2(new_n319), .ZN(new_n858));
  INV_X1    g0658(.A(new_n647), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT37), .B1(new_n311), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n853), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n853), .A2(KEYINPUT38), .A3(new_n862), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT40), .B1(new_n846), .B2(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n307), .B(new_n308), .C1(new_n617), .C2(new_n620), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n311), .A2(new_n859), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT111), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n858), .B2(new_n860), .ZN(new_n873));
  AND4_X1   g0673(.A1(new_n872), .A2(new_n860), .A3(new_n305), .A4(new_n316), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT110), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n857), .B2(new_n319), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n316), .A2(KEYINPUT110), .A3(new_n305), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n877), .A2(new_n878), .A3(new_n870), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n869), .A2(new_n871), .B1(new_n875), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n866), .B1(new_n881), .B2(KEYINPUT38), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n882), .A2(KEYINPUT40), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n868), .B1(new_n846), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n708), .ZN(new_n885));
  INV_X1    g0685(.A(new_n826), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n462), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n822), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n884), .B2(new_n887), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT39), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n882), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT109), .B1(new_n449), .B2(new_n650), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n449), .A2(KEYINPUT109), .A3(new_n650), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n891), .B(new_n895), .C1(new_n867), .C2(new_n890), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n621), .A2(new_n647), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n841), .A2(new_n845), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n785), .B1(new_n676), .B2(new_n786), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n867), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n896), .B(new_n897), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n623), .B1(new_n688), .B2(new_n462), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n903), .B(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n821), .B1(new_n889), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n905), .B2(new_n889), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n216), .A2(new_n547), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n515), .B(KEYINPUT104), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT35), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n911), .B2(new_n910), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT106), .ZN(new_n914));
  XNOR2_X1  g0714(.A(KEYINPUT105), .B(KEYINPUT36), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n914), .B(new_n915), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n218), .A2(new_n442), .A3(new_n249), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n221), .A2(G50), .ZN(new_n918));
  OAI211_X1 g0718(.A(G1), .B(new_n752), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n907), .A2(new_n916), .A3(new_n919), .ZN(G367));
  NAND2_X1  g0720(.A1(new_n624), .A2(new_n649), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n534), .B(new_n536), .C1(new_n522), .C2(new_n650), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n662), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n534), .B1(new_n922), .B2(new_n509), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n925), .A2(KEYINPUT42), .B1(new_n650), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(KEYINPUT42), .B2(new_n925), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT43), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n604), .A2(new_n650), .ZN(new_n930));
  MUX2_X1   g0730(.A(new_n684), .B(new_n628), .S(new_n930), .Z(new_n931));
  OAI21_X1  g0731(.A(new_n928), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n929), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n932), .B(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n659), .A2(new_n924), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n934), .B(new_n935), .Z(new_n936));
  INV_X1    g0736(.A(new_n661), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n662), .B1(new_n658), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n655), .B(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n710), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n662), .A2(new_n660), .A3(new_n923), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT45), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n662), .A2(new_n660), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n924), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT44), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n944), .A2(KEYINPUT44), .A3(new_n924), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n943), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n659), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n950), .B(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n710), .B1(new_n940), .B2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n665), .B(KEYINPUT41), .Z(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n936), .B(KEYINPUT113), .C1(new_n956), .C2(new_n755), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT113), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n755), .B1(new_n953), .B2(new_n955), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n934), .B(new_n935), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n957), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n931), .A2(new_n768), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n770), .B1(new_n664), .B2(new_n362), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n760), .A2(new_n239), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n775), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n724), .A2(G294), .B1(new_n732), .B2(G97), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n967), .B1(new_n466), .B2(new_n735), .C1(new_n742), .C2(new_n803), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n729), .A2(G303), .B1(new_n719), .B2(G317), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT46), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n715), .B2(new_n547), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n747), .A2(KEYINPUT46), .A3(G116), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n258), .B1(new_n798), .B2(G283), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n969), .A2(new_n971), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n731), .A2(new_n442), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G58), .B2(new_n747), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n221), .B2(new_n735), .ZN(new_n977));
  AOI22_X1  g0777(.A1(G143), .A2(new_n737), .B1(new_n724), .B2(G159), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n262), .B1(new_n729), .B2(G150), .ZN(new_n979));
  AOI22_X1  g0779(.A1(G50), .A2(new_n798), .B1(new_n719), .B2(G137), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n968), .A2(new_n974), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT47), .Z(new_n983));
  OAI211_X1 g0783(.A(new_n963), .B(new_n966), .C1(new_n713), .C2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n962), .A2(new_n984), .ZN(G387));
  NOR2_X1   g0785(.A1(new_n658), .A2(new_n773), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n236), .A2(new_n287), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT114), .Z(new_n988));
  NOR2_X1   g0788(.A1(new_n275), .A2(G50), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT50), .ZN(new_n990));
  AOI211_X1 g0790(.A(G45), .B(new_n667), .C1(G68), .C2(G77), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n761), .B(new_n988), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n757), .A2(new_n668), .B1(G107), .B2(new_n210), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n769), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n756), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n726), .A2(new_n221), .B1(new_n718), .B2(new_n801), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n262), .B(new_n996), .C1(G50), .C2(new_n729), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n715), .A2(new_n442), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n362), .A2(new_n736), .B1(new_n724), .B2(new_n339), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n737), .A2(G159), .B1(new_n732), .B2(G97), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n258), .B1(new_n719), .B2(G326), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n735), .A2(new_n813), .B1(new_n715), .B2(new_n495), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n729), .A2(G317), .B1(new_n798), .B2(G303), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n800), .B2(new_n742), .C1(new_n740), .C2(new_n803), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT48), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n1007), .B2(new_n1006), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT49), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1003), .B1(new_n547), .B2(new_n731), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1002), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n986), .B(new_n995), .C1(new_n712), .C2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n939), .B2(new_n755), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n940), .A2(new_n665), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n710), .A2(new_n939), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(G393));
  AND2_X1   g0818(.A1(new_n940), .A2(new_n952), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n665), .B1(new_n940), .B2(new_n952), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n952), .A2(new_n754), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n924), .A2(new_n768), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G317), .A2(new_n737), .B1(new_n729), .B2(G311), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT52), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n262), .B1(new_n718), .B2(new_n740), .C1(new_n495), .C2(new_n726), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n466), .A2(new_n731), .B1(new_n715), .B2(new_n813), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n800), .A2(new_n811), .B1(new_n547), .B2(new_n735), .ZN(new_n1028));
  OR4_X1    g0828(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n735), .A2(new_n442), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n800), .A2(new_n202), .B1(new_n731), .B2(new_n223), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1030), .B(new_n1031), .C1(G68), .C2(new_n747), .ZN(new_n1032));
  INV_X1    g0832(.A(G159), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n803), .A2(new_n801), .B1(new_n1033), .B2(new_n728), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT51), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n798), .A2(new_n339), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n262), .B1(new_n719), .B2(G143), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1032), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n713), .B1(new_n1029), .B2(new_n1038), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n761), .A2(new_n246), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n770), .B1(G97), .B2(new_n664), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n775), .B(new_n1039), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1022), .B1(new_n1023), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1021), .A2(new_n1043), .ZN(G390));
  OAI211_X1 g0844(.A(G330), .B(new_n786), .C1(new_n708), .C2(new_n826), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n898), .A2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g0847(.A(G330), .B(new_n786), .C1(new_n704), .C2(new_n708), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n841), .B2(new_n845), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n784), .B1(new_n687), .B2(new_n783), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n1047), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n898), .A2(new_n1046), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT116), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n898), .A2(KEYINPUT116), .A3(new_n1046), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n841), .A2(new_n845), .A3(new_n1048), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1051), .B1(new_n1057), .B2(new_n900), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n822), .B1(new_n885), .B2(new_n886), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n460), .A2(new_n461), .A3(new_n1059), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1060), .B(new_n623), .C1(new_n688), .C2(new_n462), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n891), .B1(new_n867), .B2(new_n890), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n899), .B1(new_n845), .B2(new_n841), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1063), .B1(new_n1064), .B2(new_n895), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n898), .A2(new_n1050), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT115), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n894), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1067), .B1(new_n1068), .B2(new_n892), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n893), .A2(KEYINPUT115), .A3(new_n894), .ZN(new_n1070));
  AND3_X1   g0870(.A1(new_n1069), .A2(new_n1070), .A3(new_n882), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1066), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1049), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1065), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n895), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n901), .A2(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1076), .A2(new_n1063), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1077));
  AOI21_X1  g0877(.A(KEYINPUT116), .B1(new_n898), .B2(new_n1046), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1053), .B(new_n1045), .C1(new_n841), .C2(new_n845), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1074), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n666), .B1(new_n1062), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT117), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1081), .B(new_n1084), .C1(new_n1061), .C2(new_n1058), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  OR3_X1    g0886(.A1(new_n1047), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1056), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1078), .A2(new_n1079), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1087), .B1(new_n1089), .B2(new_n899), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1061), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1084), .B1(new_n1092), .B2(new_n1081), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1083), .B1(new_n1086), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1082), .A2(new_n755), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n767), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1063), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n775), .B1(new_n275), .B2(new_n793), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n803), .A2(new_n813), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1030), .B(new_n1099), .C1(G107), .C2(new_n724), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n258), .B1(new_n798), .B2(G97), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n729), .A2(G116), .B1(new_n719), .B2(G294), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n716), .B1(G68), .B2(new_n732), .ZN(new_n1103));
  AND4_X1   g0903(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1104), .A2(KEYINPUT119), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n735), .A2(new_n1033), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n800), .A2(new_n802), .B1(new_n731), .B2(new_n202), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(G128), .C2(new_n737), .ZN(new_n1108));
  XOR2_X1   g0908(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1109));
  NAND3_X1  g0909(.A1(new_n747), .A2(G150), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1109), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n801), .B2(new_n715), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT54), .B(G143), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n728), .A2(new_n795), .B1(new_n726), .B2(new_n1113), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n262), .B(new_n1114), .C1(G125), .C2(new_n719), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1108), .A2(new_n1110), .A3(new_n1112), .A4(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1105), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(KEYINPUT119), .B2(new_n1104), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1097), .B(new_n1098), .C1(new_n713), .C2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1095), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1094), .A2(new_n1121), .ZN(G378));
  INV_X1    g0922(.A(new_n903), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n827), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n898), .A2(new_n867), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT40), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n822), .B1(new_n846), .B2(new_n883), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n349), .A2(new_n647), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n612), .B2(new_n354), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n612), .A2(new_n354), .A3(new_n1130), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1134), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1127), .A2(new_n1128), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1137), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1123), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1137), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n846), .A2(new_n883), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(G330), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1141), .B1(new_n1143), .B2(new_n868), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1127), .A2(new_n1128), .A3(new_n1137), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1144), .A2(new_n903), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1140), .A2(new_n1146), .A3(KEYINPUT122), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1091), .B1(new_n1081), .B2(new_n1058), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT122), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1144), .A2(new_n903), .A3(new_n1149), .A4(new_n1145), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT57), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1152), .B1(new_n1140), .B2(new_n1146), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n666), .B1(new_n1154), .B2(new_n1148), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1147), .A2(new_n755), .A3(new_n1150), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n803), .A2(new_n547), .B1(new_n221), .B2(new_n735), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1159), .B(KEYINPUT121), .Z(new_n1160));
  OAI211_X1 g0960(.A(new_n286), .B(new_n262), .C1(new_n728), .C2(new_n466), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n598), .A2(new_n726), .B1(new_n813), .B2(new_n718), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n999), .B1(new_n248), .B2(new_n731), .C1(new_n800), .C2(new_n519), .ZN(new_n1163));
  OR4_X1    g0963(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n255), .A2(new_n286), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT120), .ZN(new_n1167));
  AOI21_X1  g0967(.A(G50), .B1(new_n262), .B2(new_n286), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1165), .A2(KEYINPUT58), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n737), .A2(G125), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n800), .B2(new_n795), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n729), .A2(G128), .B1(new_n798), .B2(G137), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n715), .B2(new_n1113), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1171), .B(new_n1173), .C1(G150), .C2(new_n736), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1167), .B1(G124), .B2(new_n719), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT59), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1177), .B1(new_n1033), .B2(new_n731), .C1(new_n1174), .C2(new_n1178), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1169), .B1(KEYINPUT58), .B2(new_n1165), .C1(new_n1176), .C2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n712), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n775), .B1(new_n202), .B2(new_n793), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(new_n1141), .C2(new_n767), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1158), .A2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1157), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(G375));
  NAND2_X1  g0986(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1092), .A2(new_n1187), .A3(new_n955), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n547), .A2(new_n800), .B1(new_n803), .B2(new_n495), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G97), .B2(new_n747), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n728), .A2(new_n813), .B1(new_n726), .B2(new_n466), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n258), .B(new_n1191), .C1(G303), .C2(new_n719), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n975), .B1(new_n362), .B2(new_n736), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1190), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n735), .A2(new_n202), .B1(new_n715), .B2(new_n1033), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G132), .B2(new_n737), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n262), .B1(new_n719), .B2(G128), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n729), .A2(G137), .B1(new_n798), .B2(G150), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1113), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n724), .A2(new_n1199), .B1(new_n732), .B2(G58), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .A4(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n713), .B1(new_n1194), .B2(new_n1201), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n775), .B(new_n1202), .C1(new_n221), .C2(new_n793), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n766), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1203), .B1(new_n898), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n1058), .B2(new_n754), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1188), .A2(new_n1207), .ZN(G381));
  INV_X1    g1008(.A(G390), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n819), .ZN(new_n1210));
  OR2_X1    g1010(.A1(G393), .A2(G396), .ZN(new_n1211));
  NOR4_X1   g1011(.A1(G387), .A2(new_n1210), .A3(G381), .A4(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(KEYINPUT117), .B1(new_n1062), .B2(new_n1082), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n1085), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1120), .B1(new_n1214), .B2(new_n1083), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1212), .A2(new_n1215), .A3(new_n1185), .ZN(G407));
  NAND2_X1  g1016(.A1(new_n648), .A2(G213), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1185), .A2(new_n1215), .A3(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(G407), .A2(G213), .A3(new_n1219), .ZN(G409));
  XOR2_X1   g1020(.A(G393), .B(G396), .Z(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n962), .A2(new_n984), .A3(G390), .ZN(new_n1223));
  AOI21_X1  g1023(.A(G390), .B1(new_n962), .B2(new_n984), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1222), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(G387), .A2(new_n1209), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n962), .A2(new_n984), .A3(G390), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1226), .A2(new_n1221), .A3(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT61), .ZN(new_n1229));
  AND3_X1   g1029(.A1(new_n1225), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT124), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT60), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n665), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(KEYINPUT60), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1236), .A2(new_n1187), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1231), .B1(new_n1235), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n666), .B1(new_n1236), .B2(new_n1187), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(KEYINPUT124), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1238), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(G384), .B1(new_n1242), .B2(new_n1207), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n819), .B(new_n1206), .C1(new_n1238), .C2(new_n1241), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1184), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(G378), .A2(new_n1156), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1140), .A2(new_n1146), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT123), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1140), .A2(new_n1146), .A3(KEYINPUT123), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1250), .A2(new_n755), .A3(new_n1251), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1147), .A2(new_n1148), .A3(new_n955), .A4(new_n1150), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1252), .A2(new_n1183), .A3(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1215), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1218), .B1(new_n1247), .B2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1245), .A2(new_n1256), .A3(KEYINPUT63), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1230), .A2(new_n1257), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1235), .A2(new_n1237), .A3(new_n1231), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT124), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1207), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n819), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1242), .A2(G384), .A3(new_n1207), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1262), .A2(G2897), .A3(new_n1218), .A4(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1218), .A2(G2897), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1264), .B1(new_n1266), .B2(new_n1256), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT125), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1247), .A2(new_n1255), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1270), .A2(new_n1217), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT63), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1264), .B(KEYINPUT125), .C1(new_n1266), .C2(new_n1256), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1258), .A2(new_n1269), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1225), .A2(new_n1228), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1271), .A2(KEYINPUT62), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1245), .A2(new_n1256), .A3(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1264), .B(new_n1229), .C1(new_n1266), .C2(new_n1256), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1276), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1275), .A2(new_n1282), .ZN(G405));
  INV_X1    g1083(.A(KEYINPUT127), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1276), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1276), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(KEYINPUT127), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1215), .B1(new_n1157), .B2(new_n1184), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(KEYINPUT126), .A3(new_n1247), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT126), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1290), .B(new_n1215), .C1(new_n1157), .C2(new_n1184), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1289), .A2(new_n1245), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1245), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1285), .B(new_n1287), .C1(new_n1293), .C2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1294), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1296), .A2(KEYINPUT127), .A3(new_n1286), .A4(new_n1292), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1295), .A2(new_n1297), .ZN(G402));
endmodule


