//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 0 1 1 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n557, new_n558, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1257, new_n1258,
    new_n1259, new_n1260;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT68), .Z(new_n451));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n451), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n451), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n461), .A2(G137), .A3(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n470), .B1(new_n461), .B2(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n468), .B1(new_n471), .B2(new_n462), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(G125), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n469), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n467), .B1(new_n472), .B2(new_n477), .ZN(G160));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n464), .ZN(new_n480));
  NAND2_X1  g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  AOI21_X1  g056(.A(G2105), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n462), .B1(new_n480), .B2(new_n481), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OR2_X1    g064(.A1(new_n462), .A2(G114), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(G126), .B(G2105), .C1(new_n473), .C2(new_n474), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n462), .C1(new_n473), .C2(new_n474), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n482), .A2(new_n498), .A3(G138), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(G164));
  XNOR2_X1  g075(.A(KEYINPUT6), .B(G651), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(G50), .A3(G543), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n503));
  XNOR2_X1  g078(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(G75), .A2(G543), .ZN(new_n505));
  AND3_X1   g080(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n506));
  AOI21_X1  g081(.A(KEYINPUT5), .B1(KEYINPUT71), .B2(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n506), .A2(new_n507), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n510), .A2(G651), .B1(new_n514), .B2(G88), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n504), .A2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT73), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n501), .A2(G543), .ZN(new_n521));
  AOI22_X1  g096(.A1(G51), .A2(new_n521), .B1(new_n514), .B2(G89), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT71), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT5), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(G63), .A3(G651), .ZN(new_n529));
  XOR2_X1   g104(.A(new_n529), .B(KEYINPUT72), .Z(new_n530));
  NOR2_X1   g105(.A1(new_n523), .A2(new_n530), .ZN(G168));
  XOR2_X1   g106(.A(KEYINPUT74), .B(G90), .Z(new_n532));
  NAND2_X1  g107(.A1(new_n514), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n501), .A2(G543), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n528), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G651), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n536), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n508), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G651), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT75), .ZN(new_n546));
  OAI211_X1 g121(.A(G43), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  OAI211_X1 g123(.A(new_n546), .B(new_n547), .C1(new_n513), .C2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n528), .A2(G81), .A3(new_n501), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n546), .B1(new_n551), .B2(new_n547), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n545), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT77), .ZN(new_n558));
  XOR2_X1   g133(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n559));
  XNOR2_X1  g134(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  NAND3_X1  g136(.A1(new_n501), .A2(G53), .A3(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n501), .A2(new_n564), .A3(G53), .A4(G543), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n514), .A2(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT78), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(new_n526), .B2(new_n527), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n566), .A2(new_n567), .A3(new_n572), .ZN(G299));
  INV_X1    g148(.A(G168), .ZN(G286));
  NAND2_X1  g149(.A1(new_n521), .A2(G49), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n514), .A2(G87), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G288));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  OR3_X1    g154(.A1(new_n513), .A2(KEYINPUT79), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT79), .B1(new_n513), .B2(new_n579), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n528), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G48), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n583), .A2(new_n538), .B1(new_n584), .B2(new_n535), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT80), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n508), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(new_n521), .B2(G48), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT80), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n590), .A2(new_n591), .A3(new_n581), .A4(new_n580), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n586), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n595), .A2(new_n538), .ZN(new_n596));
  INV_X1    g171(.A(G47), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n535), .A2(new_n597), .B1(new_n513), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(KEYINPUT81), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT81), .ZN(new_n601));
  OAI221_X1 g176(.A(new_n601), .B1(new_n513), .B2(new_n598), .C1(new_n597), .C2(new_n535), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n596), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n508), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G651), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n521), .A2(G54), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  NAND4_X1  g186(.A1(new_n611), .A2(new_n528), .A3(G92), .A4(new_n501), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n610), .B1(new_n513), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g189(.A1(new_n608), .A2(new_n609), .A3(new_n612), .A4(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G171), .B2(new_n616), .ZN(G284));
  OAI21_X1  g193(.A(new_n617), .B1(G171), .B2(new_n616), .ZN(G321));
  NAND2_X1  g194(.A1(G299), .A2(new_n616), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G168), .B2(new_n616), .ZN(G297));
  XNOR2_X1  g196(.A(G297), .B(KEYINPUT83), .ZN(G280));
  INV_X1    g197(.A(new_n615), .ZN(new_n623));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G860), .ZN(G148));
  NOR2_X1   g200(.A1(new_n615), .A2(G559), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT84), .ZN(new_n627));
  MUX2_X1   g202(.A(new_n553), .B(new_n627), .S(G868), .Z(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XOR2_X1   g204(.A(KEYINPUT85), .B(KEYINPUT12), .Z(new_n630));
  NAND3_X1  g205(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT85), .B(KEYINPUT12), .ZN(new_n633));
  INV_X1    g208(.A(new_n631), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  INV_X1    g212(.A(G2100), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n482), .A2(G135), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n484), .A2(G123), .ZN(new_n642));
  OR2_X1    g217(.A1(G99), .A2(G2105), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n643), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2096), .Z(new_n646));
  NAND3_X1  g221(.A1(new_n639), .A2(new_n640), .A3(new_n646), .ZN(G156));
  INV_X1    g222(.A(G14), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2430), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(KEYINPUT14), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g234(.A1(new_n653), .A2(KEYINPUT14), .A3(new_n657), .A4(new_n654), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n649), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n659), .A2(new_n649), .A3(new_n660), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1341), .B(G1348), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n648), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT86), .ZN(new_n667));
  AND3_X1   g242(.A1(new_n659), .A2(new_n649), .A3(new_n660), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n668), .A2(new_n661), .ZN(new_n669));
  INV_X1    g244(.A(new_n665), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n667), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NOR4_X1   g246(.A1(new_n668), .A2(new_n661), .A3(KEYINPUT86), .A4(new_n665), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n666), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G401));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2072), .B(G2078), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  OR3_X1    g253(.A1(new_n677), .A2(KEYINPUT87), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g254(.A(KEYINPUT87), .B1(new_n677), .B2(new_n678), .ZN(new_n680));
  INV_X1    g255(.A(new_n675), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n676), .B(KEYINPUT17), .Z(new_n682));
  OAI211_X1 g257(.A(new_n679), .B(new_n680), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n678), .A2(new_n675), .A3(new_n676), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT18), .Z(new_n685));
  NAND3_X1  g260(.A1(new_n682), .A2(new_n678), .A3(new_n681), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n683), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G2096), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT88), .B(G2100), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n690), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(G227));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1956), .B(G2474), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT89), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1961), .B(G1966), .Z(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1971), .B(G1976), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT19), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n698), .A2(new_n699), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n700), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n704), .A2(new_n702), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT20), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT90), .Z(new_n712));
  NAND3_X1  g287(.A1(new_n707), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n712), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n708), .B(KEYINPUT20), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n706), .ZN(new_n716));
  XOR2_X1   g291(.A(G1991), .B(G1996), .Z(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  AND3_X1   g293(.A1(new_n713), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n718), .B1(new_n713), .B2(new_n716), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n695), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n713), .A2(new_n716), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(new_n717), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n713), .A2(new_n716), .A3(new_n718), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n723), .A2(new_n694), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n721), .A2(new_n725), .ZN(G229));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G22), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G166), .B2(new_n727), .ZN(new_n729));
  INV_X1    g304(.A(G1971), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n727), .A2(G23), .ZN(new_n732));
  INV_X1    g307(.A(G288), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(new_n727), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT33), .B(G1976), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT32), .B(G1981), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n727), .B1(new_n586), .B2(new_n592), .ZN(new_n740));
  NOR2_X1   g315(.A1(G6), .A2(G16), .ZN(new_n741));
  OR3_X1    g316(.A1(new_n740), .A2(KEYINPUT93), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(KEYINPUT93), .B1(new_n740), .B2(new_n741), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n737), .B1(new_n739), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n742), .A2(new_n738), .A3(new_n743), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(KEYINPUT34), .ZN(new_n748));
  NOR2_X1   g323(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n737), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n744), .A2(new_n739), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT34), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n751), .A2(new_n752), .A3(new_n753), .A4(new_n746), .ZN(new_n754));
  INV_X1    g329(.A(G29), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G25), .ZN(new_n756));
  INV_X1    g331(.A(G107), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G2105), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n758), .B(G2104), .C1(G95), .C2(G2105), .ZN(new_n759));
  OAI211_X1 g334(.A(G119), .B(G2105), .C1(new_n473), .C2(new_n474), .ZN(new_n760));
  OAI211_X1 g335(.A(G131), .B(new_n462), .C1(new_n473), .C2(new_n474), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n759), .B(new_n760), .C1(new_n761), .C2(KEYINPUT91), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT91), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n482), .B2(G131), .ZN(new_n764));
  OAI21_X1  g339(.A(KEYINPUT92), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n760), .A2(new_n759), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT92), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n761), .A2(KEYINPUT91), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n482), .A2(new_n763), .A3(G131), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n766), .A2(new_n767), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n765), .A2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n756), .B1(new_n772), .B2(new_n755), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT35), .B(G1991), .Z(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n773), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n727), .A2(G24), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n603), .B2(new_n727), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1986), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n748), .A2(new_n750), .A3(new_n754), .A4(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n753), .B1(new_n745), .B2(new_n746), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n754), .A2(new_n780), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n749), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n727), .A2(G20), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT23), .Z(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G299), .B2(G16), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1956), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n554), .A2(G16), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G16), .B2(G19), .ZN(new_n792));
  INV_X1    g367(.A(G1341), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n793), .B2(new_n792), .ZN(new_n795));
  NOR2_X1   g370(.A1(G16), .A2(G21), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G168), .B2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT98), .B(G1966), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n461), .A2(G127), .ZN(new_n800));
  NAND2_X1  g375(.A1(G115), .A2(G2104), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n462), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT25), .ZN(new_n804));
  NAND2_X1  g379(.A1(G103), .A2(G2104), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(G2105), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n462), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n482), .A2(G139), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n803), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(KEYINPUT97), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT97), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n803), .A2(new_n811), .A3(new_n808), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n755), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n755), .A2(G33), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n755), .A2(G35), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT101), .Z(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G162), .B2(new_n755), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT102), .B(KEYINPUT29), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(G2090), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n815), .A2(G2072), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(G164), .A2(G29), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G27), .B2(G29), .ZN(new_n824));
  INV_X1    g399(.A(G2078), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT30), .B(G28), .ZN(new_n827));
  OR2_X1    g402(.A1(KEYINPUT31), .A2(G11), .ZN(new_n828));
  NAND2_X1  g403(.A1(KEYINPUT31), .A2(G11), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n827), .A2(new_n755), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n645), .B2(new_n755), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n755), .A2(G32), .ZN(new_n832));
  NAND3_X1  g407(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT26), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n484), .A2(G129), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n465), .A2(G105), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n461), .A2(new_n462), .ZN(new_n838));
  INV_X1    g413(.A(G141), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n832), .B1(new_n841), .B2(G29), .ZN(new_n842));
  XNOR2_X1  g417(.A(KEYINPUT27), .B(G1996), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n831), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n824), .A2(new_n825), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n826), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n813), .A2(G2072), .A3(new_n814), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n755), .A2(G26), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT28), .ZN(new_n849));
  INV_X1    g424(.A(G116), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n464), .B1(new_n850), .B2(G2105), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT95), .ZN(new_n852));
  NOR3_X1   g427(.A1(new_n852), .A2(G104), .A3(G2105), .ZN(new_n853));
  INV_X1    g428(.A(G104), .ZN(new_n854));
  AOI21_X1  g429(.A(KEYINPUT95), .B1(new_n854), .B2(new_n462), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n851), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n461), .A2(G140), .A3(new_n462), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n461), .A2(G128), .A3(G2105), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n849), .B1(new_n860), .B2(new_n755), .ZN(new_n861));
  XNOR2_X1  g436(.A(KEYINPUT96), .B(G2067), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n842), .B2(new_n843), .ZN(new_n865));
  NOR4_X1   g440(.A1(new_n846), .A2(new_n847), .A3(new_n863), .A4(new_n865), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n795), .A2(new_n799), .A3(new_n822), .A4(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n820), .A2(new_n821), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT103), .ZN(new_n869));
  NOR2_X1   g444(.A1(G5), .A2(G16), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT99), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(G301), .B2(new_n727), .ZN(new_n872));
  INV_X1    g447(.A(G1961), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(G1348), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n727), .A2(G4), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n876), .B1(new_n615), .B2(G16), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n874), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT24), .ZN(new_n879));
  INV_X1    g454(.A(G34), .ZN(new_n880));
  AOI21_X1  g455(.A(G29), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(new_n879), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(G160), .B2(new_n755), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n883), .A2(G2084), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT100), .ZN(new_n885));
  INV_X1    g460(.A(new_n877), .ZN(new_n886));
  AOI22_X1  g461(.A1(new_n886), .A2(G1348), .B1(G2084), .B2(new_n883), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n878), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n867), .A2(new_n869), .A3(new_n888), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n889), .A2(KEYINPUT104), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(KEYINPUT104), .ZN(new_n891));
  AOI22_X1  g466(.A1(new_n785), .A2(new_n786), .B1(new_n890), .B2(new_n891), .ZN(G311));
  NAND2_X1  g467(.A1(new_n785), .A2(new_n786), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(new_n891), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(G150));
  NAND2_X1  g470(.A1(new_n623), .A2(G559), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT105), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(KEYINPUT38), .Z(new_n898));
  INV_X1    g473(.A(G55), .ZN(new_n899));
  INV_X1    g474(.A(G93), .ZN(new_n900));
  OAI22_X1  g475(.A1(new_n535), .A2(new_n899), .B1(new_n513), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(G67), .B1(new_n506), .B2(new_n507), .ZN(new_n902));
  NAND2_X1  g477(.A1(G80), .A2(G543), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n538), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n553), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n905), .B(new_n545), .C1(new_n552), .C2(new_n550), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n898), .B(new_n909), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n910), .A2(KEYINPUT39), .ZN(new_n911));
  INV_X1    g486(.A(G860), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(KEYINPUT39), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n905), .A2(new_n912), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(KEYINPUT37), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(G145));
  INV_X1    g492(.A(KEYINPUT109), .ZN(new_n918));
  INV_X1    g493(.A(G37), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n836), .A2(new_n840), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n499), .A2(new_n497), .ZN(new_n921));
  AOI22_X1  g496(.A1(new_n484), .A2(G126), .B1(new_n490), .B2(new_n492), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n921), .A2(new_n859), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n859), .B1(new_n921), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n806), .A2(new_n807), .ZN(new_n926));
  INV_X1    g501(.A(G139), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n926), .B1(new_n838), .B2(new_n927), .ZN(new_n928));
  OAI211_X1 g503(.A(KEYINPUT97), .B(KEYINPUT106), .C1(new_n928), .C2(new_n802), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n812), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n498), .B1(new_n482), .B2(G138), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n922), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n860), .ZN(new_n934));
  NAND2_X1  g509(.A1(G164), .A2(new_n859), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n841), .A3(new_n935), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n925), .A2(new_n930), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n809), .A2(KEYINPUT106), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n938), .B1(new_n925), .B2(new_n936), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n630), .A2(new_n631), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n633), .A2(new_n634), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n632), .A2(KEYINPUT107), .A3(new_n635), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n771), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n482), .A2(G142), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n484), .A2(G130), .ZN(new_n948));
  OR2_X1    g523(.A1(G106), .A2(G2105), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n949), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n943), .A2(new_n944), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n952), .A2(new_n765), .A3(new_n770), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n946), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n951), .B1(new_n946), .B2(new_n953), .ZN(new_n955));
  OAI22_X1  g530(.A1(new_n937), .A2(new_n939), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n938), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n923), .A2(new_n924), .A3(new_n920), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n841), .B1(new_n934), .B2(new_n935), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n925), .A2(new_n930), .A3(new_n936), .ZN(new_n961));
  INV_X1    g536(.A(new_n951), .ZN(new_n962));
  INV_X1    g537(.A(new_n953), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n952), .B1(new_n765), .B2(new_n770), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n946), .A2(new_n951), .A3(new_n953), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n960), .A2(new_n961), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  XOR2_X1   g542(.A(new_n488), .B(new_n645), .Z(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(G160), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n956), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n969), .B1(new_n956), .B2(new_n967), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n919), .B(new_n970), .C1(new_n971), .C2(KEYINPUT108), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n971), .A2(KEYINPUT108), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n918), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n956), .A2(new_n967), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n975), .B1(new_n976), .B2(new_n969), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n970), .A2(new_n919), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n971), .A2(KEYINPUT108), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n977), .A2(new_n978), .A3(KEYINPUT109), .A4(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n974), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g557(.A(new_n627), .B(new_n909), .Z(new_n983));
  OR2_X1    g558(.A1(G299), .A2(new_n615), .ZN(new_n984));
  NAND2_X1  g559(.A1(G299), .A2(new_n615), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n989));
  AND2_X1   g564(.A1(G299), .A2(new_n615), .ZN(new_n990));
  NOR2_X1   g565(.A1(G299), .A2(new_n615), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT41), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT41), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n984), .A2(new_n993), .A3(new_n985), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n989), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT111), .B1(new_n986), .B2(KEYINPUT41), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n987), .A2(new_n988), .B1(new_n983), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT110), .B1(new_n983), .B2(new_n986), .ZN(new_n999));
  AOI21_X1  g574(.A(G288), .B1(new_n586), .B2(new_n592), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n586), .A2(G288), .A3(new_n592), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n603), .A2(G303), .ZN(new_n1003));
  NAND2_X1  g578(.A1(G290), .A2(G166), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n603), .B(G303), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1002), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1006), .B1(new_n1007), .B2(new_n1000), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT42), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n998), .A2(new_n999), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n998), .B2(new_n999), .ZN(new_n1012));
  OAI21_X1  g587(.A(G868), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(G868), .B2(new_n905), .ZN(G295));
  OAI21_X1  g589(.A(new_n1013), .B1(G868), .B2(new_n905), .ZN(G331));
  INV_X1    g590(.A(KEYINPUT43), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n907), .A2(G301), .A3(new_n908), .ZN(new_n1018));
  AOI21_X1  g593(.A(G301), .B1(new_n907), .B2(new_n908), .ZN(new_n1019));
  OAI21_X1  g594(.A(G286), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n909), .A2(G171), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n907), .A2(G301), .A3(new_n908), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(G168), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n992), .A2(new_n994), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1020), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n986), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1017), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n986), .ZN(new_n1028));
  NOR3_X1   g603(.A1(new_n1018), .A2(new_n1019), .A3(G286), .ZN(new_n1029));
  AOI21_X1  g604(.A(G168), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1028), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1023), .B(new_n1020), .C1(new_n995), .C2(new_n996), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(new_n1032), .A3(new_n1009), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1027), .A2(new_n1033), .A3(new_n919), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT112), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT112), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1027), .A2(new_n1033), .A3(new_n1036), .A4(new_n919), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1016), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1033), .A2(new_n919), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1009), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(KEYINPUT43), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT44), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT43), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1027), .A2(new_n1033), .A3(new_n1016), .A4(new_n919), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT44), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1043), .A2(new_n1048), .ZN(G397));
  INV_X1    g624(.A(KEYINPUT123), .ZN(new_n1050));
  INV_X1    g625(.A(G1384), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT45), .B1(new_n933), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n467), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n462), .B1(new_n475), .B2(new_n469), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(KEYINPUT69), .ZN(new_n1055));
  AOI211_X1 g630(.A(new_n468), .B(new_n462), .C1(new_n475), .C2(new_n469), .ZN(new_n1056));
  OAI211_X1 g631(.A(G40), .B(new_n1053), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1052), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT45), .ZN(new_n1059));
  NOR3_X1   g634(.A1(G164), .A2(new_n1059), .A3(G1384), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(G1966), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G40), .ZN(new_n1063));
  AOI211_X1 g638(.A(new_n1063), .B(new_n467), .C1(new_n472), .C2(new_n477), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1065));
  INV_X1    g640(.A(G2084), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT50), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n933), .A2(new_n1067), .A3(new_n1051), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .A4(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1050), .B1(new_n1062), .B2(new_n1070), .ZN(new_n1071));
  XOR2_X1   g646(.A(KEYINPUT118), .B(G8), .Z(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1060), .A2(new_n1052), .A3(new_n1057), .ZN(new_n1074));
  OAI211_X1 g649(.A(KEYINPUT123), .B(new_n1069), .C1(new_n1074), .C2(G1966), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1071), .A2(G286), .A3(new_n1073), .A4(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1071), .A2(G8), .A3(new_n1075), .ZN(new_n1078));
  NAND2_X1  g653(.A1(G286), .A2(new_n1073), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1073), .B1(new_n1062), .B2(new_n1070), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1081), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1076), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT62), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT62), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1085), .B(new_n1076), .C1(new_n1080), .C2(new_n1082), .ZN(new_n1086));
  NAND4_X1  g661(.A1(G160), .A2(G40), .A3(new_n1051), .A4(new_n933), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n575), .A2(new_n576), .A3(G1976), .A4(new_n577), .ZN(new_n1088));
  INV_X1    g663(.A(G1976), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT52), .B1(G288), .B2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1087), .A2(new_n1073), .A3(new_n1088), .A4(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n933), .A2(new_n1051), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1073), .B(new_n1088), .C1(new_n1057), .C2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT52), .ZN(new_n1094));
  INV_X1    g669(.A(G1981), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n590), .A2(new_n1095), .A3(new_n581), .A4(new_n580), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n513), .A2(new_n579), .ZN(new_n1097));
  OAI21_X1  g672(.A(G1981), .B1(new_n585), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1096), .A2(new_n1098), .A3(KEYINPUT49), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(new_n1073), .A3(new_n1087), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT49), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1091), .B(new_n1094), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1059), .B1(G164), .B2(G1384), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT113), .B(G1384), .Z(new_n1104));
  NAND3_X1  g679(.A1(new_n933), .A2(KEYINPUT45), .A3(new_n1104), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1064), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT115), .B(G1971), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1064), .A2(new_n1068), .A3(new_n1065), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1109), .A2(G2090), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1073), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n1112));
  NAND4_X1  g687(.A1(G303), .A2(new_n1112), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1113));
  AND2_X1   g688(.A1(G303), .A2(G8), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1113), .B1(new_n1114), .B2(KEYINPUT55), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1112), .B1(new_n1114), .B2(KEYINPUT55), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1102), .B1(new_n1111), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1058), .A2(new_n1105), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1107), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(KEYINPUT116), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1110), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1120), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(new_n1126), .A3(G8), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1128), .A2(G2078), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1074), .A2(new_n1129), .B1(new_n1109), .B2(new_n873), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1064), .A2(new_n1103), .A3(new_n825), .A4(new_n1105), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n1128), .ZN(new_n1132));
  AOI21_X1  g707(.A(G301), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1118), .A2(new_n1127), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1084), .A2(new_n1086), .A3(new_n1134), .ZN(new_n1135));
  XOR2_X1   g710(.A(G299), .B(KEYINPUT57), .Z(new_n1136));
  INV_X1    g711(.A(G1956), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1109), .A2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(KEYINPUT56), .B(G2072), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1058), .A2(new_n1105), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1136), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1057), .A2(new_n1092), .ZN(new_n1142));
  INV_X1    g717(.A(G2067), .ZN(new_n1143));
  AOI22_X1  g718(.A1(new_n1109), .A2(new_n875), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1144), .A2(new_n615), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1136), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1141), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT121), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(KEYINPUT121), .B(new_n1141), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1136), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1151), .B1(new_n1152), .B2(new_n1146), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1136), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1156), .A2(KEYINPUT61), .A3(new_n1141), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n615), .B1(new_n1144), .B2(KEYINPUT60), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT60), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1109), .A2(new_n875), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1087), .A2(G2067), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1158), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1153), .A2(new_n1157), .A3(new_n1163), .ZN(new_n1164));
  XOR2_X1   g739(.A(KEYINPUT58), .B(G1341), .Z(new_n1165));
  NAND2_X1  g740(.A1(new_n1087), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1166), .B1(new_n1121), .B2(G1996), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n554), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1167), .A2(new_n1169), .A3(KEYINPUT59), .A4(new_n554), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1144), .A2(KEYINPUT60), .A3(new_n615), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1149), .B(new_n1150), .C1(new_n1164), .C2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT54), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1109), .A2(new_n873), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n933), .A2(new_n1104), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n1059), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1129), .A2(G40), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n467), .A2(new_n1054), .A3(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1179), .A2(new_n1105), .A3(new_n1181), .ZN(new_n1182));
  AND4_X1   g757(.A1(G301), .A2(new_n1132), .A3(new_n1177), .A4(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1176), .B1(new_n1133), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT124), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  OAI211_X1 g761(.A(KEYINPUT124), .B(new_n1176), .C1(new_n1133), .C2(new_n1183), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1118), .A2(new_n1127), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1058), .A2(new_n1061), .A3(new_n1129), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1132), .A2(new_n1177), .A3(new_n1190), .A4(G301), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(KEYINPUT54), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1132), .A2(new_n1177), .A3(new_n1182), .ZN(new_n1193));
  OR2_X1    g768(.A1(new_n1193), .A2(KEYINPUT125), .ZN(new_n1194));
  AOI21_X1  g769(.A(G301), .B1(new_n1193), .B2(KEYINPUT125), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1192), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1189), .A2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1175), .A2(new_n1083), .A3(new_n1188), .A4(new_n1197), .ZN(new_n1198));
  OAI211_X1 g773(.A(new_n1089), .B(new_n733), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1199));
  XOR2_X1   g774(.A(new_n1096), .B(KEYINPUT120), .Z(new_n1200));
  NAND2_X1  g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1201), .A2(new_n1073), .A3(new_n1087), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT119), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1102), .B(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1202), .B1(new_n1204), .B2(new_n1127), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT63), .ZN(new_n1206));
  OR2_X1    g781(.A1(new_n1081), .A2(G286), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1206), .B1(new_n1189), .B2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1102), .B(KEYINPUT119), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1125), .A2(G8), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1210), .A2(new_n1117), .ZN(new_n1211));
  NOR3_X1   g786(.A1(new_n1081), .A2(new_n1206), .A3(G286), .ZN(new_n1212));
  NAND4_X1  g787(.A1(new_n1209), .A2(new_n1211), .A3(new_n1127), .A4(new_n1212), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1205), .B1(new_n1208), .B2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g789(.A1(new_n1135), .A2(new_n1198), .A3(new_n1214), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n1179), .A2(new_n1057), .ZN(new_n1216));
  OR2_X1    g791(.A1(new_n1216), .A2(KEYINPUT114), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1216), .A2(KEYINPUT114), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g794(.A(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g795(.A(new_n920), .B(G1996), .ZN(new_n1221));
  XNOR2_X1  g796(.A(new_n859), .B(new_n1143), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g798(.A1(new_n771), .A2(new_n775), .ZN(new_n1224));
  NOR2_X1   g799(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g800(.A(new_n1225), .B1(new_n774), .B2(new_n772), .ZN(new_n1226));
  XOR2_X1   g801(.A(new_n603), .B(G1986), .Z(new_n1227));
  OAI21_X1  g802(.A(new_n1220), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1215), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1220), .A2(new_n1223), .ZN(new_n1230));
  AOI22_X1  g805(.A1(new_n1230), .A2(new_n1224), .B1(new_n1143), .B2(new_n860), .ZN(new_n1231));
  INV_X1    g806(.A(KEYINPUT126), .ZN(new_n1232));
  OAI21_X1  g807(.A(new_n1220), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g808(.A(new_n1233), .B1(new_n1232), .B2(new_n1231), .ZN(new_n1234));
  AOI21_X1  g809(.A(new_n1219), .B1(new_n920), .B2(new_n1222), .ZN(new_n1235));
  INV_X1    g810(.A(KEYINPUT46), .ZN(new_n1236));
  INV_X1    g811(.A(G1996), .ZN(new_n1237));
  NAND3_X1  g812(.A1(new_n1220), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  OAI21_X1  g813(.A(KEYINPUT46), .B1(new_n1219), .B2(G1996), .ZN(new_n1239));
  AOI21_X1  g814(.A(new_n1235), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  XNOR2_X1  g815(.A(new_n1240), .B(KEYINPUT47), .ZN(new_n1241));
  OR3_X1    g816(.A1(new_n1219), .A2(G1986), .A3(G290), .ZN(new_n1242));
  INV_X1    g817(.A(KEYINPUT48), .ZN(new_n1243));
  OR2_X1    g818(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g819(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1245));
  NAND2_X1  g820(.A1(new_n1220), .A2(new_n1226), .ZN(new_n1246));
  AND3_X1   g821(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  NOR3_X1   g822(.A1(new_n1234), .A2(new_n1241), .A3(new_n1247), .ZN(new_n1248));
  NAND2_X1  g823(.A1(new_n1229), .A2(new_n1248), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g824(.A(new_n459), .B1(new_n691), .B2(new_n692), .ZN(new_n1251));
  NAND4_X1  g825(.A1(new_n673), .A2(new_n1251), .A3(new_n721), .A4(new_n725), .ZN(new_n1252));
  AOI21_X1  g826(.A(new_n1252), .B1(new_n974), .B2(new_n980), .ZN(new_n1253));
  AND3_X1   g827(.A1(new_n1253), .A2(new_n1046), .A3(KEYINPUT127), .ZN(new_n1254));
  AOI21_X1  g828(.A(KEYINPUT127), .B1(new_n1253), .B2(new_n1046), .ZN(new_n1255));
  NOR2_X1   g829(.A1(new_n1254), .A2(new_n1255), .ZN(G308));
  NAND2_X1  g830(.A1(new_n1253), .A2(new_n1046), .ZN(new_n1257));
  INV_X1    g831(.A(KEYINPUT127), .ZN(new_n1258));
  NAND2_X1  g832(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g833(.A1(new_n1253), .A2(new_n1046), .A3(KEYINPUT127), .ZN(new_n1260));
  NAND2_X1  g834(.A1(new_n1259), .A2(new_n1260), .ZN(G225));
endmodule


