//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976;
  INV_X1    g000(.A(KEYINPUT34), .ZN(new_n202));
  INV_X1    g001(.A(G227gat), .ZN(new_n203));
  INV_X1    g002(.A(G233gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT69), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(G113gat), .B2(G120gat), .ZN(new_n208));
  AND2_X1   g007(.A1(G113gat), .A2(G120gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G127gat), .B(G134gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n211), .B(new_n206), .C1(new_n209), .C2(new_n208), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT28), .ZN(new_n216));
  XNOR2_X1  g015(.A(KEYINPUT27), .B(G183gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT67), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT67), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT27), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(G183gat), .ZN(new_n221));
  INV_X1    g020(.A(G183gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(KEYINPUT27), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n219), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n218), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G190gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n216), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT26), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT26), .ZN(new_n232));
  AND3_X1   g031(.A1(new_n229), .A2(KEYINPUT68), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT68), .B1(new_n229), .B2(new_n232), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n228), .B(new_n231), .C1(new_n233), .C2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT27), .B1(new_n237), .B2(new_n222), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n220), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n238), .A2(new_n239), .A3(new_n216), .A4(new_n226), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n235), .A2(new_n236), .A3(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n227), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n222), .A2(new_n226), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT24), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n236), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n245), .A2(new_n246), .A3(new_n248), .A4(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT25), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT23), .ZN(new_n252));
  NOR3_X1   g051(.A1(new_n252), .A2(G169gat), .A3(G176gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n228), .A2(KEYINPUT23), .ZN(new_n254));
  AOI211_X1 g053(.A(new_n251), .B(new_n253), .C1(new_n230), .C2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NOR3_X1   g056(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n243), .B(new_n248), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n253), .B1(new_n230), .B2(new_n254), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n250), .A2(new_n255), .B1(new_n261), .B2(new_n251), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n215), .B1(new_n242), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n251), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n260), .A2(new_n250), .A3(KEYINPUT25), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n240), .A2(new_n236), .ZN(new_n267));
  AOI21_X1  g066(.A(G190gat), .B1(new_n218), .B2(new_n224), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n267), .B(new_n235), .C1(new_n268), .C2(new_n216), .ZN(new_n269));
  INV_X1    g068(.A(new_n215), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n266), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n205), .B1(new_n263), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n202), .B1(new_n272), .B2(KEYINPUT71), .ZN(new_n273));
  INV_X1    g072(.A(new_n205), .ZN(new_n274));
  INV_X1    g073(.A(new_n271), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n270), .B1(new_n266), .B2(new_n269), .ZN(new_n276));
  OAI211_X1 g075(.A(KEYINPUT71), .B(new_n274), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n277), .A2(KEYINPUT72), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n279), .B1(new_n272), .B2(KEYINPUT71), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n273), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT34), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n272), .A2(KEYINPUT71), .A3(new_n279), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n277), .A2(KEYINPUT72), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT32), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n263), .A2(new_n205), .A3(new_n271), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT70), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT70), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n263), .A2(new_n292), .A3(new_n205), .A4(new_n271), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n289), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT33), .B1(new_n291), .B2(new_n293), .ZN(new_n295));
  XOR2_X1   g094(.A(G15gat), .B(G43gat), .Z(new_n296));
  XNOR2_X1  g095(.A(G71gat), .B(G99gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NOR3_X1   g098(.A1(new_n294), .A2(new_n295), .A3(new_n299), .ZN(new_n300));
  AOI221_X4 g099(.A(new_n289), .B1(KEYINPUT33), .B2(new_n298), .C1(new_n291), .C2(new_n293), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n288), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n291), .A2(new_n293), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT33), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n299), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n294), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n301), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n307), .A2(new_n308), .A3(new_n287), .A4(new_n281), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n302), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT36), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n307), .A2(new_n308), .B1(new_n287), .B2(new_n281), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(KEYINPUT73), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n314), .B1(new_n310), .B2(KEYINPUT73), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT36), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n312), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G78gat), .B(G106gat), .ZN(new_n318));
  INV_X1    g117(.A(G50gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n320), .B(G22gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G211gat), .B(G218gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(G197gat), .B(G204gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT22), .ZN(new_n325));
  INV_X1    g124(.A(G211gat), .ZN(new_n326));
  INV_X1    g125(.A(G218gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n323), .A2(new_n324), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n323), .B1(new_n328), .B2(new_n324), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G141gat), .ZN(new_n334));
  INV_X1    g133(.A(G148gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G141gat), .A2(G148gat), .ZN(new_n337));
  AND2_X1   g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n336), .B(new_n337), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT2), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT76), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  AND2_X1   g143(.A1(G141gat), .A2(G148gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(G141gat), .A2(G148gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G155gat), .B(G162gat), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .A4(new_n342), .ZN(new_n350));
  INV_X1    g149(.A(new_n348), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n342), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n341), .A2(KEYINPUT75), .A3(KEYINPUT2), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n353), .A2(new_n354), .A3(new_n347), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n344), .A2(new_n350), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT3), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT29), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n333), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n356), .ZN(new_n362));
  INV_X1    g161(.A(new_n331), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT29), .B1(new_n363), .B2(new_n329), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT82), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n357), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n359), .B1(new_n330), .B2(new_n331), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n367), .A2(KEYINPUT82), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n362), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G228gat), .A2(G233gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n361), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT83), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT3), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n364), .A2(KEYINPUT83), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n356), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI211_X1 g174(.A(G228gat), .B(G233gat), .C1(new_n375), .C2(new_n360), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n371), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n378), .B1(new_n371), .B2(new_n376), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n322), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n371), .A2(new_n376), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n377), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n371), .A2(new_n376), .A3(new_n378), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n321), .A3(new_n384), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G226gat), .A2(G233gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n266), .A2(new_n269), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n388), .B1(new_n389), .B2(new_n359), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n225), .A2(new_n226), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT28), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n228), .B1(new_n229), .B2(new_n232), .ZN(new_n393));
  INV_X1    g192(.A(new_n234), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n229), .A2(KEYINPUT68), .A3(new_n232), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n240), .A2(new_n236), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n392), .A2(new_n398), .B1(new_n264), .B2(new_n265), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n399), .A2(new_n387), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n390), .A2(new_n400), .A3(new_n332), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT74), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n402), .B1(new_n399), .B2(new_n387), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n389), .A2(KEYINPUT74), .A3(new_n388), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n387), .B1(new_n399), .B2(KEYINPUT29), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n401), .B1(new_n407), .B2(new_n332), .ZN(new_n408));
  XNOR2_X1  g207(.A(G8gat), .B(G36gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(G64gat), .B(G92gat), .ZN(new_n410));
  XOR2_X1   g209(.A(new_n409), .B(new_n410), .Z(new_n411));
  NAND2_X1  g210(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT30), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n389), .A2(new_n388), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n406), .A2(new_n333), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n390), .B1(new_n403), .B2(new_n404), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n416), .B1(new_n417), .B2(new_n333), .ZN(new_n418));
  INV_X1    g217(.A(new_n411), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n408), .A2(KEYINPUT30), .A3(new_n411), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n414), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n270), .B1(new_n356), .B2(new_n357), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n344), .A2(new_n350), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n355), .A2(new_n351), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n424), .A2(new_n357), .A3(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(new_n425), .A3(new_n215), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n356), .A2(KEYINPUT4), .A3(new_n215), .ZN(new_n432));
  NAND2_X1  g231(.A1(G225gat), .A2(G233gat), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n428), .A2(new_n431), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT5), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n356), .B(new_n215), .ZN(new_n436));
  INV_X1    g235(.A(new_n433), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT78), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n431), .A2(KEYINPUT77), .A3(new_n432), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT77), .B1(new_n431), .B2(new_n432), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n435), .B(new_n433), .C1(new_n423), .C2(new_n426), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n440), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT77), .ZN(new_n447));
  AND4_X1   g246(.A1(KEYINPUT4), .A2(new_n424), .A3(new_n425), .A4(new_n215), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT4), .B1(new_n356), .B2(new_n215), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n431), .A2(KEYINPUT77), .A3(new_n432), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n452), .A2(KEYINPUT78), .A3(new_n444), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n439), .B1(new_n446), .B2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(G1gat), .B(G29gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(KEYINPUT0), .ZN(new_n456));
  XNOR2_X1  g255(.A(G57gat), .B(G85gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT78), .B1(new_n452), .B2(new_n444), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n445), .A2(new_n440), .A3(new_n450), .A4(new_n451), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n458), .B1(new_n434), .B2(new_n438), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n464), .A2(KEYINPUT79), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT79), .B1(new_n464), .B2(new_n465), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n459), .B(new_n460), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT80), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n461), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT6), .B1(new_n454), .B2(new_n458), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n471), .B(KEYINPUT80), .C1(new_n467), .C2(new_n466), .ZN(new_n472));
  AOI211_X1 g271(.A(new_n386), .B(new_n422), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n386), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT38), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT37), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n411), .B1(new_n408), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n418), .A2(KEYINPUT37), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n419), .B1(new_n418), .B2(KEYINPUT37), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n417), .A2(new_n332), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n406), .A2(new_n332), .A3(new_n415), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT37), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n475), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n412), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n461), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n458), .B(KEYINPUT84), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n454), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n489), .B(new_n460), .C1(new_n466), .C2(new_n467), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n486), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n437), .B1(new_n452), .B2(new_n427), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n436), .A2(new_n437), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT39), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n488), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(KEYINPUT85), .B(KEYINPUT39), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n437), .B(new_n497), .C1(new_n452), .C2(new_n427), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT86), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n499), .A2(KEYINPUT40), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n499), .A2(KEYINPUT40), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n489), .B(new_n422), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n474), .B1(new_n491), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n317), .B1(new_n473), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n490), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT35), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n381), .A2(new_n385), .A3(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n422), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n315), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n302), .A2(new_n309), .A3(new_n386), .ZN(new_n511));
  AOI211_X1 g310(.A(new_n422), .B(new_n511), .C1(new_n470), .C2(new_n472), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n510), .B1(new_n512), .B2(new_n506), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n504), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G57gat), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT95), .B1(new_n515), .B2(G64gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT95), .ZN(new_n517));
  INV_X1    g316(.A(G64gat), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(new_n518), .A3(G57gat), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n516), .B(new_n519), .C1(G57gat), .C2(new_n518), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT96), .ZN(new_n521));
  NAND2_X1  g320(.A1(G71gat), .A2(G78gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(G71gat), .A2(G78gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT9), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n520), .A2(new_n521), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(new_n521), .B2(new_n520), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT94), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n523), .B1(new_n527), .B2(new_n522), .ZN(new_n528));
  XNOR2_X1  g327(.A(G57gat), .B(G64gat), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n527), .A2(KEYINPUT9), .ZN(new_n530));
  OAI221_X1 g329(.A(new_n528), .B1(new_n527), .B2(new_n522), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT21), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(G231gat), .A2(G233gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(G127gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G15gat), .B(G22gat), .ZN(new_n539));
  INV_X1    g338(.A(G1gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT16), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n542), .B1(G1gat), .B2(new_n539), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(G8gat), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(new_n533), .B2(new_n532), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n538), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G183gat), .B(G211gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT97), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n550));
  INV_X1    g349(.A(G155gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n549), .B(new_n552), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n547), .A2(new_n553), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G113gat), .B(G141gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(G197gat), .ZN(new_n559));
  XOR2_X1   g358(.A(KEYINPUT11), .B(G169gat), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n561), .B(KEYINPUT12), .Z(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G229gat), .A2(G233gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT14), .B(G29gat), .ZN(new_n565));
  INV_X1    g364(.A(G36gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(G29gat), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n319), .A2(G43gat), .ZN(new_n571));
  INV_X1    g370(.A(G43gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(G50gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT87), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT15), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n573), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n576), .B1(new_n577), .B2(KEYINPUT87), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n570), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT89), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n573), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n571), .A2(KEYINPUT88), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n572), .A2(KEYINPUT89), .A3(G50gat), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT88), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n584), .A2(new_n319), .A3(G43gat), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n581), .A2(new_n582), .A3(new_n583), .A4(new_n585), .ZN(new_n586));
  AOI22_X1  g385(.A1(new_n586), .A2(new_n576), .B1(new_n567), .B2(new_n569), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n578), .A2(new_n575), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n579), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n545), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT17), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n591), .B(new_n579), .C1(new_n587), .C2(new_n588), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT90), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n544), .B1(KEYINPUT17), .B2(new_n589), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n564), .B(new_n590), .C1(new_n593), .C2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT18), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT92), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n545), .A2(new_n589), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT90), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n592), .B(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n599), .B1(new_n601), .B2(new_n594), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT92), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n602), .A2(new_n603), .A3(KEYINPUT18), .A4(new_n564), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n598), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(new_n564), .B(KEYINPUT13), .Z(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n545), .A2(new_n589), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n607), .B1(new_n590), .B2(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(KEYINPUT91), .B(KEYINPUT18), .Z(new_n610));
  AOI21_X1  g409(.A(new_n609), .B1(new_n596), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n563), .B1(new_n605), .B2(new_n611), .ZN(new_n612));
  AOI211_X1 g411(.A(new_n562), .B(new_n609), .C1(new_n596), .C2(new_n610), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n605), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(KEYINPUT93), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT93), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n605), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n612), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(G85gat), .A2(G92gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT7), .ZN(new_n621));
  NAND2_X1  g420(.A1(G99gat), .A2(G106gat), .ZN(new_n622));
  INV_X1    g421(.A(G85gat), .ZN(new_n623));
  INV_X1    g422(.A(G92gat), .ZN(new_n624));
  AOI22_X1  g423(.A1(KEYINPUT8), .A2(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G99gat), .B(G106gat), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n626), .B(new_n627), .Z(new_n628));
  OAI21_X1  g427(.A(new_n619), .B1(new_n628), .B2(new_n589), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n626), .B(new_n627), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n630), .B1(new_n589), .B2(KEYINPUT17), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n629), .B1(new_n601), .B2(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G190gat), .B(G218gat), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n635), .B(KEYINPUT98), .Z(new_n636));
  XNOR2_X1  g435(.A(G134gat), .B(G162gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n633), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n632), .B(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n638), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G230gat), .A2(G233gat), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n532), .A2(new_n628), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT10), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n630), .A2(new_n526), .A3(new_n531), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n630), .A2(KEYINPUT10), .A3(new_n526), .A4(new_n531), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n646), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n645), .B1(new_n647), .B2(new_n649), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT99), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT99), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n654), .A2(new_n660), .A3(new_n657), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n657), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n663), .B1(new_n652), .B2(new_n653), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NOR4_X1   g464(.A1(new_n557), .A2(new_n618), .A3(new_n644), .A4(new_n665), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n514), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n468), .A2(new_n469), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n668), .A2(new_n472), .A3(new_n487), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g471(.A1(new_n667), .A2(new_n422), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT16), .B(G8gat), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(KEYINPUT42), .Z(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(G8gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT100), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(G1325gat));
  INV_X1    g478(.A(new_n667), .ZN(new_n680));
  OAI21_X1  g479(.A(G15gat), .B1(new_n680), .B2(new_n317), .ZN(new_n681));
  INV_X1    g480(.A(new_n315), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(G15gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n681), .B1(new_n680), .B2(new_n683), .ZN(G1326gat));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n474), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT101), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT43), .B(G22gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  INV_X1    g487(.A(new_n644), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n689), .B1(new_n504), .B2(new_n513), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n556), .A2(new_n618), .A3(new_n665), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n692), .A2(G29gat), .A3(new_n669), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT45), .Z(new_n694));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n300), .A2(new_n288), .A3(new_n301), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT73), .B1(new_n696), .B2(new_n313), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT73), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n302), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n697), .A2(new_n316), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n311), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n491), .A2(new_n502), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n386), .ZN(new_n703));
  INV_X1    g502(.A(new_n422), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n669), .A2(new_n474), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n701), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n511), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n669), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n708), .A2(KEYINPUT35), .B1(new_n315), .B2(new_n509), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n695), .B(new_n644), .C1(new_n706), .C2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(KEYINPUT102), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT102), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n713), .B1(new_n690), .B2(new_n695), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n713), .B(new_n644), .C1(new_n706), .C2(new_n709), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT44), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n691), .B(new_n712), .C1(new_n714), .C2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G29gat), .B1(new_n717), .B2(new_n669), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n694), .A2(new_n718), .ZN(G1328gat));
  AND4_X1   g518(.A1(new_n566), .A2(new_n690), .A3(new_n422), .A4(new_n691), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT46), .ZN(new_n721));
  OAI21_X1  g520(.A(G36gat), .B1(new_n717), .B2(new_n704), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT104), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n721), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(G1329gat));
  INV_X1    g526(.A(KEYINPUT47), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n682), .A2(G43gat), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  OR3_X1    g529(.A1(new_n692), .A2(KEYINPUT105), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT105), .B1(new_n692), .B2(new_n730), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n728), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT106), .B1(new_n717), .B2(new_n317), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(G43gat), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n717), .A2(KEYINPUT106), .A3(new_n317), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n733), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(G43gat), .B1(new_n717), .B2(new_n317), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n731), .A2(new_n732), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n728), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n737), .A2(new_n741), .ZN(G1330gat));
  OAI21_X1  g541(.A(new_n319), .B1(new_n692), .B2(new_n386), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n474), .A2(G50gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n717), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g545(.A(new_n618), .ZN(new_n747));
  INV_X1    g546(.A(new_n665), .ZN(new_n748));
  NOR4_X1   g547(.A1(new_n557), .A2(new_n747), .A3(new_n644), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n514), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n670), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G57gat), .ZN(G1332gat));
  INV_X1    g552(.A(KEYINPUT49), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n422), .B1(new_n754), .B2(new_n518), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT107), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n518), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1333gat));
  OAI21_X1  g558(.A(G71gat), .B1(new_n750), .B2(new_n317), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n682), .A2(G71gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n750), .B2(new_n761), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g562(.A1(new_n751), .A2(new_n474), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g564(.A1(new_n556), .A2(new_n747), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(new_n748), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n712), .B(new_n768), .C1(new_n714), .C2(new_n716), .ZN(new_n769));
  OAI21_X1  g568(.A(G85gat), .B1(new_n769), .B2(new_n669), .ZN(new_n770));
  INV_X1    g569(.A(new_n690), .ZN(new_n771));
  OR3_X1    g570(.A1(new_n771), .A2(KEYINPUT51), .A3(new_n767), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT51), .B1(new_n771), .B2(new_n767), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n772), .A2(new_n665), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n670), .A2(new_n623), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n770), .B1(new_n774), .B2(new_n775), .ZN(G1336gat));
  OAI21_X1  g575(.A(G92gat), .B1(new_n769), .B2(new_n704), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n422), .A2(new_n624), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n774), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT52), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n777), .B(new_n781), .C1(new_n774), .C2(new_n778), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(G1337gat));
  OAI21_X1  g582(.A(G99gat), .B1(new_n769), .B2(new_n317), .ZN(new_n784));
  OR2_X1    g583(.A1(new_n682), .A2(G99gat), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n774), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT108), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT108), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n784), .B(new_n788), .C1(new_n774), .C2(new_n785), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(G1338gat));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  OAI21_X1  g590(.A(G106gat), .B1(new_n769), .B2(new_n386), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n791), .B1(new_n792), .B2(KEYINPUT109), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n386), .A2(G106gat), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n792), .B1(new_n774), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  OAI221_X1 g596(.A(new_n792), .B1(KEYINPUT109), .B2(new_n791), .C1(new_n774), .C2(new_n795), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(G1339gat));
  NAND4_X1  g598(.A1(new_n556), .A2(new_n618), .A3(new_n689), .A4(new_n748), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n650), .A2(new_n651), .A3(new_n646), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n802), .A2(new_n652), .A3(new_n803), .ZN(new_n804));
  XOR2_X1   g603(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n805));
  NAND2_X1  g604(.A1(new_n652), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n663), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  AOI22_X1  g607(.A1(KEYINPUT55), .A2(new_n808), .B1(new_n659), .B2(new_n661), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n810), .B1(new_n804), .B2(new_n807), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n809), .A2(new_n644), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(new_n602), .B2(new_n564), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n590), .A2(new_n608), .A3(new_n607), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n602), .A2(new_n813), .A3(new_n564), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n561), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n605), .A2(new_n613), .A3(new_n616), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n616), .B1(new_n605), .B2(new_n613), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n812), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n665), .B(new_n818), .C1(new_n820), .C2(new_n819), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n809), .A2(new_n811), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n823), .B1(new_n618), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n822), .B1(new_n825), .B2(new_n689), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n800), .B1(new_n826), .B2(new_n556), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n827), .A2(new_n670), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n828), .A2(new_n704), .A3(new_n707), .ZN(new_n829));
  AOI21_X1  g628(.A(G113gat), .B1(new_n829), .B2(new_n747), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n827), .A2(new_n315), .A3(new_n386), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n670), .A3(new_n704), .ZN(new_n832));
  INV_X1    g631(.A(G113gat), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n832), .A2(new_n833), .A3(new_n618), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n830), .A2(new_n834), .ZN(G1340gat));
  AOI21_X1  g634(.A(G120gat), .B1(new_n829), .B2(new_n665), .ZN(new_n836));
  INV_X1    g635(.A(G120gat), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n832), .A2(new_n837), .A3(new_n748), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n836), .A2(new_n838), .ZN(G1341gat));
  NAND3_X1  g638(.A1(new_n829), .A2(new_n537), .A3(new_n556), .ZN(new_n840));
  OAI21_X1  g639(.A(G127gat), .B1(new_n832), .B2(new_n557), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XOR2_X1   g641(.A(new_n842), .B(KEYINPUT112), .Z(G1342gat));
  OAI21_X1  g642(.A(G134gat), .B1(new_n832), .B2(new_n689), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n689), .A2(new_n422), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT113), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(G134gat), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n828), .A2(new_n707), .A3(new_n847), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n848), .A2(KEYINPUT56), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(KEYINPUT56), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n844), .A2(new_n849), .A3(new_n850), .ZN(G1343gat));
  NOR2_X1   g650(.A1(new_n701), .A2(new_n386), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n828), .A2(new_n704), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n334), .B1(new_n853), .B2(new_n618), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n701), .A2(new_n669), .A3(new_n422), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n856), .B1(new_n804), .B2(new_n807), .ZN(new_n857));
  INV_X1    g656(.A(new_n652), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(KEYINPUT54), .A3(new_n801), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n859), .A2(KEYINPUT115), .A3(new_n663), .A4(new_n806), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n857), .A2(new_n810), .A3(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n857), .A2(new_n860), .A3(KEYINPUT116), .A4(new_n810), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n809), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n823), .B1(new_n865), .B2(new_n618), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n822), .B1(new_n866), .B2(new_n689), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n800), .B1(new_n867), .B2(new_n556), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(KEYINPUT57), .A3(new_n474), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT57), .B1(new_n827), .B2(new_n474), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI211_X1 g671(.A(KEYINPUT114), .B(KEYINPUT57), .C1(new_n827), .C2(new_n474), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n855), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n747), .A2(G141gat), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n854), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT58), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT58), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n876), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(G1344gat));
  NOR3_X1   g681(.A1(new_n853), .A2(G148gat), .A3(new_n748), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n665), .B(new_n855), .C1(new_n872), .C2(new_n873), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n335), .A2(KEYINPUT59), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n855), .A2(new_n665), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT57), .B1(new_n868), .B2(new_n474), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n827), .A2(KEYINPUT57), .A3(new_n474), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G148gat), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n892), .A2(KEYINPUT59), .ZN(new_n893));
  OAI211_X1 g692(.A(KEYINPUT118), .B(new_n884), .C1(new_n887), .C2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n895));
  AOI22_X1  g694(.A1(new_n885), .A2(new_n886), .B1(new_n892), .B2(KEYINPUT59), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(new_n883), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n894), .A2(new_n897), .ZN(G1345gat));
  NOR3_X1   g697(.A1(new_n874), .A2(new_n551), .A3(new_n557), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n853), .A2(new_n557), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(KEYINPUT119), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(G155gat), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(KEYINPUT119), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(G1346gat));
  NOR2_X1   g703(.A1(new_n846), .A2(G162gat), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n828), .A2(new_n852), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT120), .B1(new_n874), .B2(new_n689), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(G162gat), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n874), .A2(KEYINPUT120), .A3(new_n689), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(G1347gat));
  NOR2_X1   g709(.A1(new_n670), .A2(new_n704), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n831), .A2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(G169gat), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n912), .A2(new_n913), .A3(new_n618), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n827), .A2(new_n669), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(new_n422), .A3(new_n707), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n747), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n914), .B1(new_n913), .B2(new_n918), .ZN(G1348gat));
  OR3_X1    g718(.A1(new_n916), .A2(G176gat), .A3(new_n748), .ZN(new_n920));
  OAI21_X1  g719(.A(G176gat), .B1(new_n912), .B2(new_n748), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1349gat));
  OR3_X1    g721(.A1(new_n912), .A2(KEYINPUT121), .A3(new_n557), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT121), .B1(new_n912), .B2(new_n557), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n923), .A2(G183gat), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n917), .A2(new_n225), .A3(new_n556), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT60), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n925), .A2(new_n929), .A3(new_n926), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1350gat));
  OAI21_X1  g730(.A(G190gat), .B1(new_n912), .B2(new_n689), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n932), .A2(KEYINPUT122), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n226), .A3(new_n644), .ZN(new_n935));
  XOR2_X1   g734(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n936));
  OAI211_X1 g735(.A(new_n934), .B(new_n935), .C1(new_n932), .C2(new_n936), .ZN(G1351gat));
  NOR3_X1   g736(.A1(new_n701), .A2(new_n386), .A3(new_n704), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n915), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT123), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n939), .B(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(G197gat), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n941), .A2(new_n942), .A3(new_n747), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n911), .A2(new_n317), .A3(new_n747), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n868), .A2(new_n474), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT57), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n827), .A2(KEYINPUT57), .A3(new_n474), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT124), .ZN(new_n950));
  OR3_X1    g749(.A1(new_n889), .A2(new_n890), .A3(KEYINPUT124), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n944), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT125), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(G197gat), .B1(new_n952), .B2(new_n953), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n943), .B1(new_n954), .B2(new_n955), .ZN(G1352gat));
  AOI21_X1  g755(.A(G204gat), .B1(KEYINPUT126), .B2(KEYINPUT62), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n915), .A2(new_n665), .A3(new_n938), .A4(new_n957), .ZN(new_n958));
  NOR2_X1   g757(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n958), .B(new_n959), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n950), .A2(new_n951), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n911), .A2(new_n317), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n961), .A2(new_n748), .A3(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(G204gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n960), .B1(new_n963), .B2(new_n964), .ZN(G1353gat));
  NOR2_X1   g764(.A1(new_n962), .A2(new_n557), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n326), .B1(new_n949), .B2(new_n966), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n967), .B(KEYINPUT63), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n557), .A2(G211gat), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n941), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n969), .B1(new_n941), .B2(new_n970), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(G1354gat));
  AOI21_X1  g772(.A(G218gat), .B1(new_n941), .B2(new_n644), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n961), .A2(new_n962), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n689), .A2(new_n327), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(G1355gat));
endmodule


