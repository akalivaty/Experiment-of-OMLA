//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XOR2_X1   g0002(.A(new_n202), .B(KEYINPUT64), .Z(G355));
  NAND2_X1  g0003(.A1(G1), .A2(G20), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT65), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  INV_X1    g0009(.A(KEYINPUT1), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n211));
  INV_X1    g0011(.A(G50), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G116), .ZN(new_n214));
  INV_X1    g0014(.A(G270), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT66), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(new_n216), .A2(new_n217), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G97), .A2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G58), .A2(G232), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n206), .B1(KEYINPUT67), .B2(new_n210), .C1(new_n222), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n210), .A2(KEYINPUT67), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(G58), .A2(G68), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n209), .B(new_n228), .C1(new_n231), .C2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n215), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  INV_X1    g0045(.A(G107), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n214), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G68), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT68), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT68), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G41), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT5), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n254), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G45), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G1), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n253), .A2(KEYINPUT5), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT69), .ZN(new_n263));
  AND2_X1   g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n263), .B1(new_n264), .B2(new_n229), .ZN(new_n265));
  AND2_X1   g0065(.A1(G1), .A2(G13), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(KEYINPUT69), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n262), .A2(G264), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n224), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(G257), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G1698), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n272), .A2(new_n274), .A3(new_n276), .A4(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G294), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n264), .A2(new_n229), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT88), .ZN(new_n284));
  AND3_X1   g0084(.A1(new_n270), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n284), .B1(new_n270), .B2(new_n283), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n261), .A2(G274), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NOR3_X1   g0088(.A1(new_n264), .A2(new_n263), .A3(new_n229), .ZN(new_n289));
  AOI21_X1  g0089(.A(KEYINPUT69), .B1(new_n266), .B2(new_n267), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n258), .A2(new_n260), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT82), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n258), .A2(KEYINPUT82), .A3(new_n260), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n291), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n285), .A2(new_n286), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n287), .B1(new_n265), .B2(new_n268), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n258), .A2(KEYINPUT82), .A3(new_n260), .ZN(new_n299));
  AOI21_X1  g0099(.A(KEYINPUT82), .B1(new_n258), .B2(new_n260), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(new_n283), .A3(new_n270), .ZN(new_n302));
  OAI22_X1  g0102(.A1(new_n297), .A2(G200), .B1(G190), .B2(new_n302), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n274), .A2(new_n276), .A3(new_n230), .A4(G87), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT22), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT3), .B(G33), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n307), .A2(KEYINPUT22), .A3(new_n230), .A4(G87), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  AND2_X1   g0110(.A1(KEYINPUT72), .A2(G107), .ZN(new_n311));
  NOR2_X1   g0111(.A1(KEYINPUT72), .A2(G107), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT23), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT23), .B1(new_n246), .B2(G20), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G20), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G33), .A2(G116), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n310), .A2(new_n320), .A3(KEYINPUT24), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT24), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n316), .A2(G20), .B1(new_n314), .B2(new_n318), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(new_n309), .ZN(new_n324));
  NAND3_X1  g0124(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n229), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n321), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n325), .A2(new_n229), .ZN(new_n328));
  INV_X1    g0128(.A(G1), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G33), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(G13), .A3(G20), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n328), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G107), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n331), .A2(G107), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n334), .B(KEYINPUT25), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n327), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n303), .A2(KEYINPUT90), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT90), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n270), .A2(new_n283), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n339), .A2(new_n296), .A3(G190), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(KEYINPUT88), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n270), .A2(new_n283), .A3(new_n284), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n341), .A2(new_n301), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G200), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n340), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n327), .A2(new_n333), .A3(new_n335), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n338), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT89), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n297), .A2(new_n348), .A3(G179), .ZN(new_n349));
  INV_X1    g0149(.A(G179), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT89), .B1(new_n343), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n302), .A2(G169), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n337), .A2(new_n347), .B1(new_n353), .B2(new_n346), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT71), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n328), .A2(new_n355), .B1(G1), .B2(new_n230), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n356), .B1(new_n355), .B2(new_n328), .ZN(new_n357));
  OAI21_X1  g0157(.A(G20), .B1(new_n233), .B2(G50), .ZN(new_n358));
  INV_X1    g0158(.A(G150), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n230), .A2(new_n273), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n230), .A2(G33), .ZN(new_n361));
  XNOR2_X1  g0161(.A(KEYINPUT8), .B(G58), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n358), .B1(new_n359), .B2(new_n360), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n357), .A2(G50), .B1(new_n363), .B2(new_n326), .ZN(new_n364));
  INV_X1    g0164(.A(new_n331), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n212), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT74), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n364), .B(new_n366), .C1(new_n367), .C2(KEYINPUT9), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(KEYINPUT9), .ZN(new_n369));
  XOR2_X1   g0169(.A(new_n368), .B(new_n369), .Z(new_n370));
  INV_X1    g0170(.A(KEYINPUT10), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n307), .A2(G222), .A3(new_n271), .ZN(new_n372));
  INV_X1    g0172(.A(G77), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n372), .B1(new_n373), .B2(new_n307), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n307), .A2(G1698), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT70), .ZN(new_n376));
  XNOR2_X1  g0176(.A(new_n375), .B(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n374), .B1(new_n377), .B2(G223), .ZN(new_n378));
  INV_X1    g0178(.A(new_n282), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n329), .A2(G274), .ZN(new_n381));
  XNOR2_X1  g0181(.A(KEYINPUT68), .B(G41), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n263), .B(new_n381), .C1(new_n382), .C2(G45), .ZN(new_n383));
  AOI21_X1  g0183(.A(G1), .B1(new_n253), .B2(new_n259), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n265), .B2(new_n268), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n383), .B1(new_n386), .B2(new_n213), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n380), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G200), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(G190), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n370), .A2(new_n371), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n391), .B1(new_n344), .B2(new_n388), .ZN(new_n393));
  XNOR2_X1  g0193(.A(new_n368), .B(new_n369), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT10), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT76), .ZN(new_n397));
  INV_X1    g0197(.A(G68), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(G20), .ZN(new_n399));
  OAI221_X1 g0199(.A(new_n399), .B1(new_n361), .B2(new_n373), .C1(new_n212), .C2(new_n360), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n326), .ZN(new_n401));
  XNOR2_X1  g0201(.A(new_n401), .B(KEYINPUT11), .ZN(new_n402));
  INV_X1    g0202(.A(G13), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n399), .A2(G1), .A3(new_n403), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n404), .B(KEYINPUT12), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n326), .B1(new_n329), .B2(G20), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n405), .B1(G68), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n307), .A2(G226), .A3(new_n271), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G97), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT75), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(KEYINPUT75), .A2(G33), .A3(G97), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n274), .A2(new_n276), .A3(G232), .A4(G1698), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n410), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n282), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n385), .A2(G238), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n418), .A2(new_n383), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT13), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n417), .A2(new_n282), .B1(G238), .B2(new_n385), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT13), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(new_n423), .A3(new_n383), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n421), .A2(G190), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n409), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n344), .B1(new_n421), .B2(new_n424), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n397), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n427), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n429), .A2(KEYINPUT76), .A3(new_n425), .A4(new_n409), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT78), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n408), .B(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT14), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n421), .A2(new_n424), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n434), .B1(new_n435), .B2(G169), .ZN(new_n436));
  INV_X1    g0236(.A(G169), .ZN(new_n437));
  AOI211_X1 g0237(.A(KEYINPUT14), .B(new_n437), .C1(new_n421), .C2(new_n424), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT77), .B1(new_n435), .B2(new_n350), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT77), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n421), .A2(new_n441), .A3(G179), .A4(new_n424), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n433), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n431), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n388), .A2(new_n350), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n364), .A2(new_n366), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n446), .B(new_n447), .C1(G169), .C2(new_n388), .ZN(new_n448));
  INV_X1    g0248(.A(G244), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n383), .B1(new_n386), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n377), .A2(G238), .ZN(new_n451));
  XNOR2_X1  g0251(.A(KEYINPUT72), .B(G107), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n274), .A2(new_n276), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n307), .A2(G232), .A3(new_n271), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n451), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n450), .B1(new_n457), .B2(new_n282), .ZN(new_n458));
  OR2_X1    g0258(.A1(new_n458), .A2(G169), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n331), .A2(G77), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G20), .A2(G77), .ZN(new_n461));
  XOR2_X1   g0261(.A(KEYINPUT15), .B(G87), .Z(new_n462));
  XNOR2_X1  g0262(.A(new_n462), .B(KEYINPUT73), .ZN(new_n463));
  OAI221_X1 g0263(.A(new_n461), .B1(new_n360), .B2(new_n362), .C1(new_n463), .C2(new_n361), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n460), .B1(new_n464), .B2(new_n326), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n406), .A2(G77), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n458), .A2(new_n350), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n459), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n396), .A2(new_n445), .A3(new_n448), .A4(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT79), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT7), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n307), .B2(G20), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n275), .A2(G33), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n475));
  OAI211_X1 g0275(.A(KEYINPUT7), .B(new_n230), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n398), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G58), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(new_n398), .ZN(new_n479));
  OAI21_X1  g0279(.A(G20), .B1(new_n479), .B2(new_n232), .ZN(new_n480));
  INV_X1    g0280(.A(G159), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n480), .B1(new_n481), .B2(new_n360), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n471), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT16), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT16), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n471), .B(new_n485), .C1(new_n477), .C2(new_n482), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(new_n326), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n362), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(new_n331), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n489), .B1(new_n357), .B2(new_n488), .ZN(new_n490));
  INV_X1    g0290(.A(new_n384), .ZN(new_n491));
  OAI211_X1 g0291(.A(G232), .B(new_n491), .C1(new_n289), .C2(new_n290), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n383), .ZN(new_n493));
  OR2_X1    g0293(.A1(G223), .A2(G1698), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n213), .A2(G1698), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n274), .A2(new_n494), .A3(new_n276), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G87), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n379), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n344), .B1(new_n493), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n496), .A2(new_n497), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n282), .ZN(new_n501));
  INV_X1    g0301(.A(G190), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n501), .A2(new_n502), .A3(new_n492), .A4(new_n383), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n499), .A2(KEYINPUT80), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT80), .B1(new_n499), .B2(new_n503), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n487), .B(new_n490), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT17), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n499), .A2(new_n503), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT80), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n499), .A2(KEYINPUT80), .A3(new_n503), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n513), .A2(KEYINPUT17), .A3(new_n490), .A4(new_n487), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n487), .A2(new_n490), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n501), .A2(new_n350), .A3(new_n492), .A4(new_n383), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n493), .A2(new_n498), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(G169), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT18), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n516), .A2(new_n520), .A3(KEYINPUT18), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n458), .A2(new_n344), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n465), .A2(new_n466), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n458), .A2(G190), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n515), .B(new_n525), .C1(new_n526), .C2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n470), .A2(new_n530), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n262), .A2(G257), .A3(new_n269), .ZN(new_n532));
  OAI21_X1  g0332(.A(KEYINPUT83), .B1(new_n296), .B2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n274), .A2(new_n276), .A3(G244), .A4(new_n271), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT4), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(KEYINPUT81), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n307), .A2(G244), .A3(new_n271), .A4(new_n536), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n307), .A2(G250), .A3(G1698), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n535), .A2(KEYINPUT81), .B1(G33), .B2(G283), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n282), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT83), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n262), .A2(G257), .A3(new_n269), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n301), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n533), .A2(new_n350), .A3(new_n544), .A4(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n544), .A2(new_n301), .A3(new_n546), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n437), .ZN(new_n550));
  INV_X1    g0350(.A(new_n332), .ZN(new_n551));
  INV_X1    g0351(.A(G97), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n331), .A2(G97), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n452), .B1(new_n473), .B2(new_n476), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n360), .A2(new_n373), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT6), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n552), .A2(new_n246), .ZN(new_n560));
  NOR2_X1   g0360(.A1(G97), .A2(G107), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n246), .A2(KEYINPUT6), .A3(G97), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n230), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NOR3_X1   g0364(.A1(new_n557), .A2(new_n558), .A3(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n554), .B(new_n556), .C1(new_n565), .C2(new_n328), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n548), .A2(new_n550), .A3(new_n566), .ZN(new_n567));
  AND4_X1   g0367(.A1(G190), .A2(new_n544), .A3(new_n301), .A4(new_n546), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n533), .A2(new_n544), .A3(new_n547), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n568), .B1(new_n569), .B2(G200), .ZN(new_n570));
  INV_X1    g0370(.A(new_n566), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT19), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n230), .B1(new_n415), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(G87), .A2(G97), .ZN(new_n575));
  AOI21_X1  g0375(.A(KEYINPUT85), .B1(new_n452), .B2(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(KEYINPUT85), .B(new_n575), .C1(new_n311), .C2(new_n312), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n574), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n307), .A2(new_n230), .A3(G68), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n573), .B1(new_n361), .B2(new_n552), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n326), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n463), .A2(new_n365), .ZN(new_n584));
  OR2_X1    g0384(.A1(new_n463), .A2(new_n551), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT86), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(G250), .B1(new_n329), .B2(G45), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n259), .A2(G1), .A3(G274), .ZN(new_n590));
  AOI211_X1 g0390(.A(new_n589), .B(new_n590), .C1(new_n265), .C2(new_n268), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n274), .A2(new_n276), .A3(G238), .A4(new_n271), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT84), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT84), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n307), .A2(new_n594), .A3(G238), .A4(new_n271), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n307), .A2(G244), .A3(G1698), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n593), .A2(new_n595), .A3(new_n318), .A4(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n591), .B1(new_n597), .B2(new_n282), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G179), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n437), .B2(new_n598), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n583), .A2(KEYINPUT86), .A3(new_n584), .A4(new_n585), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n588), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n598), .A2(G190), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n332), .A2(G87), .ZN(new_n604));
  AND4_X1   g0404(.A1(new_n603), .A2(new_n583), .A3(new_n584), .A4(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n598), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G200), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  AND4_X1   g0408(.A1(new_n567), .A2(new_n572), .A3(new_n602), .A4(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT87), .ZN(new_n610));
  NAND2_X1  g0410(.A1(G264), .A2(G1698), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n307), .B(new_n611), .C1(new_n277), .C2(G1698), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n612), .B(new_n282), .C1(G303), .C2(new_n307), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n262), .A2(G270), .A3(new_n269), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n301), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n332), .A2(G116), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n329), .A2(new_n214), .A3(G13), .A4(G20), .ZN(new_n617));
  NAND2_X1  g0417(.A1(G33), .A2(G283), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n618), .B(new_n230), .C1(G33), .C2(new_n552), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n214), .A2(G20), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n326), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT20), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n621), .A2(new_n622), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n616), .B(new_n617), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n615), .A2(new_n626), .A3(G169), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT21), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n610), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n621), .A2(new_n622), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n630), .A2(new_n623), .B1(G116), .B2(new_n332), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n437), .B1(new_n631), .B2(new_n617), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n632), .A2(KEYINPUT87), .A3(KEYINPUT21), .A4(new_n615), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n627), .A2(new_n628), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n301), .A2(new_n613), .A3(new_n614), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n635), .A2(G179), .A3(new_n626), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n629), .A2(new_n633), .A3(new_n634), .A4(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n626), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n615), .A2(new_n502), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n639), .B1(G200), .B2(new_n615), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n637), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  AND4_X1   g0441(.A1(new_n354), .A2(new_n531), .A3(new_n609), .A4(new_n641), .ZN(G372));
  NAND2_X1  g0442(.A1(new_n508), .A2(new_n514), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n431), .A2(new_n469), .ZN(new_n644));
  INV_X1    g0444(.A(new_n433), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n440), .A2(new_n442), .ZN(new_n646));
  INV_X1    g0446(.A(new_n424), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n423), .B1(new_n422), .B2(new_n383), .ZN(new_n648));
  OAI21_X1  g0448(.A(G169), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT14), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n435), .A2(new_n434), .A3(G169), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n645), .B1(new_n646), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n643), .B1(new_n644), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(KEYINPUT18), .B1(new_n516), .B2(new_n520), .ZN(new_n655));
  AOI211_X1 g0455(.A(new_n522), .B(new_n519), .C1(new_n487), .C2(new_n490), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n396), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n658), .A2(new_n448), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n600), .A2(new_n586), .ZN(new_n660));
  AOI21_X1  g0460(.A(KEYINPUT7), .B1(new_n454), .B2(new_n230), .ZN(new_n661));
  AOI211_X1 g0461(.A(new_n472), .B(G20), .C1(new_n274), .C2(new_n276), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n453), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n558), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n562), .A2(new_n563), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(G20), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n663), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n553), .B1(new_n667), .B2(new_n326), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n668), .A2(new_n556), .B1(new_n437), .B2(new_n549), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n570), .A2(new_n571), .B1(new_n669), .B2(new_n548), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n605), .A2(new_n607), .B1(new_n600), .B2(new_n586), .ZN(new_n671));
  AOI21_X1  g0471(.A(KEYINPUT90), .B1(new_n303), .B2(new_n336), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n345), .A2(new_n346), .A3(new_n338), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n670), .B(new_n671), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n637), .B1(new_n346), .B2(new_n353), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n660), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n567), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n602), .A2(new_n677), .A3(new_n608), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT26), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n669), .A2(KEYINPUT91), .A3(new_n548), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT91), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n567), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n671), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n679), .B1(KEYINPUT26), .B2(new_n683), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n676), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n531), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n659), .A2(new_n686), .ZN(G369));
  NAND3_X1  g0487(.A1(new_n329), .A2(new_n230), .A3(G13), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G213), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G343), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n641), .B1(new_n638), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n637), .A2(new_n626), .A3(new_n693), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n353), .A2(new_n346), .ZN(new_n699));
  OR3_X1    g0499(.A1(new_n699), .A2(KEYINPUT92), .A3(new_n694), .ZN(new_n700));
  OAI21_X1  g0500(.A(KEYINPUT92), .B1(new_n699), .B2(new_n694), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n346), .A2(new_n693), .ZN(new_n702));
  AOI22_X1  g0502(.A1(new_n700), .A2(new_n701), .B1(new_n354), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n699), .A2(new_n693), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n637), .A2(new_n694), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n707), .B1(new_n703), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n705), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT93), .ZN(G399));
  INV_X1    g0512(.A(new_n207), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(new_n382), .ZN(new_n714));
  OR3_X1    g0514(.A1(new_n576), .A2(new_n578), .A3(G116), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n714), .A2(new_n329), .A3(new_n715), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n716), .A2(KEYINPUT94), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n714), .A2(new_n235), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(KEYINPUT94), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  INV_X1    g0521(.A(G330), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT95), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT30), .ZN(new_n724));
  AOI211_X1 g0524(.A(new_n350), .B(new_n591), .C1(new_n597), .C2(new_n282), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n725), .A2(new_n635), .A3(new_n341), .A4(new_n342), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n296), .A2(new_n532), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n727), .B(new_n544), .C1(new_n723), .C2(KEYINPUT30), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n724), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n635), .A2(G179), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n730), .A2(new_n569), .A3(new_n343), .A4(new_n606), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n615), .A2(new_n285), .A3(new_n286), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n723), .A2(KEYINPUT30), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n549), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n724), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n732), .A2(new_n734), .A3(new_n725), .A4(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n729), .A2(new_n731), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n693), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(KEYINPUT31), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT31), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n737), .A2(new_n740), .A3(new_n693), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n609), .A2(new_n354), .A3(new_n641), .A4(new_n694), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n722), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n685), .A2(new_n694), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT29), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n683), .A2(KEYINPUT26), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT26), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n602), .A2(new_n677), .A3(new_n608), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g0551(.A(KEYINPUT29), .B(new_n694), .C1(new_n676), .C2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n744), .B1(new_n747), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n721), .B1(new_n753), .B2(G1), .ZN(G364));
  NOR2_X1   g0554(.A1(G13), .A2(G33), .ZN(new_n755));
  XOR2_X1   g0555(.A(new_n755), .B(KEYINPUT97), .Z(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n695), .A2(new_n696), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n344), .A2(G179), .ZN(new_n759));
  NAND2_X1  g0559(.A1(G20), .A2(G190), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n230), .A2(G190), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n759), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n307), .B1(new_n762), .B2(new_n223), .C1(new_n246), .C2(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT100), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G179), .A2(G200), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n230), .B1(new_n767), .B2(G190), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n552), .ZN(new_n769));
  NOR4_X1   g0569(.A1(new_n230), .A2(new_n350), .A3(new_n344), .A4(G190), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n760), .A2(new_n350), .A3(new_n344), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n771), .A2(new_n398), .B1(new_n773), .B2(new_n212), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n766), .A2(new_n769), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n350), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n763), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G77), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n760), .A2(new_n350), .A3(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G58), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n763), .A2(new_n767), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n481), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT99), .B(KEYINPUT32), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n775), .A2(new_n779), .A3(new_n781), .A4(new_n785), .ZN(new_n786));
  XOR2_X1   g0586(.A(KEYINPUT33), .B(G317), .Z(new_n787));
  INV_X1    g0587(.A(new_n780), .ZN(new_n788));
  INV_X1    g0588(.A(G322), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n771), .A2(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT102), .ZN(new_n791));
  INV_X1    g0591(.A(new_n782), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n791), .B1(G329), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G303), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n454), .B1(new_n762), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT101), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n795), .A2(new_n796), .B1(G326), .B2(new_n772), .ZN(new_n798));
  INV_X1    g0598(.A(new_n764), .ZN(new_n799));
  INV_X1    g0599(.A(new_n768), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G283), .A2(new_n799), .B1(new_n800), .B2(G294), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n793), .A2(new_n797), .A3(new_n798), .A4(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G311), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n777), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n786), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n229), .B1(G20), .B2(new_n437), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT98), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n713), .A2(new_n307), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT96), .Z(new_n811));
  NAND2_X1  g0611(.A1(new_n251), .A2(G45), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n811), .B(new_n812), .C1(G45), .C2(new_n234), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n207), .A2(G355), .A3(new_n307), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n813), .B(new_n814), .C1(G116), .C2(new_n207), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n808), .A2(new_n757), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n403), .A2(G20), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n329), .B1(new_n818), .B2(G45), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n714), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n758), .A2(new_n809), .A3(new_n817), .A4(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n821), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n698), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n697), .A2(G330), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(G396));
  OR2_X1    g0626(.A1(new_n469), .A2(new_n693), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n529), .A2(new_n526), .B1(new_n527), .B2(new_n694), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n469), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n745), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n469), .A2(new_n693), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n469), .B2(new_n828), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n833), .B(new_n694), .C1(new_n676), .C2(new_n684), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(new_n744), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n823), .ZN(new_n837));
  INV_X1    g0637(.A(new_n756), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n830), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n808), .A2(new_n838), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n373), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G87), .A2(new_n799), .B1(new_n792), .B2(G311), .ZN(new_n842));
  INV_X1    g0642(.A(G294), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n843), .B2(new_n788), .ZN(new_n844));
  INV_X1    g0644(.A(new_n762), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n769), .B(new_n844), .C1(G107), .C2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n773), .A2(new_n794), .ZN(new_n847));
  INV_X1    g0647(.A(G283), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n771), .A2(new_n848), .B1(new_n214), .B2(new_n777), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n307), .B(new_n847), .C1(new_n849), .C2(KEYINPUT103), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n846), .B(new_n850), .C1(KEYINPUT103), .C2(new_n849), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n764), .A2(new_n398), .B1(new_n762), .B2(new_n212), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n454), .B(new_n852), .C1(G58), .C2(new_n800), .ZN(new_n853));
  INV_X1    g0653(.A(G132), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n853), .B1(new_n854), .B2(new_n782), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT105), .ZN(new_n856));
  XNOR2_X1  g0656(.A(KEYINPUT104), .B(G143), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n778), .A2(G159), .B1(new_n780), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(G137), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n858), .B1(new_n859), .B2(new_n773), .C1(new_n359), .C2(new_n771), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT34), .Z(new_n861));
  OAI21_X1  g0661(.A(new_n851), .B1(new_n856), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n808), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n839), .A2(new_n821), .A3(new_n841), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n837), .A2(new_n864), .ZN(G384));
  INV_X1    g0665(.A(new_n691), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n516), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n515), .B2(new_n525), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n521), .A2(new_n867), .A3(new_n506), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n521), .A2(new_n867), .A3(KEYINPUT37), .A4(new_n506), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT38), .B1(new_n868), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n867), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n657), .B2(new_n643), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT38), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(new_n871), .A4(new_n872), .ZN(new_n878));
  NOR2_X1   g0678(.A1(KEYINPUT108), .A2(KEYINPUT38), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n874), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n876), .A2(new_n871), .A3(new_n872), .A4(new_n879), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n742), .A2(new_n743), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n428), .A2(new_n430), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n433), .A2(new_n694), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n653), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n886), .B1(new_n431), .B2(new_n444), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n830), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n883), .A2(KEYINPUT40), .A3(new_n884), .A4(new_n890), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n890), .A2(new_n884), .A3(new_n874), .A4(new_n878), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT40), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n893), .A2(KEYINPUT109), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(KEYINPUT109), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n892), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n891), .A2(new_n897), .A3(G330), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n531), .A2(new_n744), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n531), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n891), .A2(new_n897), .A3(new_n884), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n747), .A2(new_n531), .A3(new_n752), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n659), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n903), .B(new_n905), .Z(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n881), .A2(new_n907), .A3(new_n882), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n874), .A2(KEYINPUT39), .A3(new_n878), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT107), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT107), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n874), .A2(new_n911), .A3(new_n878), .A4(KEYINPUT39), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n908), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n653), .A2(new_n693), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n913), .A2(new_n914), .B1(new_n657), .B2(new_n691), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n834), .A2(new_n827), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n889), .A2(new_n888), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n916), .A2(new_n874), .A3(new_n878), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n906), .B(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n329), .B2(new_n818), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n214), .B1(new_n665), .B2(KEYINPUT35), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n922), .B(new_n231), .C1(KEYINPUT35), .C2(new_n665), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT36), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n234), .A2(new_n373), .A3(new_n479), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT106), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(G50), .B2(new_n398), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(G1), .A3(new_n403), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n921), .A2(new_n924), .A3(new_n928), .ZN(G367));
  NOR2_X1   g0729(.A1(new_n703), .A2(new_n708), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n566), .A2(new_n693), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n670), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(KEYINPUT42), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n567), .B1(new_n932), .B2(new_n699), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n694), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT42), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n930), .A2(new_n938), .A3(new_n933), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n935), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n583), .A2(new_n584), .A3(new_n604), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n693), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n671), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n660), .A2(new_n942), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n940), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n947), .B1(new_n940), .B2(new_n948), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n932), .B1(new_n567), .B2(new_n694), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n705), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n949), .A2(new_n950), .A3(new_n954), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n935), .A2(new_n939), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT43), .ZN(new_n957));
  INV_X1    g0757(.A(new_n945), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n956), .A2(new_n957), .A3(new_n958), .A4(new_n937), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n940), .A2(new_n947), .A3(new_n948), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n953), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n955), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n819), .B(KEYINPUT110), .Z(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n753), .ZN(new_n965));
  OAI21_X1  g0765(.A(KEYINPUT44), .B1(new_n710), .B2(new_n951), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT44), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n709), .A2(new_n967), .A3(new_n952), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n707), .B(new_n951), .C1(new_n703), .C2(new_n708), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT45), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n966), .B(new_n968), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n698), .A2(new_n708), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(new_n703), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n965), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n714), .B(KEYINPUT41), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n964), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n962), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n782), .A2(new_n859), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n771), .A2(new_n481), .B1(new_n212), .B2(new_n777), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n981), .B(new_n982), .C1(new_n772), .C2(new_n857), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n764), .A2(new_n373), .B1(new_n762), .B2(new_n478), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n454), .B(new_n984), .C1(G150), .C2(new_n780), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n983), .B(new_n985), .C1(new_n398), .C2(new_n768), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT111), .Z(new_n987));
  NAND2_X1  g0787(.A1(new_n778), .A2(G283), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n762), .A2(new_n214), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT46), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n454), .B1(new_n794), .B2(new_n788), .C1(new_n771), .C2(new_n843), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n453), .B2(new_n800), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n792), .A2(G317), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(new_n552), .C2(new_n764), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n990), .B(new_n994), .C1(G311), .C2(new_n772), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n987), .B1(new_n988), .B2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT47), .Z(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n808), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n958), .A2(new_n757), .ZN(new_n999));
  INV_X1    g0799(.A(new_n811), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n816), .B1(new_n207), .B2(new_n463), .C1(new_n1000), .C2(new_n243), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n998), .A2(new_n821), .A3(new_n999), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n980), .A2(new_n1002), .ZN(G387));
  NAND2_X1  g0803(.A1(new_n975), .A2(new_n963), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n788), .A2(new_n212), .B1(new_n764), .B2(new_n552), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n463), .A2(new_n768), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(G68), .C2(new_n778), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n845), .A2(G77), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n454), .B1(new_n792), .B2(G150), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n770), .A2(new_n488), .B1(G159), .B2(new_n772), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G294), .A2(new_n845), .B1(new_n800), .B2(G283), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n778), .A2(G303), .B1(new_n780), .B2(G317), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n803), .B2(new_n771), .C1(new_n789), .C2(new_n773), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT48), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT112), .Z(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n1015), .B2(new_n1014), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(KEYINPUT49), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n799), .A2(G116), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n792), .A2(G326), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1019), .A2(new_n454), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1018), .A2(KEYINPUT49), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1011), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n808), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n488), .A2(new_n212), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT50), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n398), .A2(new_n373), .ZN(new_n1028));
  NOR4_X1   g0828(.A1(new_n1027), .A2(new_n715), .A3(G45), .A4(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n811), .B1(new_n259), .B2(new_n240), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n715), .A2(new_n207), .A3(new_n307), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n207), .A2(G107), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n816), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n703), .A2(new_n757), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1025), .A2(new_n821), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n753), .A2(new_n975), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n714), .B1(new_n753), .B2(new_n975), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1004), .B(new_n1036), .C1(new_n1038), .C2(new_n1039), .ZN(G393));
  OR2_X1    g0840(.A1(new_n971), .A2(new_n972), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1041), .A2(new_n705), .A3(new_n966), .A4(new_n968), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n973), .A2(new_n704), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n1037), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1038), .A2(new_n973), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1045), .A2(new_n714), .A3(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1042), .A2(new_n1043), .A3(new_n963), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n816), .B1(new_n552), .B2(new_n207), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n811), .B2(new_n248), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G150), .A2(new_n772), .B1(new_n780), .B2(G159), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT51), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n454), .B1(new_n792), .B2(new_n857), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n373), .B2(new_n768), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n362), .A2(new_n777), .B1(new_n764), .B2(new_n223), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1052), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n212), .B2(new_n771), .C1(new_n398), .C2(new_n762), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G317), .A2(new_n772), .B1(new_n780), .B2(G311), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT52), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n307), .B(new_n1059), .C1(G303), .C2(new_n770), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n800), .A2(G116), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n792), .A2(G322), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n799), .A2(G107), .B1(new_n845), .B2(G283), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n777), .A2(new_n843), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1057), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1050), .B1(new_n1066), .B2(new_n808), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n757), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n821), .B(new_n1067), .C1(new_n951), .C2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1048), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1047), .A2(new_n1071), .ZN(G390));
  OAI211_X1 g0872(.A(new_n694), .B(new_n829), .C1(new_n676), .C2(new_n751), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n827), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n917), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n914), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1075), .A2(new_n1076), .A3(new_n883), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1077), .B1(new_n913), .B2(new_n1078), .ZN(new_n1079));
  AND4_X1   g0879(.A1(G330), .A2(new_n884), .A3(new_n917), .A4(new_n833), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n744), .A2(new_n833), .A3(new_n917), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1077), .B(new_n1082), .C1(new_n913), .C2(new_n1078), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n963), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n823), .B1(new_n362), .B2(new_n840), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT114), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n845), .A2(G150), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n1088));
  NOR2_X1   g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n454), .B1(new_n792), .B2(G125), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n772), .A2(G128), .ZN(new_n1091));
  XOR2_X1   g0891(.A(KEYINPUT54), .B(G143), .Z(new_n1092));
  NAND2_X1  g0892(.A1(new_n778), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1090), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1089), .B(new_n1094), .C1(G50), .C2(new_n799), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1087), .A2(new_n1088), .B1(new_n800), .B2(G159), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n1097), .B1(new_n854), .B2(new_n788), .C1(new_n859), .C2(new_n771), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n771), .A2(new_n452), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n454), .B1(new_n788), .B2(new_n214), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n764), .A2(new_n398), .B1(new_n762), .B2(new_n223), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n777), .A2(new_n552), .B1(new_n768), .B2(new_n373), .ZN(new_n1102));
  NOR4_X1   g0902(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1103), .B1(new_n848), .B2(new_n773), .C1(new_n843), .C2(new_n782), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1098), .A2(new_n1104), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1086), .B1(new_n807), .B2(new_n1105), .C1(new_n913), .C2(new_n756), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n917), .B1(new_n744), .B2(new_n833), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n916), .B1(new_n1080), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT113), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OR3_X1    g0910(.A1(new_n1080), .A2(new_n1107), .A3(new_n1074), .ZN(new_n1111));
  OAI211_X1 g0911(.A(KEYINPUT113), .B(new_n916), .C1(new_n1080), .C2(new_n1107), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n904), .A2(new_n659), .A3(new_n899), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1081), .A2(new_n1083), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n714), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1081), .A2(new_n1083), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1084), .B(new_n1106), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT116), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1123), .A2(new_n714), .A3(new_n1115), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1124), .A2(KEYINPUT116), .A3(new_n1084), .A4(new_n1106), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1120), .A2(new_n1125), .ZN(G378));
  XOR2_X1   g0926(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n396), .A2(new_n448), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1128), .B1(new_n396), .B2(new_n448), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n447), .A2(new_n866), .ZN(new_n1131));
  OR3_X1    g0931(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1131), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n898), .A2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n891), .A2(new_n897), .A3(new_n1134), .A4(G330), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n919), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1136), .A2(new_n1137), .A3(new_n918), .A4(new_n915), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n768), .A2(new_n398), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n773), .A2(new_n214), .B1(new_n764), .B2(new_n478), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n1142), .B(new_n1143), .C1(G97), .C2(new_n770), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1008), .B1(new_n848), .B2(new_n782), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n254), .A2(new_n256), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n454), .B(new_n1146), .C1(new_n788), .C2(new_n246), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1144), .B(new_n1148), .C1(new_n463), .C2(new_n777), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT58), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n273), .A2(new_n253), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT117), .ZN(new_n1152));
  AOI211_X1 g0952(.A(G50), .B(new_n1152), .C1(new_n454), .C2(new_n1146), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT118), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(G137), .A2(new_n778), .B1(new_n845), .B2(new_n1092), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n800), .A2(G150), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n772), .A2(G125), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n770), .A2(G132), .B1(G128), .B2(new_n780), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1159), .B(KEYINPUT59), .Z(new_n1160));
  NAND2_X1  g0960(.A1(new_n799), .A2(G159), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n792), .A2(G124), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1160), .A2(new_n1152), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1150), .A2(new_n1154), .A3(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT119), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1165), .A2(new_n808), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1135), .A2(new_n756), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(new_n212), .C2(new_n840), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1141), .A2(new_n963), .B1(new_n821), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1115), .A2(new_n1114), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1170), .A2(KEYINPUT57), .A3(new_n1140), .A4(new_n1139), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n714), .ZN(new_n1172));
  AOI21_X1  g0972(.A(KEYINPUT57), .B1(new_n1141), .B2(new_n1170), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1169), .B1(new_n1172), .B2(new_n1173), .ZN(G375));
  AOI21_X1  g0974(.A(new_n1006), .B1(new_n453), .B2(new_n778), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n848), .B2(new_n788), .C1(new_n843), .C2(new_n773), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n762), .A2(new_n552), .B1(new_n782), .B2(new_n794), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1177), .A2(KEYINPUT120), .B1(G116), .B2(new_n770), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(KEYINPUT120), .B2(new_n1177), .C1(new_n373), .C2(new_n764), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1176), .A2(new_n307), .A3(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G159), .A2(new_n845), .B1(new_n792), .B2(G128), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1181), .A2(KEYINPUT122), .B1(new_n770), .B2(new_n1092), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n359), .B2(new_n777), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n772), .A2(G132), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT121), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n454), .B1(G137), .B2(new_n780), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1186), .B1(new_n212), .B2(new_n768), .C1(new_n478), .C2(new_n764), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1181), .A2(KEYINPUT122), .ZN(new_n1188));
  NOR4_X1   g0988(.A1(new_n1183), .A2(new_n1185), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n808), .B1(new_n1180), .B2(new_n1189), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n821), .B(new_n1190), .C1(new_n917), .C2(new_n756), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n398), .B2(new_n840), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n1113), .B2(new_n963), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1122), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n977), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1193), .B1(new_n1194), .B2(new_n1195), .ZN(G381));
  NAND2_X1  g0996(.A1(new_n1168), .A2(new_n821), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1197), .B1(new_n1198), .B2(new_n964), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1171), .A2(new_n714), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT57), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1170), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1201), .B1(new_n1202), .B2(new_n1198), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1199), .B1(new_n1200), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1118), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1046), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n1044), .B2(new_n1037), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1070), .B1(new_n1208), .B2(new_n714), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1002), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n962), .B2(new_n979), .ZN(new_n1211));
  INV_X1    g1011(.A(G384), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(G393), .A2(G396), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1209), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  OR3_X1    g1014(.A1(new_n1206), .A2(G381), .A3(new_n1214), .ZN(G407));
  OAI211_X1 g1015(.A(G407), .B(G213), .C1(G343), .C2(new_n1206), .ZN(G409));
  INV_X1    g1016(.A(KEYINPUT126), .ZN(new_n1217));
  OAI21_X1  g1017(.A(KEYINPUT123), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n714), .B(new_n1122), .C1(new_n1218), .C2(KEYINPUT60), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1218), .A2(KEYINPUT60), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1193), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n1212), .ZN(new_n1222));
  OAI211_X1 g1022(.A(G384), .B(new_n1193), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1223));
  INV_X1    g1023(.A(G213), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1224), .A2(G343), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(G2897), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1222), .A2(new_n1223), .A3(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1226), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1141), .A2(new_n977), .A3(new_n1170), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1118), .B1(new_n1169), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1204), .B2(G378), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1229), .B1(new_n1232), .B2(new_n1225), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1203), .A2(new_n714), .A3(new_n1171), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(G378), .A2(new_n1169), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1169), .A2(new_n1230), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n1205), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n1234), .B(new_n1225), .C1(new_n1236), .C2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT62), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1233), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT61), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1120), .A2(new_n1125), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1238), .B1(new_n1243), .B2(G375), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1234), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1225), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1242), .B1(new_n1247), .B2(KEYINPUT62), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1217), .B1(new_n1241), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1247), .A2(KEYINPUT62), .B1(new_n1250), .B2(new_n1229), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT61), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1251), .A2(new_n1252), .A3(KEYINPUT126), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT125), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(G390), .B2(new_n1211), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(G390), .A2(new_n1211), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  XOR2_X1   g1057(.A(G393), .B(G396), .Z(new_n1258));
  NOR2_X1   g1058(.A1(G390), .A2(new_n1211), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1258), .B1(new_n1259), .B2(KEYINPUT125), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1258), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(new_n1259), .B2(KEYINPUT124), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G387), .A2(new_n1209), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT124), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(new_n1256), .A3(new_n1264), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n1257), .A2(new_n1260), .B1(new_n1262), .B2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1249), .A2(new_n1253), .A3(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(KEYINPUT61), .B1(new_n1239), .B2(KEYINPUT63), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1262), .A2(new_n1265), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(G387), .A2(new_n1209), .A3(KEYINPUT125), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1270), .A2(new_n1255), .A3(new_n1256), .A4(new_n1261), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1233), .A2(KEYINPUT63), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1268), .B(new_n1272), .C1(new_n1273), .C2(new_n1239), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1267), .A2(new_n1274), .ZN(G405));
  INV_X1    g1075(.A(new_n1236), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1204), .A2(new_n1118), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1266), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1277), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1272), .A2(new_n1236), .A3(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT127), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1278), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1281), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1234), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(KEYINPUT127), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1278), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1286), .A2(new_n1245), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1284), .A2(new_n1288), .ZN(G402));
endmodule


