//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n807,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n203));
  INV_X1    g002(.A(G134gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(KEYINPUT68), .ZN(new_n205));
  XNOR2_X1  g004(.A(G113gat), .B(G120gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n206), .B2(KEYINPUT1), .ZN(new_n207));
  INV_X1    g006(.A(G127gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n209));
  INV_X1    g008(.A(G113gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(G120gat), .ZN(new_n211));
  INV_X1    g010(.A(G120gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n212), .A2(G113gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n209), .B(new_n204), .C1(new_n211), .C2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n207), .A2(new_n208), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n208), .B1(new_n207), .B2(new_n214), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n203), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n207), .A2(new_n214), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G127gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n220), .A2(KEYINPUT69), .A3(new_n215), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT70), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT25), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g029(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n227), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT23), .B1(new_n233), .B2(KEYINPUT65), .ZN(new_n234));
  NAND2_X1  g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT23), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n236), .B(new_n237), .C1(G169gat), .C2(G176gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n234), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n224), .B1(new_n232), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n224), .B1(new_n227), .B2(new_n228), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n243), .A2(new_n234), .A3(new_n235), .A4(new_n238), .ZN(new_n244));
  OAI211_X1 g043(.A(KEYINPUT66), .B(new_n224), .C1(new_n232), .C2(new_n239), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT27), .B(G183gat), .ZN(new_n247));
  INV_X1    g046(.A(G190gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT67), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT28), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(KEYINPUT67), .A3(KEYINPUT28), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT26), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n233), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n235), .A3(new_n256), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n252), .A2(new_n226), .A3(new_n253), .A4(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n222), .A2(new_n223), .A3(new_n246), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n246), .A2(new_n258), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n218), .A2(new_n221), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT70), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G227gat), .A2(G233gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n260), .A2(new_n261), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n259), .A2(new_n262), .A3(new_n263), .A4(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT34), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n259), .A2(new_n262), .A3(new_n264), .ZN(new_n267));
  INV_X1    g066(.A(new_n263), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT32), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n267), .A2(new_n268), .B1(new_n269), .B2(KEYINPUT33), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT71), .B(G71gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(G99gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(G15gat), .B(G43gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n274), .A2(KEYINPUT72), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT33), .B1(new_n274), .B2(KEYINPUT72), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI211_X1 g077(.A(new_n269), .B(new_n278), .C1(new_n267), .C2(new_n268), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n266), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n275), .A2(new_n266), .A3(new_n279), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n202), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n270), .A2(new_n274), .ZN(new_n284));
  INV_X1    g083(.A(new_n279), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT34), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n265), .B(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n284), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(KEYINPUT36), .A3(new_n280), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G225gat), .A2(G233gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT82), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n220), .A2(new_n215), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT81), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT77), .ZN(new_n297));
  INV_X1    g096(.A(G141gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G148gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n298), .A2(G148gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n297), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n301), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n303), .A2(new_n299), .A3(KEYINPUT77), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT2), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G155gat), .B(G162gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT2), .ZN(new_n310));
  INV_X1    g109(.A(G148gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n298), .A2(KEYINPUT78), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT78), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G141gat), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n311), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n310), .B(new_n307), .C1(new_n315), .C2(new_n301), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT80), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT78), .B(G141gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n303), .B1(new_n319), .B2(new_n311), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n320), .A2(KEYINPUT80), .A3(new_n310), .A4(new_n307), .ZN(new_n321));
  AOI221_X4 g120(.A(new_n296), .B1(new_n306), .B2(new_n308), .C1(new_n318), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(new_n321), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT81), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n293), .B(new_n295), .C1(new_n322), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n323), .A2(new_n324), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n296), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n318), .A2(new_n321), .B1(new_n308), .B2(new_n306), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT81), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n294), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n293), .B1(new_n329), .B2(new_n294), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n292), .B(new_n326), .C1(new_n331), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT83), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT3), .B1(new_n322), .B2(new_n325), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT3), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n329), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n338), .A3(new_n295), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n329), .A2(new_n294), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT4), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n222), .A2(KEYINPUT4), .A3(new_n329), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n339), .A2(new_n291), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT84), .B(KEYINPUT5), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n295), .B1(new_n322), .B2(new_n325), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(new_n332), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT83), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n347), .A2(new_n348), .A3(new_n292), .A4(new_n326), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n335), .A2(new_n344), .A3(new_n345), .A4(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n341), .B1(new_n261), .B2(new_n327), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n329), .A2(KEYINPUT4), .A3(new_n294), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n339), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n345), .A2(new_n292), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  XOR2_X1   g155(.A(G1gat), .B(G29gat), .Z(new_n357));
  XNOR2_X1  g156(.A(G57gat), .B(G85gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT85), .B(KEYINPUT0), .ZN(new_n360));
  XOR2_X1   g159(.A(new_n359), .B(new_n360), .Z(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n356), .A2(KEYINPUT6), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n350), .A2(new_n361), .A3(new_n355), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT6), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n361), .B1(new_n350), .B2(new_n355), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n363), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G8gat), .B(G36gat), .ZN(new_n369));
  INV_X1    g168(.A(G64gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G92gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  XOR2_X1   g173(.A(KEYINPUT73), .B(G204gat), .Z(new_n375));
  INV_X1    g174(.A(G197gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT22), .ZN(new_n378));
  INV_X1    g177(.A(G211gat), .ZN(new_n379));
  INV_X1    g178(.A(G218gat), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT73), .B(G204gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G197gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n377), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT74), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G211gat), .B(G218gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT29), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n260), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G226gat), .A2(G233gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n394), .B1(new_n246), .B2(new_n258), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n391), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n260), .A2(new_n392), .B1(G226gat), .B2(G233gat), .ZN(new_n399));
  INV_X1    g198(.A(new_n391), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n399), .A2(new_n400), .A3(new_n396), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n374), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT76), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT30), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n395), .A2(new_n391), .A3(new_n397), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n400), .B1(new_n399), .B2(new_n396), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n408), .A2(KEYINPUT76), .A3(new_n374), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n404), .A2(new_n405), .A3(new_n409), .ZN(new_n410));
  XOR2_X1   g209(.A(new_n373), .B(KEYINPUT75), .Z(new_n411));
  OR2_X1    g210(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n408), .A2(KEYINPUT30), .A3(new_n374), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n410), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n368), .A2(new_n414), .A3(KEYINPUT86), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT86), .B1(new_n368), .B2(new_n414), .ZN(new_n416));
  XNOR2_X1  g215(.A(G78gat), .B(G106gat), .ZN(new_n417));
  XOR2_X1   g216(.A(new_n417), .B(KEYINPUT31), .Z(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n384), .A2(new_n387), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n392), .B1(new_n384), .B2(new_n387), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n337), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n327), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT87), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G228gat), .A2(G233gat), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n323), .A2(new_n337), .A3(new_n324), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n391), .B1(new_n427), .B2(KEYINPUT29), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n422), .A2(KEYINPUT87), .A3(new_n327), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n425), .A2(new_n426), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT88), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n431), .B1(new_n427), .B2(KEYINPUT29), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n338), .A2(KEYINPUT88), .A3(new_n392), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n391), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n337), .B1(new_n391), .B2(KEYINPUT29), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n435), .B1(new_n325), .B2(new_n322), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n419), .B(new_n430), .C1(new_n437), .C2(new_n426), .ZN(new_n438));
  XNOR2_X1  g237(.A(G22gat), .B(G50gat), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n426), .B1(new_n434), .B2(new_n436), .ZN(new_n440));
  INV_X1    g239(.A(new_n430), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n418), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n438), .A2(new_n439), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n439), .B1(new_n438), .B2(new_n442), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n415), .A2(new_n416), .A3(new_n446), .ZN(new_n447));
  AOI211_X1 g246(.A(new_n365), .B(new_n361), .C1(new_n350), .C2(new_n355), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT89), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n356), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n350), .A2(KEYINPUT89), .A3(new_n355), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(new_n362), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n366), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n448), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT37), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n408), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n373), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n408), .A2(new_n455), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT38), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n404), .A2(new_n409), .ZN(new_n460));
  INV_X1    g259(.A(new_n458), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n411), .A2(KEYINPUT38), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n456), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n454), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n353), .A2(new_n292), .ZN(new_n467));
  OR2_X1    g266(.A1(new_n467), .A2(KEYINPUT39), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n347), .A2(new_n326), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n467), .B(KEYINPUT39), .C1(new_n292), .C2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n470), .A3(new_n361), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT40), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n410), .A2(new_n412), .A3(new_n413), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n468), .A2(new_n470), .A3(KEYINPUT40), .A4(new_n361), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n452), .A2(new_n473), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n445), .B1(new_n466), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n290), .B1(new_n447), .B2(new_n477), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n288), .B(new_n280), .C1(new_n443), .C2(new_n444), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n454), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT35), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(new_n414), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n415), .A2(new_n416), .A3(new_n479), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n482), .B1(new_n483), .B2(new_n481), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  XOR2_X1   g284(.A(G71gat), .B(G78gat), .Z(new_n486));
  INV_X1    g285(.A(KEYINPUT9), .ZN(new_n487));
  XNOR2_X1  g286(.A(G57gat), .B(G64gat), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT94), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(G71gat), .ZN(new_n492));
  INV_X1    g291(.A(G78gat), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n487), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n494), .A2(KEYINPUT95), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n495), .A2(new_n486), .A3(new_n488), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(KEYINPUT95), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n491), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(KEYINPUT96), .A2(G85gat), .A3(G92gat), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT7), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G99gat), .A2(G106gat), .ZN(new_n503));
  INV_X1    g302(.A(G85gat), .ZN(new_n504));
  AOI22_X1  g303(.A1(KEYINPUT8), .A2(new_n503), .B1(new_n504), .B2(new_n372), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n500), .A2(new_n501), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n502), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  XOR2_X1   g306(.A(G99gat), .B(G106gat), .Z(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n499), .B(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT10), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n510), .A2(KEYINPUT10), .A3(new_n498), .A4(new_n491), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G230gat), .ZN(new_n516));
  INV_X1    g315(.A(G233gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n511), .A2(new_n519), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G120gat), .B(G148gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(G204gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT97), .ZN(new_n525));
  INV_X1    g324(.A(G176gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n527), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n520), .A2(new_n521), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G15gat), .B(G22gat), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT16), .ZN(new_n534));
  AOI21_X1  g333(.A(G1gat), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(KEYINPUT92), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(KEYINPUT93), .A2(G8gat), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n533), .B(KEYINPUT92), .C1(new_n534), .C2(G1gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(KEYINPUT93), .A2(G8gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT21), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n542), .B1(new_n543), .B2(new_n499), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(G183gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(G231gat), .A2(G233gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G127gat), .B(G155gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(new_n379), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n547), .B(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n499), .A2(new_n543), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n551), .B(new_n552), .Z(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  OR2_X1    g353(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n550), .A2(new_n554), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n558), .A2(KEYINPUT41), .ZN(new_n559));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT14), .ZN(new_n563));
  INV_X1    g362(.A(G29gat), .ZN(new_n564));
  INV_X1    g363(.A(G36gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n566), .A2(new_n567), .B1(G29gat), .B2(G36gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(G43gat), .B(G50gat), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n568), .B1(KEYINPUT15), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(KEYINPUT15), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  OR2_X1    g371(.A1(new_n572), .A2(KEYINPUT17), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT91), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(KEYINPUT17), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(new_n509), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G134gat), .B(G162gat), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n572), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n579), .A2(new_n510), .B1(KEYINPUT41), .B2(new_n558), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n576), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n578), .B1(new_n576), .B2(new_n580), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n562), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n583), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(new_n561), .A3(new_n581), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n557), .A2(new_n588), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n542), .A2(new_n572), .ZN(new_n590));
  NAND2_X1  g389(.A1(G229gat), .A2(G233gat), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT91), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n573), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n542), .A2(new_n575), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n590), .B(new_n591), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT18), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n574), .A2(new_n542), .A3(new_n575), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n598), .A2(KEYINPUT18), .A3(new_n590), .A4(new_n591), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n542), .A2(new_n572), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n590), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n591), .B(KEYINPUT13), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n597), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G113gat), .B(G141gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G169gat), .B(G197gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n609), .B(KEYINPUT12), .Z(new_n610));
  NAND2_X1  g409(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n610), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n597), .A2(new_n599), .A3(new_n603), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n589), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n485), .A2(new_n532), .A3(new_n616), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n617), .A2(KEYINPUT98), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(KEYINPUT98), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n368), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g422(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n624));
  INV_X1    g423(.A(G8gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n534), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n620), .A2(new_n474), .A3(new_n624), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT42), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n414), .B1(new_n618), .B2(new_n619), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT42), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n629), .A2(new_n630), .A3(new_n624), .A4(new_n626), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n618), .A2(new_n619), .ZN(new_n633));
  OAI211_X1 g432(.A(KEYINPUT99), .B(G8gat), .C1(new_n633), .C2(new_n414), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n635), .B1(new_n629), .B2(new_n625), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n632), .A2(new_n637), .ZN(G1325gat));
  INV_X1    g437(.A(G15gat), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n283), .A2(new_n640), .A3(new_n289), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n640), .B1(new_n283), .B2(new_n289), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n633), .A2(new_n639), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n281), .A2(new_n282), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n620), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n639), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n647), .A2(KEYINPUT100), .A3(new_n639), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n645), .B1(new_n650), .B2(new_n651), .ZN(G1326gat));
  NAND2_X1  g451(.A1(new_n620), .A2(new_n445), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT43), .B(G22gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1327gat));
  AOI21_X1  g454(.A(new_n588), .B1(new_n478), .B2(new_n484), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n557), .A2(new_n531), .A3(new_n615), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n659), .A2(new_n564), .A3(new_n621), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n660), .A2(KEYINPUT102), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(KEYINPUT102), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT45), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n361), .B1(new_n356), .B2(new_n449), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n366), .B1(new_n667), .B2(new_n451), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n668), .A2(new_n464), .A3(new_n448), .ZN(new_n669));
  INV_X1    g468(.A(new_n476), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n446), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n368), .A2(new_n414), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT86), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n368), .A2(new_n414), .A3(KEYINPUT86), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(new_n445), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n643), .B1(new_n671), .B2(new_n676), .ZN(new_n677));
  NOR4_X1   g476(.A1(new_n454), .A2(KEYINPUT35), .A3(new_n474), .A4(new_n479), .ZN(new_n678));
  INV_X1    g477(.A(new_n479), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n674), .A2(new_n675), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n678), .B1(new_n680), .B2(KEYINPUT35), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n666), .B(new_n587), .C1(new_n677), .C2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n656), .B2(new_n666), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n657), .ZN(new_n684));
  OAI21_X1  g483(.A(G29gat), .B1(new_n684), .B2(new_n368), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n661), .A2(KEYINPUT45), .A3(new_n662), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n665), .A2(new_n685), .A3(new_n686), .ZN(G1328gat));
  NAND3_X1  g486(.A1(new_n683), .A2(new_n474), .A3(new_n657), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n683), .A2(KEYINPUT104), .A3(new_n474), .A4(new_n657), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n690), .A2(G36gat), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT103), .B(KEYINPUT46), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n659), .A2(new_n565), .A3(new_n474), .A4(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n656), .A2(new_n474), .A3(new_n657), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n693), .B1(new_n696), .B2(G36gat), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n692), .A2(KEYINPUT105), .A3(new_n698), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(G1329gat));
  INV_X1    g502(.A(KEYINPUT47), .ZN(new_n704));
  INV_X1    g503(.A(new_n646), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n658), .A2(G43gat), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n684), .A2(new_n644), .ZN(new_n709));
  INV_X1    g508(.A(G43gat), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n704), .B1(new_n708), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n706), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n683), .A2(new_n643), .A3(new_n657), .ZN(new_n716));
  OAI21_X1  g515(.A(G43gat), .B1(new_n716), .B2(KEYINPUT107), .ZN(new_n717));
  OAI211_X1 g516(.A(KEYINPUT47), .B(new_n713), .C1(new_n715), .C2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n712), .A2(new_n718), .ZN(G1330gat));
  OAI21_X1  g518(.A(G50gat), .B1(new_n684), .B2(new_n446), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n721), .A2(KEYINPUT48), .ZN(new_n722));
  OR3_X1    g521(.A1(new_n658), .A2(G50gat), .A3(new_n446), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n720), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(KEYINPUT48), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1331gat));
  NOR2_X1   g525(.A1(new_n677), .A2(new_n681), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n532), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n557), .A2(new_n588), .A3(new_n615), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(new_n368), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(G57gat), .Z(G1332gat));
  AOI211_X1 g532(.A(new_n414), .B(new_n731), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n734));
  NOR2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1333gat));
  OAI21_X1  g535(.A(new_n492), .B1(new_n731), .B2(new_n705), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n728), .A2(G71gat), .A3(new_n730), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n644), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g539(.A1(new_n731), .A2(new_n446), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(new_n493), .ZN(G1335gat));
  NOR2_X1   g541(.A1(new_n557), .A2(new_n614), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n683), .A2(new_n531), .A3(new_n743), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n744), .A2(new_n504), .A3(new_n368), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n587), .B(new_n743), .C1(new_n677), .C2(new_n681), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n748), .A2(new_n621), .A3(new_n531), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n745), .B1(new_n504), .B2(new_n749), .ZN(G1336gat));
  OR2_X1    g549(.A1(new_n744), .A2(new_n414), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G92gat), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n414), .A2(new_n532), .A3(G92gat), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT52), .B1(new_n748), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n748), .A2(new_n757), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n753), .A2(new_n756), .ZN(new_n759));
  AOI22_X1  g558(.A1(G92gat), .A2(new_n751), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n755), .B1(new_n760), .B2(new_n761), .ZN(G1337gat));
  XOR2_X1   g561(.A(KEYINPUT110), .B(G99gat), .Z(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(new_n744), .B2(new_n644), .ZN(new_n764));
  INV_X1    g563(.A(new_n763), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n748), .A2(new_n531), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n764), .B1(new_n766), .B2(new_n705), .ZN(G1338gat));
  OAI21_X1  g566(.A(G106gat), .B1(new_n744), .B2(new_n446), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n446), .A2(G106gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n748), .A2(new_n531), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g571(.A(new_n557), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n513), .A2(new_n514), .A3(new_n518), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n520), .A2(KEYINPUT54), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n518), .B1(new_n513), .B2(new_n514), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n529), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n775), .A2(KEYINPUT55), .A3(new_n778), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(new_n530), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT111), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n781), .A2(new_n785), .A3(new_n530), .A4(new_n782), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n784), .A2(new_n614), .A3(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n590), .A2(new_n600), .A3(new_n602), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n788), .B(KEYINPUT112), .Z(new_n789));
  AOI21_X1  g588(.A(new_n591), .B1(new_n598), .B2(new_n590), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n609), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n531), .A2(new_n791), .A3(new_n613), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n587), .B1(new_n787), .B2(new_n792), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n587), .A2(new_n613), .A3(new_n791), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(new_n784), .A3(new_n786), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n773), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n797), .B1(new_n531), .B2(new_n729), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n798), .A2(new_n679), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n368), .A2(new_n474), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n614), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n531), .ZN(new_n804));
  XOR2_X1   g603(.A(KEYINPUT113), .B(G120gat), .Z(new_n805));
  XNOR2_X1  g604(.A(new_n804), .B(new_n805), .ZN(G1341gat));
  NAND2_X1  g605(.A1(new_n801), .A2(new_n557), .ZN(new_n807));
  XOR2_X1   g606(.A(KEYINPUT68), .B(G127gat), .Z(new_n808));
  XNOR2_X1  g607(.A(new_n807), .B(new_n808), .ZN(G1342gat));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT56), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n801), .B(new_n587), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n812), .A2(G134gat), .B1(KEYINPUT114), .B2(KEYINPUT56), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n801), .A2(new_n587), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n814), .A2(new_n810), .A3(new_n811), .A4(new_n204), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n813), .B(new_n815), .C1(new_n204), .C2(new_n814), .ZN(G1343gat));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n643), .A2(new_n368), .A3(new_n474), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n615), .A2(G141gat), .ZN(new_n819));
  AND4_X1   g618(.A1(new_n445), .A2(new_n798), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n798), .A2(new_n821), .A3(new_n445), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n775), .B2(new_n778), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n824), .A2(new_n780), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n780), .ZN(new_n826));
  AND4_X1   g625(.A1(new_n530), .A2(new_n825), .A3(new_n614), .A4(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n792), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n531), .A2(new_n791), .A3(new_n613), .A4(KEYINPUT115), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n588), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n557), .B1(new_n832), .B2(new_n795), .ZN(new_n833));
  AND4_X1   g632(.A1(new_n532), .A2(new_n557), .A3(new_n588), .A4(new_n615), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n445), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT57), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n822), .A2(new_n836), .A3(new_n614), .A4(new_n818), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n820), .B1(new_n837), .B2(new_n319), .ZN(new_n838));
  AOI211_X1 g637(.A(new_n817), .B(KEYINPUT58), .C1(new_n838), .C2(KEYINPUT118), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(KEYINPUT118), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT117), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n842), .B1(new_n838), .B2(new_n817), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n839), .B1(new_n841), .B2(new_n843), .ZN(G1344gat));
  AND2_X1   g643(.A1(new_n798), .A2(new_n445), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n818), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n846), .A2(G148gat), .A3(new_n532), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT119), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n849));
  INV_X1    g648(.A(new_n783), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n794), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n557), .B1(new_n832), .B2(new_n851), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n821), .B(new_n445), .C1(new_n852), .C2(new_n834), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n853), .B1(new_n845), .B2(new_n821), .ZN(new_n854));
  INV_X1    g653(.A(new_n818), .ZN(new_n855));
  OR3_X1    g654(.A1(new_n854), .A2(new_n532), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n849), .B1(new_n856), .B2(G148gat), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n822), .A2(new_n836), .A3(new_n818), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n849), .B1(new_n858), .B2(new_n532), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n859), .A2(new_n311), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n848), .B1(new_n857), .B2(new_n860), .ZN(G1345gat));
  XOR2_X1   g660(.A(KEYINPUT79), .B(G155gat), .Z(new_n862));
  NOR3_X1   g661(.A1(new_n858), .A2(new_n862), .A3(new_n773), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n845), .A2(new_n557), .A3(new_n818), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n863), .B1(new_n862), .B2(new_n864), .ZN(G1346gat));
  NOR3_X1   g664(.A1(new_n846), .A2(G162gat), .A3(new_n588), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n866), .B(KEYINPUT120), .Z(new_n867));
  OAI21_X1  g666(.A(G162gat), .B1(new_n858), .B2(new_n588), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1347gat));
  NOR2_X1   g668(.A1(new_n621), .A2(new_n414), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n799), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(new_n615), .ZN(new_n872));
  XOR2_X1   g671(.A(new_n872), .B(G169gat), .Z(G1348gat));
  NOR2_X1   g672(.A1(new_n871), .A2(new_n532), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(new_n526), .ZN(G1349gat));
  NAND4_X1  g674(.A1(new_n799), .A2(new_n247), .A3(new_n557), .A4(new_n870), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n798), .A2(new_n679), .A3(new_n557), .A4(new_n870), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(G183gat), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT60), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n876), .A2(KEYINPUT121), .A3(new_n879), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n880), .A2(new_n881), .A3(KEYINPUT60), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(G1350gat));
  XNOR2_X1  g686(.A(KEYINPUT61), .B(G190gat), .ZN(new_n888));
  NAND2_X1  g687(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n871), .A2(new_n588), .ZN(new_n890));
  MUX2_X1   g689(.A(new_n888), .B(new_n889), .S(new_n890), .Z(G1351gat));
  NAND2_X1  g690(.A1(new_n644), .A2(new_n870), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n853), .B(new_n893), .C1(new_n845), .C2(new_n821), .ZN(new_n894));
  OAI21_X1  g693(.A(G197gat), .B1(new_n894), .B2(new_n615), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n845), .A2(new_n893), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n376), .A3(new_n614), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(G1352gat));
  XOR2_X1   g697(.A(KEYINPUT123), .B(G204gat), .Z(new_n899));
  OR2_X1    g698(.A1(new_n854), .A2(new_n532), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(new_n892), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n532), .A2(new_n899), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n896), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT62), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n903), .A2(KEYINPUT62), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n903), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n901), .A2(new_n906), .A3(new_n907), .A4(new_n908), .ZN(G1353gat));
  NOR2_X1   g708(.A1(new_n894), .A2(new_n773), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n912));
  OR2_X1    g711(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n911), .A2(G211gat), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n896), .A2(new_n379), .A3(new_n557), .ZN(new_n915));
  OAI211_X1 g714(.A(KEYINPUT125), .B(KEYINPUT63), .C1(new_n910), .C2(new_n379), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(G1354gat));
  OAI21_X1  g716(.A(G218gat), .B1(new_n894), .B2(new_n588), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n896), .A2(new_n380), .A3(new_n587), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT126), .ZN(G1355gat));
endmodule


