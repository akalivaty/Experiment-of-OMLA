//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  XNOR2_X1  g004(.A(G110), .B(G140), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n192), .A2(G227), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n191), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT65), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(new_n199), .A3(G143), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n200), .A2(new_n201), .A3(G128), .A4(new_n203), .ZN(new_n204));
  AND2_X1   g018(.A1(new_n200), .A2(new_n203), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n202), .A2(G146), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n206), .B1(new_n208), .B2(KEYINPUT1), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n204), .B1(new_n205), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G104), .ZN(new_n212));
  AND2_X1   g026(.A1(KEYINPUT79), .A2(G107), .ZN(new_n213));
  NOR2_X1   g027(.A1(KEYINPUT79), .A2(G107), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n212), .B1(new_n215), .B2(G104), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G101), .ZN(new_n217));
  INV_X1    g031(.A(G104), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(KEYINPUT3), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n220), .B1(new_n211), .B2(G104), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n215), .A2(new_n219), .B1(new_n212), .B2(new_n221), .ZN(new_n222));
  XOR2_X1   g036(.A(KEYINPUT80), .B(G101), .Z(new_n223));
  AOI21_X1  g037(.A(KEYINPUT81), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n214), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT79), .A2(G107), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n219), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n221), .A2(new_n212), .ZN(new_n228));
  AND4_X1   g042(.A1(KEYINPUT81), .A2(new_n227), .A3(new_n223), .A4(new_n228), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n210), .B(new_n217), .C1(new_n224), .C2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n222), .A2(KEYINPUT81), .A3(new_n223), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n227), .A2(new_n223), .A3(new_n228), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT81), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n231), .A2(new_n234), .B1(G101), .B2(new_n216), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n206), .B1(new_n200), .B2(KEYINPUT1), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n197), .A2(new_n199), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n207), .B1(new_n237), .B2(new_n202), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n204), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n230), .B1(new_n235), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G134), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT67), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G134), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(new_n244), .A3(G137), .ZN(new_n245));
  INV_X1    g059(.A(G137), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT68), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G137), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n247), .A2(new_n249), .A3(KEYINPUT11), .A4(G134), .ZN(new_n250));
  AOI21_X1  g064(.A(G137), .B1(new_n242), .B2(new_n244), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n245), .B(new_n250), .C1(new_n251), .C2(KEYINPUT11), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G131), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT67), .B(G134), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n254), .B1(new_n255), .B2(G137), .ZN(new_n256));
  INV_X1    g070(.A(G131), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n256), .A2(new_n257), .A3(new_n245), .A4(new_n250), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n240), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT12), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n240), .A2(KEYINPUT12), .A3(new_n259), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n200), .A2(KEYINPUT0), .A3(G128), .A4(new_n203), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT0), .B(G128), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n265), .B1(new_n238), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n227), .A2(new_n228), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(G101), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n270), .B1(new_n269), .B2(G101), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n272), .B1(new_n224), .B2(new_n229), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT82), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n231), .A2(new_n234), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT82), .B1(new_n276), .B2(new_n272), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n268), .B(new_n271), .C1(new_n275), .C2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n259), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT10), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT65), .B(G146), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n208), .B1(new_n281), .B2(G143), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n201), .B1(new_n281), .B2(G143), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n282), .B1(new_n283), .B2(new_n206), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n280), .B1(new_n284), .B2(new_n204), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n230), .A2(new_n280), .B1(new_n235), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n278), .A2(new_n279), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n195), .B1(new_n264), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n268), .A2(new_n271), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n273), .A2(new_n274), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n276), .A2(KEYINPUT82), .A3(new_n272), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n230), .A2(new_n280), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n235), .A2(new_n285), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n259), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n287), .A2(new_n296), .A3(new_n195), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n190), .B1(new_n288), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G469), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT73), .B(G902), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n279), .B1(new_n278), .B2(new_n286), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n292), .A2(new_n295), .A3(new_n259), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n194), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n264), .A2(new_n287), .A3(new_n195), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n301), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT83), .B(G469), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n189), .B1(new_n299), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G214), .B1(G237), .B2(G902), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n267), .A2(KEYINPUT86), .A3(G125), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT86), .B1(new_n267), .B2(G125), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT87), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n314), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT87), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(new_n312), .ZN(new_n318));
  INV_X1    g132(.A(G125), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n284), .A2(new_n319), .A3(new_n204), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n315), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(G224), .A3(new_n192), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n192), .A2(G224), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n315), .A2(new_n318), .A3(new_n323), .A4(new_n320), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(G110), .B(G122), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G119), .ZN(new_n328));
  OR3_X1    g142(.A1(new_n328), .A2(KEYINPUT71), .A3(G116), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT71), .B1(new_n328), .B2(G116), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XOR2_X1   g145(.A(KEYINPUT2), .B(G113), .Z(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT70), .B(G119), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G116), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n332), .B1(new_n331), .B2(new_n334), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n271), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n337), .B1(new_n290), .B2(new_n291), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n334), .A2(KEYINPUT5), .A3(new_n329), .A4(new_n330), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n334), .A2(KEYINPUT5), .ZN(new_n340));
  INV_X1    g154(.A(G113), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n335), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n235), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n327), .B1(new_n338), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n337), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n347), .B1(new_n275), .B2(new_n277), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n344), .A3(new_n326), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n346), .A2(new_n349), .A3(KEYINPUT6), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n326), .B1(new_n348), .B2(new_n344), .ZN(new_n351));
  XOR2_X1   g165(.A(KEYINPUT84), .B(KEYINPUT6), .Z(new_n352));
  AOI21_X1  g166(.A(KEYINPUT85), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n327), .B(new_n352), .C1(new_n338), .C2(new_n345), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT85), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n325), .B(new_n350), .C1(new_n353), .C2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT89), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n339), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n342), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n339), .A2(new_n358), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n235), .B1(new_n362), .B2(new_n335), .ZN(new_n363));
  XOR2_X1   g177(.A(KEYINPUT88), .B(KEYINPUT8), .Z(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(new_n326), .ZN(new_n365));
  INV_X1    g179(.A(new_n235), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n365), .B1(new_n366), .B2(new_n343), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n323), .A2(KEYINPUT7), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n316), .A2(new_n320), .A3(new_n312), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n363), .A2(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n370), .B(new_n349), .C1(new_n321), .C2(new_n368), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n371), .A2(new_n190), .ZN(new_n372));
  OAI21_X1  g186(.A(G210), .B1(G237), .B2(G902), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n357), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n373), .B1(new_n357), .B2(new_n372), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n311), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n310), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT90), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT72), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(G237), .ZN(new_n380));
  INV_X1    g194(.A(G237), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(KEYINPUT72), .ZN(new_n382));
  OAI211_X1 g196(.A(G214), .B(new_n192), .C1(new_n380), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n202), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(KEYINPUT72), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n379), .A2(G237), .ZN(new_n386));
  AOI21_X1  g200(.A(G953), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(G143), .A3(G214), .ZN(new_n388));
  NAND2_X1  g202(.A1(KEYINPUT18), .A2(G131), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n384), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G140), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G125), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n319), .A2(G140), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n281), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n396), .B1(new_n196), .B2(new_n395), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n390), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n389), .B1(new_n384), .B2(new_n388), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n378), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n385), .A2(new_n386), .ZN(new_n401));
  AND4_X1   g215(.A1(G143), .A2(new_n401), .A3(G214), .A4(new_n192), .ZN(new_n402));
  AOI21_X1  g216(.A(G143), .B1(new_n387), .B2(G214), .ZN(new_n403));
  OAI211_X1 g217(.A(KEYINPUT18), .B(G131), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n404), .A2(KEYINPUT90), .A3(new_n397), .A4(new_n390), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g220(.A(KEYINPUT17), .B(G131), .C1(new_n402), .C2(new_n403), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT91), .ZN(new_n408));
  OAI21_X1  g222(.A(G131), .B1(new_n402), .B2(new_n403), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT17), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n384), .A2(new_n257), .A3(new_n388), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n257), .B1(new_n384), .B2(new_n388), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT91), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT17), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT16), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(new_n391), .A3(G125), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n417), .B1(new_n394), .B2(new_n416), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n196), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT75), .ZN(new_n420));
  OAI211_X1 g234(.A(G146), .B(new_n417), .C1(new_n394), .C2(new_n416), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n418), .A2(KEYINPUT75), .A3(new_n196), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n408), .A2(new_n412), .A3(new_n415), .A4(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(G113), .B(G122), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n426), .B(new_n218), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n406), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT92), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n406), .A2(new_n425), .A3(KEYINPUT92), .A4(new_n427), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n427), .B1(new_n406), .B2(new_n425), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT93), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n436), .A3(new_n190), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n433), .B1(new_n430), .B2(new_n431), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT93), .B1(new_n438), .B2(G902), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n437), .A2(G475), .A3(new_n439), .ZN(new_n440));
  XOR2_X1   g254(.A(new_n421), .B(KEYINPUT76), .Z(new_n441));
  NAND2_X1  g255(.A1(new_n409), .A2(new_n411), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n394), .B(KEYINPUT19), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n441), .B(new_n442), .C1(new_n237), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n406), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n427), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n432), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT20), .ZN(new_n449));
  NOR2_X1   g263(.A1(G475), .A2(G902), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n430), .A2(new_n431), .B1(new_n446), .B2(new_n445), .ZN(new_n452));
  INV_X1    g266(.A(new_n450), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT20), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n440), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT94), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n440), .A2(KEYINPUT94), .A3(new_n455), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G952), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n461), .A2(KEYINPUT99), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(KEYINPUT99), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n192), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n464), .B1(G234), .B2(G237), .ZN(new_n465));
  AOI211_X1 g279(.A(new_n192), .B(new_n300), .C1(G234), .C2(G237), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(G898), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G478), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(KEYINPUT15), .ZN(new_n471));
  XNOR2_X1  g285(.A(G116), .B(G122), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n215), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n472), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(KEYINPUT14), .ZN(new_n475));
  INV_X1    g289(.A(G116), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(KEYINPUT14), .A3(G122), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G107), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n206), .A2(G143), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(KEYINPUT95), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n202), .A2(G128), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n255), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n255), .B1(new_n480), .B2(new_n481), .ZN(new_n484));
  OAI221_X1 g298(.A(new_n473), .B1(new_n475), .B2(new_n478), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT13), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n481), .A2(new_n486), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n480), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n487), .B1(new_n490), .B2(KEYINPUT96), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT96), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n241), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT97), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n225), .A2(new_n226), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n474), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n482), .A2(new_n495), .B1(new_n473), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n498), .B1(new_n495), .B2(new_n482), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n485), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G217), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n187), .A2(new_n501), .A3(G953), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n502), .B(new_n485), .C1(new_n494), .C2(new_n499), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n301), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT98), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI211_X1 g322(.A(KEYINPUT98), .B(new_n301), .C1(new_n504), .C2(new_n505), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n471), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI22_X1  g324(.A1(new_n506), .A2(new_n507), .B1(KEYINPUT15), .B2(new_n470), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n377), .A2(new_n460), .A3(new_n469), .A4(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n335), .A2(new_n336), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n259), .A2(new_n268), .ZN(new_n517));
  AOI21_X1  g331(.A(G134), .B1(new_n247), .B2(new_n249), .ZN(new_n518));
  OAI21_X1  g332(.A(G131), .B1(new_n251), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n239), .A2(new_n258), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(KEYINPUT30), .A3(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n519), .B1(new_n252), .B2(G131), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT69), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n522), .A2(new_n523), .B1(new_n204), .B2(new_n284), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n258), .A2(KEYINPUT69), .A3(new_n519), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT66), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n258), .A2(new_n253), .B1(new_n267), .B2(new_n526), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n265), .B(KEYINPUT66), .C1(new_n238), .C2(new_n266), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n524), .A2(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n516), .B(new_n521), .C1(new_n529), .C2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT29), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n387), .A2(G210), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(KEYINPUT27), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT26), .B(G101), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n520), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n267), .B1(new_n253), .B2(new_n258), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n537), .B1(new_n515), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n532), .A2(new_n533), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n522), .A2(new_n523), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n543), .A2(new_n525), .A3(new_n239), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n267), .A2(new_n526), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n259), .A2(new_n545), .A3(new_n528), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n516), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT28), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n549), .B1(new_n540), .B2(new_n515), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n517), .A2(new_n515), .A3(new_n520), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n551), .A2(KEYINPUT28), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n548), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n537), .B1(new_n553), .B2(KEYINPUT29), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n540), .A2(new_n549), .A3(new_n515), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n551), .A2(KEYINPUT28), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n516), .B1(new_n538), .B2(new_n539), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n533), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n300), .B(new_n542), .C1(new_n554), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G472), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n543), .A2(new_n525), .A3(new_n239), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n531), .B1(new_n562), .B2(new_n546), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT30), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n538), .A2(new_n539), .A3(new_n564), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n563), .A2(new_n515), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n537), .A2(new_n551), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT31), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  XOR2_X1   g382(.A(new_n535), .B(new_n536), .Z(new_n569));
  NAND2_X1  g383(.A1(new_n553), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT31), .ZN(new_n571));
  INV_X1    g385(.A(new_n567), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n532), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n568), .A2(new_n570), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT32), .ZN(new_n575));
  NOR2_X1   g389(.A1(G472), .A2(G902), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n575), .B1(new_n574), .B2(new_n576), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n561), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT74), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT23), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n581), .B1(new_n333), .B2(G128), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n328), .A2(new_n206), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n333), .B2(new_n206), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n582), .B1(new_n584), .B2(new_n581), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT24), .B(G110), .Z(new_n586));
  OAI22_X1  g400(.A1(new_n585), .A2(G110), .B1(new_n586), .B2(new_n584), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n441), .A2(new_n587), .A3(new_n396), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n585), .A2(G110), .B1(new_n586), .B2(new_n584), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n589), .A2(new_n423), .A3(new_n422), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT22), .B(G137), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n588), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n588), .A2(new_n590), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n593), .B(KEYINPUT77), .Z(new_n596));
  OAI211_X1 g410(.A(new_n300), .B(new_n594), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT25), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n501), .B1(new_n300), .B2(G234), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OR2_X1    g415(.A1(new_n595), .A2(new_n596), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n602), .A2(new_n594), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n600), .A2(G902), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT74), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n608), .B(new_n561), .C1(new_n577), .C2(new_n578), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n580), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT78), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n580), .A2(KEYINPUT78), .A3(new_n607), .A4(new_n609), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n514), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(new_n223), .ZN(G3));
  NOR2_X1   g429(.A1(new_n506), .A2(G478), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n504), .A2(new_n505), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT33), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n301), .A2(new_n470), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n460), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n532), .A2(new_n571), .A3(new_n572), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n571), .B1(new_n532), .B2(new_n572), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n537), .B1(new_n557), .B2(new_n548), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n576), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(G472), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n574), .B2(new_n300), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n309), .A2(new_n630), .A3(new_n607), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n469), .B(new_n311), .C1(new_n374), .C2(new_n375), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n621), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT34), .B(G104), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  NOR2_X1   g450(.A1(new_n513), .A2(new_n456), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G107), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  AND3_X1   g454(.A1(new_n440), .A2(KEYINPUT94), .A3(new_n455), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT94), .B1(new_n440), .B2(new_n455), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n469), .B(new_n513), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n357), .A2(new_n372), .ZN(new_n645));
  INV_X1    g459(.A(new_n373), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n357), .A2(new_n372), .A3(new_n373), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT36), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n596), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n595), .B(new_n651), .Z(new_n652));
  INV_X1    g466(.A(new_n604), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n600), .B2(new_n599), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n649), .A2(new_n309), .A3(new_n311), .A4(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n630), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n644), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT37), .B(G110), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  OAI21_X1  g476(.A(KEYINPUT32), .B1(new_n625), .B2(new_n626), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n608), .B1(new_n665), .B2(new_n561), .ZN(new_n666));
  INV_X1    g480(.A(new_n609), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n657), .ZN(new_n669));
  INV_X1    g483(.A(G900), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n465), .B1(new_n466), .B2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n668), .A2(new_n669), .A3(new_n637), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  NAND2_X1  g488(.A1(new_n541), .A2(new_n558), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n190), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n569), .B1(new_n532), .B2(new_n551), .ZN(new_n677));
  OAI21_X1  g491(.A(G472), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n665), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n512), .A2(new_n655), .A3(new_n311), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n641), .A2(new_n642), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n684), .B(KEYINPUT101), .Z(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n649), .B(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(KEYINPUT102), .B1(new_n683), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n687), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n689), .A2(new_n690), .A3(new_n682), .A4(new_n681), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n671), .B(new_n692), .Z(new_n693));
  NAND2_X1  g507(.A1(new_n309), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n694), .B(KEYINPUT40), .Z(new_n695));
  NAND3_X1  g509(.A1(new_n688), .A2(new_n691), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G143), .ZN(G45));
  NOR3_X1   g511(.A1(new_n657), .A2(new_n666), .A3(new_n667), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n699));
  INV_X1    g513(.A(new_n620), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n682), .A2(new_n699), .A3(new_n700), .A4(new_n672), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n458), .A2(new_n459), .A3(new_n700), .A4(new_n672), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(KEYINPUT104), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n698), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT105), .B(G146), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G48));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n304), .A2(new_n305), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n300), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n707), .B1(new_n709), .B2(G469), .ZN(new_n710));
  INV_X1    g524(.A(G469), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n306), .A2(KEYINPUT106), .A3(new_n711), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n188), .B(new_n308), .C1(new_n710), .C2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n714), .A2(new_n580), .A3(new_n607), .A4(new_n609), .ZN(new_n715));
  INV_X1    g529(.A(new_n632), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n682), .A2(new_n716), .A3(new_n700), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT41), .B(G113), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(KEYINPUT107), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n718), .B(new_n720), .ZN(G15));
  NAND2_X1  g535(.A1(new_n716), .A2(new_n637), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n715), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT108), .B(G116), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G18));
  NOR3_X1   g539(.A1(new_n713), .A2(new_n376), .A3(new_n655), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n644), .A2(new_n668), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  NOR2_X1   g542(.A1(new_n713), .A2(new_n468), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n649), .A2(new_n512), .A3(new_n311), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n622), .A2(new_n623), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n557), .A2(new_n558), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n569), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n626), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n606), .A2(new_n735), .A3(new_n629), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n729), .A2(new_n731), .A3(new_n682), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NOR2_X1   g552(.A1(new_n735), .A2(new_n629), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n656), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n713), .A2(new_n740), .A3(new_n376), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n701), .A2(new_n703), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G125), .ZN(G27));
  INV_X1    g557(.A(KEYINPUT42), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n580), .A2(new_n607), .A3(new_n609), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n647), .A2(new_n311), .A3(new_n648), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n310), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n701), .A2(new_n703), .A3(new_n745), .A4(new_n747), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n701), .A2(new_n703), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n606), .B1(new_n665), .B2(new_n561), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n747), .A2(KEYINPUT42), .A3(new_n750), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n744), .A2(new_n748), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n257), .ZN(G33));
  NAND4_X1  g567(.A1(new_n512), .A2(new_n440), .A3(new_n455), .A4(new_n672), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(KEYINPUT109), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n745), .A2(new_n755), .A3(new_n747), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G134), .ZN(G36));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n460), .B(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(KEYINPUT43), .A3(new_n700), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n761), .B1(new_n682), .B2(new_n620), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n658), .A3(new_n656), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n763), .A2(KEYINPUT44), .A3(new_n658), .A4(new_n656), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n287), .A2(new_n296), .A3(new_n195), .ZN(new_n768));
  INV_X1    g582(.A(new_n263), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT12), .B1(new_n240), .B2(new_n259), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n303), .ZN(new_n772));
  OAI211_X1 g586(.A(KEYINPUT45), .B(new_n768), .C1(new_n772), .C2(new_n195), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n774), .B1(new_n288), .B2(new_n297), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(new_n775), .A3(G469), .ZN(new_n776));
  NAND2_X1  g590(.A1(G469), .A2(G902), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT46), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n308), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT46), .B1(new_n776), .B2(new_n777), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n189), .ZN(new_n784));
  INV_X1    g598(.A(new_n746), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n784), .A2(new_n693), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n766), .A2(new_n767), .A3(new_n786), .ZN(new_n787));
  XOR2_X1   g601(.A(KEYINPUT111), .B(G137), .Z(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(G39));
  NAND2_X1  g603(.A1(new_n784), .A2(KEYINPUT47), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT47), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n791), .B1(new_n783), .B2(new_n189), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n668), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n746), .A2(new_n607), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n793), .A2(new_n794), .A3(new_n749), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G140), .ZN(G42));
  OAI21_X1  g611(.A(new_n513), .B1(new_n641), .B2(new_n642), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n458), .A2(new_n459), .A3(new_n620), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n633), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n727), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n612), .A2(new_n613), .ZN(new_n802));
  INV_X1    g616(.A(new_n514), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n729), .A2(new_n736), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n460), .A2(new_n730), .ZN(new_n806));
  AOI22_X1  g620(.A1(new_n805), .A2(new_n806), .B1(new_n644), .B2(new_n659), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n610), .A2(new_n713), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n808), .B(new_n716), .C1(new_n621), .C2(new_n637), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n801), .A2(new_n804), .A3(new_n807), .A4(new_n809), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n740), .A2(new_n310), .A3(new_n746), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n701), .A2(new_n703), .A3(new_n811), .ZN(new_n812));
  NOR4_X1   g626(.A1(new_n456), .A2(new_n512), .A3(new_n655), .A4(new_n671), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n668), .A2(new_n747), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n812), .A2(new_n756), .A3(new_n814), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n810), .A2(new_n752), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n309), .A2(new_n655), .A3(new_n672), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n679), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n806), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n704), .A2(new_n742), .A3(new_n673), .A4(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n816), .A2(new_n822), .A3(KEYINPUT53), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n748), .A2(new_n744), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n749), .A2(new_n751), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n815), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n806), .A2(new_n818), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n827), .B1(new_n749), .B2(new_n698), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n742), .A2(new_n673), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n829), .A3(new_n821), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n727), .A2(new_n660), .A3(new_n737), .A4(new_n800), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n715), .B1(new_n717), .B2(new_n722), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n831), .A2(new_n614), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n820), .A2(KEYINPUT52), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n826), .A2(new_n830), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n823), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT112), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n840), .B1(new_n835), .B2(new_n836), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n816), .A2(new_n822), .A3(KEYINPUT112), .A4(KEYINPUT53), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n841), .A2(new_n837), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n839), .B1(KEYINPUT54), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n465), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n760), .B2(new_n762), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n713), .A2(new_n376), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n847), .A3(new_n736), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n679), .A2(new_n607), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n713), .A2(new_n746), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n850), .A2(new_n465), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n464), .B1(new_n852), .B2(new_n621), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n848), .A2(new_n849), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n849), .B1(new_n848), .B2(new_n853), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n846), .A2(new_n750), .A3(new_n851), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n856), .A2(KEYINPUT48), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(KEYINPUT48), .ZN(new_n858));
  OAI22_X1  g672(.A1(new_n854), .A2(new_n855), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n740), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n846), .A2(new_n860), .A3(new_n851), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n852), .A2(new_n460), .A3(new_n620), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n846), .A2(new_n736), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n709), .A2(new_n707), .A3(G469), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT106), .B1(new_n306), .B2(new_n711), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n781), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n866), .A2(new_n189), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n785), .B1(new_n793), .B2(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n861), .B(new_n862), .C1(new_n863), .C2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT51), .ZN(new_n871));
  OR3_X1    g685(.A1(new_n713), .A2(KEYINPUT113), .A3(new_n311), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT113), .B1(new_n713), .B2(new_n311), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(new_n687), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT114), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n846), .A3(new_n736), .ZN(new_n876));
  XOR2_X1   g690(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n875), .A2(new_n846), .A3(new_n736), .A4(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n870), .A2(new_n871), .A3(new_n878), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n878), .A2(new_n880), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT51), .B1(new_n882), .B2(new_n869), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n859), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n844), .A2(KEYINPUT117), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n461), .A2(new_n192), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT117), .B1(new_n844), .B2(new_n884), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n759), .A2(new_n700), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT49), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n188), .B(new_n311), .C1(new_n866), .C2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(new_n890), .B2(new_n866), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(new_n687), .A3(new_n850), .ZN(new_n893));
  OAI22_X1  g707(.A1(new_n887), .A2(new_n888), .B1(new_n889), .B2(new_n893), .ZN(G75));
  AOI21_X1  g708(.A(new_n300), .B1(new_n823), .B2(new_n837), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT56), .B1(new_n895), .B2(new_n646), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n350), .B1(new_n353), .B2(new_n356), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(new_n325), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT55), .ZN(new_n899));
  OAI22_X1  g713(.A1(new_n896), .A2(new_n899), .B1(G952), .B2(new_n192), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n896), .A2(new_n899), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n901), .A2(KEYINPUT118), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(KEYINPUT118), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(G51));
  NOR2_X1   g718(.A1(new_n192), .A2(G952), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n823), .A2(new_n837), .A3(new_n838), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT120), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n823), .A2(new_n837), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT54), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n823), .A2(new_n837), .A3(new_n910), .A4(new_n838), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n907), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n777), .B(KEYINPUT119), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT57), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n708), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n895), .A2(G469), .A3(new_n773), .A4(new_n775), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n905), .B1(new_n916), .B2(new_n917), .ZN(G54));
  NAND3_X1  g732(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n919), .A2(new_n452), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(new_n452), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n920), .A2(new_n921), .A3(new_n905), .ZN(G60));
  NAND2_X1  g736(.A1(G478), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT59), .Z(new_n924));
  NAND2_X1  g738(.A1(new_n843), .A2(KEYINPUT54), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n924), .B1(new_n925), .B2(new_n906), .ZN(new_n926));
  OAI21_X1  g740(.A(KEYINPUT121), .B1(new_n926), .B2(new_n618), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT121), .ZN(new_n928));
  INV_X1    g742(.A(new_n618), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n928), .B(new_n929), .C1(new_n844), .C2(new_n924), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n924), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n905), .B1(new_n912), .B2(new_n931), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n927), .A2(new_n930), .A3(new_n932), .ZN(G63));
  NAND2_X1  g747(.A1(G217), .A2(G902), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT60), .Z(new_n935));
  NAND2_X1  g749(.A1(new_n908), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n603), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n905), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n652), .B(KEYINPUT122), .Z(new_n939));
  OAI21_X1  g753(.A(new_n938), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(G66));
  INV_X1    g756(.A(G224), .ZN(new_n943));
  OAI21_X1  g757(.A(G953), .B1(new_n467), .B2(new_n943), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT123), .Z(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n833), .B2(G953), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n897), .B1(G898), .B2(new_n192), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(G69));
  AOI21_X1  g762(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n704), .A2(new_n673), .A3(new_n742), .ZN(new_n951));
  INV_X1    g765(.A(new_n752), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n784), .A2(new_n693), .A3(new_n806), .A4(new_n750), .ZN(new_n953));
  AND4_X1   g767(.A1(new_n952), .A2(new_n796), .A3(new_n756), .A4(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n787), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n955), .A2(G953), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n563), .A2(new_n565), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(new_n443), .Z(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(new_n670), .B2(new_n192), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n798), .A2(new_n799), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n802), .A2(new_n693), .A3(new_n747), .A4(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n796), .B1(KEYINPUT124), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(KEYINPUT124), .B2(new_n961), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n787), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n951), .A2(new_n696), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT62), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n967), .A2(G953), .ZN(new_n968));
  OAI221_X1 g782(.A(new_n950), .B1(new_n956), .B2(new_n959), .C1(new_n968), .C2(new_n958), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n964), .A2(new_n966), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n958), .B1(new_n970), .B2(new_n192), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n956), .A2(new_n959), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n949), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n969), .A2(new_n973), .ZN(G72));
  NOR3_X1   g788(.A1(new_n964), .A2(new_n810), .A3(new_n966), .ZN(new_n975));
  NAND2_X1  g789(.A1(G472), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT63), .Z(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT125), .Z(new_n978));
  OAI21_X1  g792(.A(new_n677), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n978), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n955), .B2(new_n810), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n532), .A2(new_n541), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT126), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n905), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n979), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n982), .A2(new_n977), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n986), .A2(new_n677), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n843), .A2(new_n987), .ZN(new_n988));
  OR2_X1    g802(.A1(new_n988), .A2(KEYINPUT127), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(KEYINPUT127), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n985), .B1(new_n989), .B2(new_n990), .ZN(G57));
endmodule


