//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 0 1 1 0 1 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n551, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1139, new_n1140, new_n1141, new_n1142;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT66), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT67), .Z(new_n459));
  NAND2_X1  g034(.A1(new_n455), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  XNOR2_X1  g037(.A(KEYINPUT68), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n466), .B1(new_n463), .B2(new_n465), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n471), .A2(new_n475), .ZN(G160));
  INV_X1    g051(.A(new_n467), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n470), .ZN(new_n478));
  INV_X1    g053(.A(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(new_n470), .B2(G112), .ZN(new_n481));
  OAI22_X1  g056(.A1(new_n478), .A2(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n467), .A2(new_n470), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(G124), .B2(new_n483), .ZN(G162));
  AND2_X1   g059(.A1(new_n470), .A2(G138), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n466), .B(new_n485), .C1(new_n463), .C2(new_n465), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G2104), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n489), .A2(KEYINPUT68), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(KEYINPUT68), .ZN(new_n491));
  OAI21_X1  g066(.A(KEYINPUT3), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n492), .A2(KEYINPUT69), .A3(new_n466), .A4(new_n485), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n488), .A2(KEYINPUT4), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n472), .A2(new_n495), .A3(new_n485), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  AND3_X1   g072(.A1(new_n470), .A2(G102), .A3(G2104), .ZN(new_n498));
  NAND2_X1  g073(.A1(G114), .A2(G2104), .ZN(new_n499));
  INV_X1    g074(.A(G126), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n467), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n498), .B1(new_n501), .B2(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n497), .A2(KEYINPUT70), .A3(new_n502), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(G164));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n515), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  INV_X1    g098(.A(new_n517), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G89), .ZN(new_n525));
  INV_X1    g100(.A(new_n519), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n525), .A2(new_n527), .A3(new_n528), .A4(new_n530), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(KEYINPUT71), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(KEYINPUT71), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(G168));
  AOI22_X1  g109(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n514), .ZN(new_n536));
  XNOR2_X1  g111(.A(KEYINPUT72), .B(G90), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n517), .A2(new_n537), .B1(new_n519), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  XNOR2_X1  g116(.A(KEYINPUT73), .B(G43), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n517), .A2(new_n541), .B1(new_n519), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n543), .B(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n514), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  INV_X1    g130(.A(KEYINPUT75), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n556), .B(new_n557), .C1(new_n519), .C2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(G91), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n561));
  OAI221_X1 g136(.A(new_n559), .B1(new_n560), .B2(new_n517), .C1(new_n514), .C2(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(KEYINPUT75), .B1(new_n526), .B2(G53), .ZN(new_n563));
  NOR3_X1   g138(.A1(new_n519), .A2(new_n556), .A3(new_n558), .ZN(new_n564));
  NOR3_X1   g139(.A1(new_n563), .A2(new_n557), .A3(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  INV_X1    g143(.A(G168), .ZN(G286));
  NAND2_X1  g144(.A1(new_n524), .A2(G87), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n526), .A2(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(new_n526), .A2(G48), .ZN(new_n574));
  INV_X1    g149(.A(G86), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n517), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n512), .A2(G61), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT76), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n514), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n576), .A2(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n582), .A2(new_n514), .ZN(new_n583));
  INV_X1    g158(.A(G85), .ZN(new_n584));
  INV_X1    g159(.A(G47), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n517), .A2(new_n584), .B1(new_n519), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT77), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n587), .A2(KEYINPUT77), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n583), .B1(new_n589), .B2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n524), .A2(G92), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT10), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(new_n512), .ZN(new_n596));
  XNOR2_X1  g171(.A(KEYINPUT78), .B(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n594), .B1(G651), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n526), .A2(G54), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n601), .A2(KEYINPUT79), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(KEYINPUT79), .ZN(new_n603));
  AND2_X1   g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n592), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n592), .B1(new_n604), .B2(G868), .ZN(G321));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G868), .B2(new_n566), .ZN(G297));
  OAI21_X1  g183(.A(new_n607), .B1(G868), .B2(new_n566), .ZN(G280));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n604), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n604), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g190(.A(G135), .ZN(new_n616));
  NOR2_X1   g191(.A1(G99), .A2(G2105), .ZN(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(new_n470), .B2(G111), .ZN(new_n618));
  OAI22_X1  g193(.A1(new_n478), .A2(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(G123), .B2(new_n483), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT81), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NOR3_X1   g197(.A1(new_n490), .A2(new_n491), .A3(G2105), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(new_n472), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT80), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G2100), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT13), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n625), .B(new_n628), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n622), .B(new_n629), .C1(new_n626), .C2(G2100), .ZN(G156));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT15), .B(G2435), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(KEYINPUT14), .ZN(new_n635));
  XOR2_X1   g210(.A(G2451), .B(G2454), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G1341), .B(G1348), .Z(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT82), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n643), .B(G14), .C1(new_n641), .C2(new_n640), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(G401));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2072), .B(G2078), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT18), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(KEYINPUT83), .ZN(new_n651));
  OAI21_X1  g226(.A(KEYINPUT17), .B1(new_n651), .B2(new_n646), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(new_n648), .Z(new_n653));
  AND2_X1   g228(.A1(new_n651), .A2(new_n646), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2096), .B(G2100), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(G227));
  XNOR2_X1  g232(.A(G1971), .B(G1976), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  XOR2_X1   g234(.A(G1956), .B(G2474), .Z(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n659), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  AOI22_X1  g240(.A1(new_n663), .A2(KEYINPUT20), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n667), .A2(new_n659), .A3(new_n662), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n666), .B(new_n668), .C1(KEYINPUT20), .C2(new_n663), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1986), .B(G1996), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G1981), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G1991), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(G229));
  INV_X1    g250(.A(G16), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G23), .ZN(new_n677));
  INV_X1    g252(.A(G288), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n677), .B1(new_n678), .B2(new_n676), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT33), .Z(new_n680));
  OR2_X1    g255(.A1(new_n680), .A2(G1976), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(G1976), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n676), .A2(G6), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n576), .A2(new_n580), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(new_n684), .B2(new_n676), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT32), .B(G1981), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n676), .A2(G22), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G166), .B2(new_n676), .ZN(new_n689));
  INV_X1    g264(.A(G1971), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND4_X1  g266(.A1(new_n681), .A2(new_n682), .A3(new_n687), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(KEYINPUT34), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT85), .Z(new_n694));
  NAND2_X1  g269(.A1(new_n676), .A2(G24), .ZN(new_n695));
  INV_X1    g270(.A(G290), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n676), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT84), .B(G1986), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n692), .A2(KEYINPUT34), .ZN(new_n700));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G25), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n483), .A2(G119), .ZN(new_n703));
  OR2_X1    g278(.A1(G95), .A2(G2105), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n704), .B(G2104), .C1(G107), .C2(new_n470), .ZN(new_n705));
  INV_X1    g280(.A(G131), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n703), .B(new_n705), .C1(new_n478), .C2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n702), .B1(new_n708), .B2(new_n701), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT35), .B(G1991), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n709), .B(new_n710), .Z(new_n711));
  NAND4_X1  g286(.A1(new_n694), .A2(new_n699), .A3(new_n700), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT36), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT31), .B(G11), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n676), .A2(G4), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(new_n604), .B2(new_n676), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n716), .A2(G1348), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(G1348), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n719));
  NAND2_X1  g294(.A1(new_n701), .A2(G26), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n483), .A2(G128), .ZN(new_n722));
  OR2_X1    g297(.A1(G104), .A2(G2105), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n723), .B(G2104), .C1(G116), .C2(new_n470), .ZN(new_n724));
  INV_X1    g299(.A(G140), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n722), .B(new_n724), .C1(new_n478), .C2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n721), .B1(new_n727), .B2(new_n701), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G2067), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n676), .A2(G19), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n549), .B2(new_n676), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n731), .A2(G1341), .ZN(new_n732));
  NOR4_X1   g307(.A1(new_n717), .A2(new_n718), .A3(new_n729), .A4(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT25), .Z(new_n735));
  INV_X1    g310(.A(G139), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n478), .B2(new_n736), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT87), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n472), .A2(G127), .ZN(new_n739));
  INV_X1    g314(.A(G115), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(new_n489), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n738), .B1(G2105), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G29), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G29), .B2(G33), .ZN(new_n744));
  INV_X1    g319(.A(G2072), .ZN(new_n745));
  OR2_X1    g320(.A1(KEYINPUT24), .A2(G34), .ZN(new_n746));
  NAND2_X1  g321(.A1(KEYINPUT24), .A2(G34), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n746), .A2(new_n701), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G160), .B2(new_n701), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT88), .Z(new_n750));
  AOI22_X1  g325(.A1(new_n744), .A2(new_n745), .B1(G2084), .B2(new_n750), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(G2084), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n701), .A2(G35), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G162), .B2(new_n701), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT29), .Z(new_n755));
  INV_X1    g330(.A(G2090), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AND3_X1   g332(.A1(new_n751), .A2(new_n752), .A3(new_n757), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n731), .A2(G1341), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n744), .A2(new_n745), .ZN(new_n760));
  NOR2_X1   g335(.A1(G168), .A2(new_n676), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n676), .B2(G21), .ZN(new_n762));
  INV_X1    g337(.A(G1966), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT91), .ZN(new_n765));
  INV_X1    g340(.A(G28), .ZN(new_n766));
  NOR3_X1   g341(.A1(new_n765), .A2(new_n766), .A3(KEYINPUT30), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n765), .B1(new_n766), .B2(KEYINPUT30), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(new_n701), .ZN(new_n769));
  AOI211_X1 g344(.A(new_n767), .B(new_n769), .C1(KEYINPUT30), .C2(new_n766), .ZN(new_n770));
  NAND2_X1  g345(.A1(G171), .A2(G16), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G5), .B2(G16), .ZN(new_n772));
  INV_X1    g347(.A(G1961), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n764), .B(new_n774), .C1(new_n773), .C2(new_n772), .ZN(new_n775));
  OAI22_X1  g350(.A1(new_n762), .A2(new_n763), .B1(new_n701), .B2(new_n621), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n760), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n733), .A2(new_n758), .A3(new_n759), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n676), .A2(G20), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT23), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(KEYINPUT23), .B1(new_n566), .B2(new_n676), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(new_n779), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1956), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n756), .B2(new_n755), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT92), .Z(new_n786));
  NOR2_X1   g361(.A1(G27), .A2(G29), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G164), .B2(G29), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G2078), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n477), .A2(G141), .A3(new_n470), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT89), .Z(new_n791));
  NAND3_X1  g366(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT26), .Z(new_n793));
  AOI22_X1  g368(.A1(new_n483), .A2(G129), .B1(G105), .B2(new_n623), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n791), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  MUX2_X1   g370(.A(G32), .B(new_n795), .S(G29), .Z(new_n796));
  XOR2_X1   g371(.A(KEYINPUT27), .B(G1996), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT90), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n796), .B(new_n798), .ZN(new_n799));
  NOR4_X1   g374(.A1(new_n778), .A2(new_n786), .A3(new_n789), .A4(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n713), .A2(new_n714), .A3(new_n800), .ZN(G150));
  INV_X1    g376(.A(G150), .ZN(G311));
  AOI22_X1  g377(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n803), .A2(new_n514), .ZN(new_n804));
  INV_X1    g379(.A(G93), .ZN(new_n805));
  INV_X1    g380(.A(G55), .ZN(new_n806));
  OAI22_X1  g381(.A1(new_n517), .A2(new_n805), .B1(new_n519), .B2(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT93), .B(G860), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT37), .Z(new_n811));
  NAND2_X1  g386(.A1(new_n604), .A2(G559), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT38), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n549), .A2(new_n808), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n549), .A2(new_n808), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n813), .B(new_n818), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(KEYINPUT94), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(KEYINPUT94), .ZN(new_n822));
  INV_X1    g397(.A(new_n809), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n811), .B1(new_n824), .B2(new_n825), .ZN(G145));
  XNOR2_X1  g401(.A(new_n742), .B(new_n503), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n795), .B(new_n708), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n726), .B(new_n625), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  XOR2_X1   g406(.A(G162), .B(G160), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n621), .ZN(new_n833));
  INV_X1    g408(.A(G142), .ZN(new_n834));
  NOR2_X1   g409(.A1(G106), .A2(G2105), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(new_n470), .B2(G118), .ZN(new_n836));
  OAI22_X1  g411(.A1(new_n478), .A2(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(G130), .B2(new_n483), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n833), .B(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n831), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(G37), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g420(.A(new_n612), .B(new_n818), .ZN(new_n846));
  AOI21_X1  g421(.A(G299), .B1(new_n599), .B2(new_n600), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT98), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n599), .A2(G299), .A3(new_n600), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT97), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n846), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT41), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT99), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n849), .A2(KEYINPUT41), .A3(new_n851), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n852), .A2(KEYINPUT99), .A3(new_n855), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(new_n846), .ZN(new_n862));
  XNOR2_X1  g437(.A(G303), .B(G288), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n863), .A2(G305), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(G305), .ZN(new_n865));
  NOR3_X1   g440(.A1(new_n864), .A2(new_n865), .A3(G290), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(G290), .B1(new_n864), .B2(new_n865), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT42), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(KEYINPUT100), .A3(new_n868), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(KEYINPUT100), .B1(new_n867), .B2(new_n868), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT42), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n870), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n854), .A2(new_n862), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n876), .B1(new_n854), .B2(new_n862), .ZN(new_n878));
  OAI21_X1  g453(.A(G868), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n808), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n879), .B1(G868), .B2(new_n880), .ZN(G295));
  OAI21_X1  g456(.A(new_n879), .B1(G868), .B2(new_n880), .ZN(G331));
  INV_X1    g457(.A(KEYINPUT44), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(new_n872), .B2(new_n873), .ZN(new_n886));
  INV_X1    g461(.A(new_n873), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n887), .A2(KEYINPUT102), .A3(new_n871), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n817), .A2(G168), .ZN(new_n890));
  OAI21_X1  g465(.A(G286), .B1(new_n815), .B2(new_n816), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n890), .A2(new_n891), .A3(G171), .ZN(new_n892));
  AOI21_X1  g467(.A(G171), .B1(new_n890), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n852), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n859), .A2(new_n860), .A3(new_n894), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n889), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n884), .B1(new_n898), .B2(G37), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n896), .A2(new_n897), .ZN(new_n900));
  OAI211_X1 g475(.A(KEYINPUT103), .B(new_n843), .C1(new_n900), .C2(new_n889), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n896), .A2(new_n897), .A3(new_n874), .ZN(new_n902));
  XOR2_X1   g477(.A(KEYINPUT101), .B(KEYINPUT43), .Z(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n899), .A2(new_n901), .A3(new_n902), .A4(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n889), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n895), .B1(new_n856), .B2(new_n858), .ZN(new_n907));
  INV_X1    g482(.A(new_n896), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n909), .A2(new_n843), .A3(new_n902), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT43), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n883), .B1(new_n905), .B2(new_n911), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n899), .A2(new_n901), .A3(new_n902), .A4(new_n903), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n904), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT44), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n912), .A2(new_n915), .ZN(G397));
  NAND2_X1  g491(.A1(G160), .A2(G40), .ZN(new_n917));
  AOI21_X1  g492(.A(G1384), .B1(new_n497), .B2(new_n502), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n917), .A2(new_n918), .A3(KEYINPUT45), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n726), .B(G2067), .ZN(new_n921));
  XOR2_X1   g496(.A(new_n921), .B(KEYINPUT104), .Z(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n795), .B(G1996), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n707), .A2(new_n710), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT123), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n726), .A2(G2067), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n920), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n919), .B1(new_n923), .B2(new_n795), .ZN(new_n931));
  INV_X1    g506(.A(G1996), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n919), .B(new_n932), .C1(KEYINPUT124), .C2(KEYINPUT46), .ZN(new_n933));
  XNOR2_X1  g508(.A(KEYINPUT124), .B(KEYINPUT46), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(new_n920), .B2(G1996), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n931), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  XOR2_X1   g511(.A(new_n936), .B(KEYINPUT47), .Z(new_n937));
  NAND2_X1  g512(.A1(new_n707), .A2(new_n710), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n925), .A2(new_n938), .A3(new_n926), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n919), .ZN(new_n940));
  NOR2_X1   g515(.A1(G290), .A2(G1986), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n919), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(KEYINPUT48), .ZN(new_n943));
  AOI211_X1 g518(.A(new_n930), .B(new_n937), .C1(new_n940), .C2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT50), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n917), .B1(new_n918), .B2(new_n945), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n497), .A2(KEYINPUT70), .A3(new_n502), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT70), .B1(new_n497), .B2(new_n502), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n947), .A2(new_n948), .A3(G1384), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n946), .B1(new_n949), .B2(new_n945), .ZN(new_n950));
  INV_X1    g525(.A(G1348), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G40), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n471), .A2(new_n953), .A3(new_n475), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n918), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n955), .A2(G2067), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT112), .B1(new_n952), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(G1384), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n505), .A2(new_n959), .A3(new_n506), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT50), .ZN(new_n961));
  AOI21_X1  g536(.A(G1348), .B1(new_n961), .B2(new_n946), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n962), .A2(new_n963), .A3(new_n956), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT60), .B1(new_n958), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n602), .A2(new_n603), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(KEYINPUT116), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n952), .A2(KEYINPUT112), .A3(new_n957), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n963), .B1(new_n962), .B2(new_n956), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n970), .A2(KEYINPUT60), .ZN(new_n971));
  OR2_X1    g546(.A1(new_n966), .A2(KEYINPUT116), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n966), .A2(KEYINPUT116), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n970), .A2(new_n972), .A3(KEYINPUT60), .A4(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n967), .A2(new_n971), .A3(new_n974), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n505), .A2(new_n945), .A3(new_n959), .A4(new_n506), .ZN(new_n976));
  INV_X1    g551(.A(new_n918), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT50), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n976), .A2(new_n954), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G1956), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n960), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n918), .A2(KEYINPUT45), .ZN(new_n984));
  XNOR2_X1  g559(.A(KEYINPUT56), .B(G2072), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n983), .A2(new_n954), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  AND3_X1   g561(.A1(G299), .A2(KEYINPUT111), .A3(KEYINPUT57), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT57), .B1(G299), .B2(KEYINPUT111), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n981), .A2(new_n986), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n989), .B1(new_n981), .B2(new_n986), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n981), .A2(new_n986), .A3(new_n989), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT61), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n992), .B(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n954), .B(new_n984), .C1(new_n949), .C2(KEYINPUT45), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n997), .B1(new_n998), .B2(G1996), .ZN(new_n999));
  XOR2_X1   g574(.A(KEYINPUT58), .B(G1341), .Z(new_n1000));
  NAND2_X1  g575(.A1(new_n955), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n917), .B1(new_n960), .B2(new_n982), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n1002), .A2(KEYINPUT113), .A3(new_n932), .A4(new_n984), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n548), .A2(KEYINPUT114), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n1004), .A2(KEYINPUT59), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT59), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n975), .A2(new_n996), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n970), .A2(new_n966), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n993), .B1(new_n1010), .B2(new_n991), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n917), .B1(new_n977), .B2(new_n982), .ZN(new_n1013));
  INV_X1    g588(.A(G2078), .ZN(new_n1014));
  AND4_X1   g589(.A1(KEYINPUT53), .A2(new_n1013), .A3(new_n1014), .A4(new_n984), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n1015), .A2(KEYINPUT121), .ZN(new_n1016));
  AOI21_X1  g591(.A(G1961), .B1(new_n961), .B2(new_n946), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n1015), .B2(KEYINPUT121), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(new_n998), .B2(G2078), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT120), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1002), .A2(new_n1014), .A3(new_n984), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT120), .B1(new_n1023), .B2(new_n1019), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1016), .B(new_n1018), .C1(new_n1022), .C2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(G171), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1020), .B(new_n1021), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n959), .A4(new_n506), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1013), .A2(new_n1029), .A3(KEYINPUT53), .A4(new_n1014), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1028), .B1(new_n1031), .B2(new_n1017), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n950), .A2(new_n773), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1033), .A2(KEYINPUT119), .A3(new_n1030), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1027), .A2(G301), .A3(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1026), .A2(new_n1036), .A3(KEYINPUT54), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n998), .A2(new_n690), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n756), .B(new_n946), .C1(new_n949), .C2(new_n945), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT105), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n961), .A2(KEYINPUT105), .A3(new_n756), .A4(new_n946), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1038), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(G303), .A2(G8), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT106), .ZN(new_n1047));
  NAND3_X1  g622(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT106), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1044), .A2(new_n1049), .A3(new_n1045), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1047), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT107), .ZN(new_n1052));
  XNOR2_X1  g627(.A(new_n1051), .B(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1043), .A2(G8), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(G1971), .B1(new_n1002), .B2(new_n984), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n979), .A2(G2090), .ZN(new_n1056));
  OAI21_X1  g631(.A(G8), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1051), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G8), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1060), .B1(new_n918), .B2(new_n954), .ZN(new_n1061));
  INV_X1    g636(.A(G1976), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(new_n1062), .B2(G288), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT52), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1064), .B1(new_n678), .B2(G1976), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1061), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT49), .ZN(new_n1068));
  NAND3_X1  g643(.A1(G305), .A2(new_n1068), .A3(G1981), .ZN(new_n1069));
  INV_X1    g644(.A(G1981), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT49), .B1(new_n684), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT109), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1073), .B1(new_n684), .B2(new_n1070), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1069), .A2(new_n1074), .A3(new_n1071), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1067), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1063), .A2(KEYINPUT52), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT108), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1063), .A2(KEYINPUT108), .A3(KEYINPUT52), .ZN(new_n1082));
  AOI211_X1 g657(.A(new_n1066), .B(new_n1078), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1054), .A2(new_n1059), .A3(new_n1083), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1037), .A2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(G168), .A2(new_n1060), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(KEYINPUT117), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(G1966), .B1(new_n1013), .B2(new_n1029), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G2084), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1091), .B(new_n946), .C1(new_n949), .C2(new_n945), .ZN(new_n1092));
  NAND2_X1  g667(.A1(KEYINPUT118), .A2(KEYINPUT51), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1088), .A2(new_n1090), .A3(new_n1092), .A4(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1092), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1096), .B(G8), .C1(new_n1097), .C2(new_n1089), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1087), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1093), .B1(new_n1100), .B2(G8), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1095), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1035), .B1(new_n1024), .B2(new_n1022), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(G171), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(G171), .B2(new_n1025), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1102), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1012), .A2(new_n1085), .A3(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1083), .A2(G8), .A3(new_n1043), .A4(new_n1053), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1102), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(G301), .B1(new_n1027), .B2(new_n1035), .ZN(new_n1112));
  OAI211_X1 g687(.A(KEYINPUT62), .B(new_n1095), .C1(new_n1099), .C2(new_n1101), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1111), .A2(new_n1084), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT63), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1043), .A2(G8), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1115), .B1(new_n1116), .B2(new_n1058), .ZN(new_n1117));
  AOI211_X1 g692(.A(new_n1060), .B(G286), .C1(new_n1090), .C2(new_n1092), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1117), .A2(new_n1054), .A3(new_n1083), .A4(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1054), .A2(new_n1059), .A3(new_n1083), .A4(new_n1118), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1115), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(G288), .A2(G1976), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1123), .B(KEYINPUT110), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1076), .A2(new_n1077), .A3(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(G1981), .B2(G305), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n1061), .ZN(new_n1127));
  AND4_X1   g702(.A1(new_n1109), .A2(new_n1114), .A3(new_n1122), .A4(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1108), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n939), .B1(G1986), .B2(G290), .ZN(new_n1130));
  INV_X1    g705(.A(new_n941), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n920), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT122), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n1135));
  AOI211_X1 g710(.A(new_n1135), .B(new_n1132), .C1(new_n1108), .C2(new_n1128), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n944), .B1(new_n1134), .B2(new_n1136), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g712(.A1(G227), .A2(new_n461), .ZN(new_n1139));
  AOI21_X1  g713(.A(G229), .B1(new_n1139), .B2(KEYINPUT125), .ZN(new_n1140));
  OAI211_X1 g714(.A(new_n644), .B(new_n1140), .C1(KEYINPUT125), .C2(new_n1139), .ZN(new_n1141));
  XNOR2_X1  g715(.A(new_n1141), .B(KEYINPUT126), .ZN(new_n1142));
  NAND4_X1  g716(.A1(new_n913), .A2(new_n914), .A3(new_n844), .A4(new_n1142), .ZN(G225));
  INV_X1    g717(.A(G225), .ZN(G308));
endmodule


