

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770;

  AND2_X1 U380 ( .A1(n632), .A2(n633), .ZN(n377) );
  XNOR2_X2 U381 ( .A(G116), .B(KEYINPUT3), .ZN(n422) );
  INV_X2 U382 ( .A(G104), .ZN(n416) );
  XNOR2_X2 U383 ( .A(n552), .B(KEYINPUT19), .ZN(n594) );
  NOR2_X2 U384 ( .A1(n658), .A2(n743), .ZN(n659) );
  XNOR2_X2 U385 ( .A(n416), .B(G113), .ZN(n502) );
  XNOR2_X1 U386 ( .A(n411), .B(n366), .ZN(n586) );
  NOR2_X1 U387 ( .A1(n695), .A2(n584), .ZN(n585) );
  AND2_X1 U388 ( .A1(n616), .A2(n653), .ZN(n633) );
  XNOR2_X1 U389 ( .A(n555), .B(KEYINPUT117), .ZN(n765) );
  OR2_X1 U390 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U391 ( .A(n491), .B(n490), .ZN(n686) );
  XNOR2_X1 U392 ( .A(n756), .B(G146), .ZN(n392) );
  XNOR2_X2 U393 ( .A(n441), .B(KEYINPUT88), .ZN(n552) );
  NAND2_X1 U394 ( .A1(n404), .A2(n402), .ZN(n541) );
  NOR2_X1 U395 ( .A1(n770), .A2(n533), .ZN(n402) );
  XNOR2_X1 U396 ( .A(n518), .B(n445), .ZN(n756) );
  XNOR2_X1 U397 ( .A(KEYINPUT4), .B(G137), .ZN(n444) );
  XNOR2_X1 U398 ( .A(G131), .B(KEYINPUT70), .ZN(n443) );
  NAND2_X1 U399 ( .A1(n660), .A2(n505), .ZN(n454) );
  INV_X1 U400 ( .A(KEYINPUT106), .ZN(n560) );
  OR2_X1 U401 ( .A1(n559), .A2(n558), .ZN(n561) );
  NOR2_X1 U402 ( .A1(n622), .A2(n614), .ZN(n697) );
  XNOR2_X1 U403 ( .A(n599), .B(n549), .ZN(n617) );
  NOR2_X1 U404 ( .A1(n541), .A2(n540), .ZN(n548) );
  XNOR2_X1 U405 ( .A(n765), .B(n393), .ZN(n410) );
  INV_X1 U406 ( .A(KEYINPUT84), .ZN(n393) );
  NOR2_X1 U407 ( .A1(n587), .A2(n760), .ZN(n462) );
  NAND2_X1 U408 ( .A1(n585), .A2(n643), .ZN(n395) );
  XNOR2_X1 U409 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n429) );
  XOR2_X1 U410 ( .A(KEYINPUT18), .B(KEYINPUT89), .Z(n430) );
  XNOR2_X1 U411 ( .A(G146), .B(G125), .ZN(n466) );
  INV_X1 U412 ( .A(n442), .ZN(n368) );
  XNOR2_X1 U413 ( .A(n438), .B(n437), .ZN(n525) );
  XNOR2_X1 U414 ( .A(n436), .B(KEYINPUT90), .ZN(n437) );
  NAND2_X1 U415 ( .A1(n525), .A2(n575), .ZN(n441) );
  XNOR2_X1 U416 ( .A(n392), .B(n487), .ZN(n647) );
  XOR2_X1 U417 ( .A(KEYINPUT5), .B(G113), .Z(n484) );
  NAND2_X1 U418 ( .A1(n386), .A2(n585), .ZN(n391) );
  INV_X1 U419 ( .A(n586), .ZN(n386) );
  XNOR2_X1 U420 ( .A(n415), .B(G107), .ZN(n426) );
  INV_X1 U421 ( .A(G122), .ZN(n415) );
  XNOR2_X1 U422 ( .A(G110), .B(G107), .ZN(n448) );
  XNOR2_X1 U423 ( .A(G104), .B(G101), .ZN(n446) );
  XNOR2_X1 U424 ( .A(n645), .B(KEYINPUT76), .ZN(n729) );
  NAND2_X1 U425 ( .A1(n585), .A2(KEYINPUT2), .ZN(n387) );
  XNOR2_X1 U426 ( .A(n409), .B(KEYINPUT110), .ZN(n576) );
  INV_X1 U427 ( .A(KEYINPUT1), .ZN(n382) );
  INV_X1 U428 ( .A(n702), .ZN(n370) );
  BUF_X1 U429 ( .A(n525), .Z(n582) );
  NAND2_X1 U430 ( .A1(n384), .A2(n360), .ZN(n572) );
  AND2_X1 U431 ( .A1(n531), .A2(n385), .ZN(n384) );
  XNOR2_X1 U432 ( .A(n481), .B(n480), .ZN(n622) );
  XNOR2_X1 U433 ( .A(n479), .B(n420), .ZN(n480) );
  XNOR2_X1 U434 ( .A(n417), .B(n364), .ZN(n621) );
  AND2_X1 U435 ( .A1(n715), .A2(n419), .ZN(n418) );
  NAND2_X1 U436 ( .A1(n734), .A2(n588), .ZN(n407) );
  INV_X1 U437 ( .A(KEYINPUT80), .ZN(n405) );
  NOR2_X1 U438 ( .A1(n769), .A2(n767), .ZN(n374) );
  NOR2_X1 U439 ( .A1(n556), .A2(KEYINPUT71), .ZN(n398) );
  NAND2_X1 U440 ( .A1(G234), .A2(G237), .ZN(n457) );
  XNOR2_X1 U441 ( .A(KEYINPUT14), .B(KEYINPUT92), .ZN(n458) );
  NOR2_X1 U442 ( .A1(n590), .A2(n358), .ZN(n528) );
  INV_X1 U443 ( .A(n614), .ZN(n419) );
  XNOR2_X1 U444 ( .A(n469), .B(n468), .ZN(n510) );
  XOR2_X1 U445 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n468) );
  XNOR2_X1 U446 ( .A(G110), .B(KEYINPUT24), .ZN(n471) );
  XNOR2_X1 U447 ( .A(G128), .B(G137), .ZN(n470) );
  XNOR2_X1 U448 ( .A(G116), .B(KEYINPUT7), .ZN(n515) );
  XOR2_X1 U449 ( .A(KEYINPUT9), .B(KEYINPUT104), .Z(n516) );
  INV_X1 U450 ( .A(KEYINPUT103), .ZN(n511) );
  XNOR2_X1 U451 ( .A(n426), .B(n414), .ZN(n512) );
  INV_X1 U452 ( .A(KEYINPUT102), .ZN(n414) );
  XNOR2_X1 U453 ( .A(n442), .B(G134), .ZN(n518) );
  XNOR2_X1 U454 ( .A(n466), .B(KEYINPUT10), .ZN(n500) );
  XNOR2_X1 U455 ( .A(G143), .B(G131), .ZN(n496) );
  XOR2_X1 U456 ( .A(G122), .B(G140), .Z(n497) );
  XNOR2_X1 U457 ( .A(n373), .B(n372), .ZN(n646) );
  INV_X1 U458 ( .A(KEYINPUT65), .ZN(n372) );
  NAND2_X1 U459 ( .A1(n396), .A2(n365), .ZN(n373) );
  XNOR2_X1 U460 ( .A(n369), .B(n368), .ZN(n433) );
  AND2_X1 U461 ( .A1(n698), .A2(n697), .ZN(n367) );
  XNOR2_X1 U462 ( .A(n564), .B(KEYINPUT41), .ZN(n733) );
  XNOR2_X1 U463 ( .A(n383), .B(n573), .ZN(n583) );
  NOR2_X1 U464 ( .A1(n572), .A2(n713), .ZN(n383) );
  XNOR2_X1 U465 ( .A(n376), .B(n375), .ZN(n566) );
  INV_X1 U466 ( .A(KEYINPUT28), .ZN(n375) );
  NOR2_X1 U467 ( .A1(n550), .A2(n700), .ZN(n376) );
  OR2_X1 U468 ( .A1(n647), .A2(G902), .ZN(n488) );
  INV_X1 U469 ( .A(n759), .ZN(n390) );
  BUF_X1 U470 ( .A(n665), .Z(n739) );
  XNOR2_X1 U471 ( .A(n392), .B(n452), .ZN(n660) );
  NOR2_X1 U472 ( .A1(n576), .A2(n552), .ZN(n553) );
  NOR2_X1 U473 ( .A1(n619), .A2(n615), .ZN(n620) );
  NAND2_X1 U474 ( .A1(n371), .A2(n363), .ZN(n619) );
  XNOR2_X1 U475 ( .A(n403), .B(KEYINPUT114), .ZN(n770) );
  NOR2_X1 U476 ( .A1(n572), .A2(n532), .ZN(n403) );
  NAND2_X1 U477 ( .A1(n380), .A2(n378), .ZN(n653) );
  NOR2_X1 U478 ( .A1(n702), .A2(n379), .ZN(n378) );
  INV_X1 U479 ( .A(n615), .ZN(n379) );
  AND2_X1 U480 ( .A1(n408), .A2(n406), .ZN(n735) );
  NOR2_X1 U481 ( .A1(n731), .A2(n407), .ZN(n406) );
  XNOR2_X1 U482 ( .A(n730), .B(KEYINPUT82), .ZN(n408) );
  XOR2_X1 U483 ( .A(KEYINPUT109), .B(n464), .Z(n358) );
  NOR2_X1 U484 ( .A1(n708), .A2(n707), .ZN(n359) );
  XOR2_X1 U485 ( .A(n527), .B(n526), .Z(n360) );
  NOR2_X1 U486 ( .A1(n557), .A2(n524), .ZN(n361) );
  AND2_X1 U487 ( .A1(n551), .A2(n689), .ZN(n362) );
  NOR2_X1 U488 ( .A1(n618), .A2(n370), .ZN(n363) );
  XOR2_X1 U489 ( .A(KEYINPUT75), .B(KEYINPUT22), .Z(n364) );
  XNOR2_X1 U490 ( .A(KEYINPUT66), .B(n644), .ZN(n365) );
  XOR2_X1 U491 ( .A(KEYINPUT48), .B(KEYINPUT83), .Z(n366) );
  OR2_X1 U492 ( .A1(n760), .A2(G952), .ZN(n671) );
  INV_X1 U493 ( .A(KEYINPUT2), .ZN(n388) );
  XNOR2_X1 U494 ( .A(n381), .B(KEYINPUT86), .ZN(n380) );
  NAND2_X1 U495 ( .A1(n367), .A2(n617), .ZN(n604) );
  NAND2_X1 U496 ( .A1(n760), .A2(G224), .ZN(n369) );
  INV_X1 U497 ( .A(n621), .ZN(n371) );
  NAND2_X1 U498 ( .A1(n583), .A2(n689), .ZN(n574) );
  XNOR2_X1 U499 ( .A(n374), .B(KEYINPUT46), .ZN(n412) );
  NAND2_X1 U500 ( .A1(n377), .A2(n640), .ZN(n641) );
  INV_X1 U501 ( .A(n556), .ZN(n401) );
  NAND2_X1 U502 ( .A1(n548), .A2(n547), .ZN(n556) );
  XNOR2_X1 U503 ( .A(n458), .B(n457), .ZN(n460) );
  NOR2_X1 U504 ( .A1(n621), .A2(n617), .ZN(n381) );
  XNOR2_X2 U505 ( .A(n565), .B(n382), .ZN(n698) );
  INV_X1 U506 ( .A(n528), .ZN(n385) );
  NOR2_X1 U507 ( .A1(n586), .A2(n387), .ZN(n421) );
  NAND2_X1 U508 ( .A1(n389), .A2(n744), .ZN(n727) );
  INV_X1 U509 ( .A(n391), .ZN(n389) );
  XNOR2_X1 U510 ( .A(n391), .B(n390), .ZN(n761) );
  NAND2_X1 U511 ( .A1(n362), .A2(n617), .ZN(n409) );
  XNOR2_X2 U512 ( .A(n488), .B(G472), .ZN(n599) );
  NAND2_X1 U513 ( .A1(n394), .A2(n744), .ZN(n396) );
  XNOR2_X2 U514 ( .A(n641), .B(KEYINPUT45), .ZN(n744) );
  NOR2_X1 U515 ( .A1(n586), .A2(n395), .ZN(n394) );
  NAND2_X1 U516 ( .A1(n399), .A2(n397), .ZN(n413) );
  NAND2_X1 U517 ( .A1(n398), .A2(n410), .ZN(n397) );
  NAND2_X1 U518 ( .A1(n400), .A2(KEYINPUT71), .ZN(n399) );
  NAND2_X1 U519 ( .A1(n401), .A2(n410), .ZN(n400) );
  INV_X1 U520 ( .A(n686), .ZN(n543) );
  NAND2_X1 U521 ( .A1(n686), .A2(n405), .ZN(n404) );
  NAND2_X1 U522 ( .A1(n413), .A2(n412), .ZN(n411) );
  XNOR2_X1 U523 ( .A(n502), .B(G110), .ZN(n425) );
  NAND2_X1 U524 ( .A1(n418), .A2(n605), .ZN(n417) );
  XNOR2_X2 U525 ( .A(n596), .B(n595), .ZN(n605) );
  XNOR2_X1 U526 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X2 U527 ( .A(n454), .B(n453), .ZN(n565) );
  BUF_X1 U528 ( .A(n666), .Z(n668) );
  NAND2_X1 U529 ( .A1(n715), .A2(n563), .ZN(n564) );
  XOR2_X1 U530 ( .A(KEYINPUT25), .B(KEYINPUT96), .Z(n420) );
  INV_X1 U531 ( .A(KEYINPUT116), .ZN(n570) );
  NOR2_X2 U532 ( .A1(n557), .A2(n559), .ZN(n689) );
  INV_X1 U533 ( .A(n422), .ZN(n424) );
  XNOR2_X1 U534 ( .A(G101), .B(G119), .ZN(n423) );
  XNOR2_X1 U535 ( .A(n424), .B(n423), .ZN(n486) );
  XNOR2_X1 U536 ( .A(n425), .B(n486), .ZN(n428) );
  XOR2_X1 U537 ( .A(KEYINPUT16), .B(n426), .Z(n427) );
  XNOR2_X1 U538 ( .A(n428), .B(n427), .ZN(n751) );
  XNOR2_X1 U539 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U540 ( .A(n466), .B(n431), .ZN(n434) );
  INV_X1 U541 ( .A(KEYINPUT64), .ZN(n432) );
  XNOR2_X2 U542 ( .A(n432), .B(G953), .ZN(n760) );
  XNOR2_X2 U543 ( .A(G143), .B(G128), .ZN(n442) );
  XNOR2_X1 U544 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U545 ( .A(n751), .B(n435), .ZN(n666) );
  XNOR2_X1 U546 ( .A(KEYINPUT15), .B(G902), .ZN(n642) );
  NAND2_X1 U547 ( .A1(n666), .A2(n642), .ZN(n438) );
  OR2_X1 U548 ( .A1(G237), .A2(G902), .ZN(n439) );
  AND2_X1 U549 ( .A1(G210), .A2(n439), .ZN(n436) );
  NAND2_X1 U550 ( .A1(G214), .A2(n439), .ZN(n440) );
  XOR2_X1 U551 ( .A(KEYINPUT91), .B(n440), .Z(n575) );
  XNOR2_X1 U552 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U553 ( .A(KEYINPUT69), .B(G140), .Z(n467) );
  XNOR2_X1 U554 ( .A(n446), .B(KEYINPUT94), .ZN(n447) );
  XNOR2_X1 U555 ( .A(n467), .B(n447), .ZN(n451) );
  NAND2_X1 U556 ( .A1(n760), .A2(G227), .ZN(n449) );
  XNOR2_X1 U557 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U558 ( .A(n451), .B(n450), .ZN(n452) );
  INV_X1 U559 ( .A(G902), .ZN(n505) );
  XNOR2_X1 U560 ( .A(KEYINPUT73), .B(G469), .ZN(n453) );
  INV_X1 U561 ( .A(n565), .ZN(n530) );
  NAND2_X1 U562 ( .A1(n594), .A2(n530), .ZN(n489) );
  NAND2_X1 U563 ( .A1(n642), .A2(G234), .ZN(n455) );
  XNOR2_X1 U564 ( .A(n455), .B(KEYINPUT20), .ZN(n478) );
  NAND2_X1 U565 ( .A1(n478), .A2(G221), .ZN(n456) );
  XNOR2_X1 U566 ( .A(KEYINPUT21), .B(n456), .ZN(n703) );
  NAND2_X1 U567 ( .A1(n460), .A2(G952), .ZN(n459) );
  XOR2_X1 U568 ( .A(KEYINPUT93), .B(n459), .Z(n726) );
  NOR2_X1 U569 ( .A1(G953), .A2(n726), .ZN(n590) );
  NAND2_X1 U570 ( .A1(G902), .A2(n460), .ZN(n587) );
  INV_X1 U571 ( .A(KEYINPUT108), .ZN(n461) );
  XNOR2_X1 U572 ( .A(n462), .B(n461), .ZN(n463) );
  NOR2_X1 U573 ( .A1(G900), .A2(n463), .ZN(n464) );
  NOR2_X1 U574 ( .A1(n703), .A2(n528), .ZN(n465) );
  XNOR2_X1 U575 ( .A(n465), .B(KEYINPUT72), .ZN(n482) );
  XOR2_X1 U576 ( .A(n467), .B(n500), .Z(n755) );
  NAND2_X1 U577 ( .A1(G234), .A2(n760), .ZN(n469) );
  NAND2_X1 U578 ( .A1(n510), .A2(G221), .ZN(n476) );
  XNOR2_X1 U579 ( .A(n470), .B(G119), .ZN(n474) );
  XOR2_X1 U580 ( .A(KEYINPUT23), .B(KEYINPUT95), .Z(n472) );
  XNOR2_X1 U581 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U582 ( .A(n474), .B(n473), .Z(n475) );
  XNOR2_X1 U583 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U584 ( .A(n477), .B(n755), .ZN(n740) );
  NOR2_X1 U585 ( .A1(n740), .A2(G902), .ZN(n481) );
  NAND2_X1 U586 ( .A1(n478), .A2(G217), .ZN(n479) );
  NAND2_X1 U587 ( .A1(n482), .A2(n622), .ZN(n550) );
  NOR2_X1 U588 ( .A1(G953), .A2(G237), .ZN(n492) );
  NAND2_X1 U589 ( .A1(n492), .A2(G210), .ZN(n483) );
  XNOR2_X1 U590 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U591 ( .A(n486), .B(n485), .ZN(n487) );
  INV_X1 U592 ( .A(n599), .ZN(n700) );
  NOR2_X1 U593 ( .A1(n489), .A2(n566), .ZN(n491) );
  INV_X1 U594 ( .A(KEYINPUT79), .ZN(n490) );
  NAND2_X1 U595 ( .A1(G214), .A2(n492), .ZN(n494) );
  XOR2_X1 U596 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n493) );
  XNOR2_X1 U597 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U598 ( .A(n495), .B(KEYINPUT98), .Z(n499) );
  XNOR2_X1 U599 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U600 ( .A(n499), .B(n498), .ZN(n504) );
  INV_X1 U601 ( .A(n500), .ZN(n501) );
  XOR2_X1 U602 ( .A(n502), .B(n501), .Z(n503) );
  XNOR2_X1 U603 ( .A(n504), .B(n503), .ZN(n655) );
  NAND2_X1 U604 ( .A1(n655), .A2(n505), .ZN(n509) );
  XOR2_X1 U605 ( .A(KEYINPUT100), .B(KEYINPUT13), .Z(n507) );
  XNOR2_X1 U606 ( .A(KEYINPUT99), .B(G475), .ZN(n506) );
  XNOR2_X1 U607 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X2 U608 ( .A(n509), .B(n508), .ZN(n557) );
  NAND2_X1 U609 ( .A1(G217), .A2(n510), .ZN(n514) );
  XNOR2_X1 U610 ( .A(n514), .B(n513), .ZN(n521) );
  XNOR2_X1 U611 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U612 ( .A(n517), .B(KEYINPUT101), .ZN(n519) );
  XNOR2_X1 U613 ( .A(n518), .B(n519), .ZN(n520) );
  XNOR2_X1 U614 ( .A(n521), .B(n520), .ZN(n736) );
  INV_X1 U615 ( .A(n736), .ZN(n522) );
  NAND2_X1 U616 ( .A1(n522), .A2(n505), .ZN(n523) );
  XNOR2_X1 U617 ( .A(n523), .B(G478), .ZN(n559) );
  AND2_X1 U618 ( .A1(n557), .A2(n559), .ZN(n691) );
  NOR2_X1 U619 ( .A1(n689), .A2(n691), .ZN(n712) );
  INV_X1 U620 ( .A(n712), .ZN(n542) );
  AND2_X1 U621 ( .A1(KEYINPUT81), .A2(n542), .ZN(n533) );
  INV_X1 U622 ( .A(n559), .ZN(n524) );
  NAND2_X1 U623 ( .A1(n361), .A2(n582), .ZN(n532) );
  XOR2_X1 U624 ( .A(KEYINPUT113), .B(KEYINPUT30), .Z(n527) );
  NAND2_X1 U625 ( .A1(n599), .A2(n575), .ZN(n526) );
  INV_X1 U626 ( .A(KEYINPUT97), .ZN(n529) );
  XNOR2_X1 U627 ( .A(n703), .B(n529), .ZN(n614) );
  NAND2_X1 U628 ( .A1(n697), .A2(n530), .ZN(n600) );
  INV_X1 U629 ( .A(n600), .ZN(n531) );
  INV_X1 U630 ( .A(KEYINPUT47), .ZN(n537) );
  AND2_X1 U631 ( .A1(n542), .A2(n537), .ZN(n534) );
  AND2_X1 U632 ( .A1(n686), .A2(n534), .ZN(n539) );
  INV_X1 U633 ( .A(KEYINPUT81), .ZN(n535) );
  NAND2_X1 U634 ( .A1(KEYINPUT80), .A2(n535), .ZN(n536) );
  AND2_X1 U635 ( .A1(n537), .A2(n536), .ZN(n538) );
  OR2_X1 U636 ( .A1(n542), .A2(KEYINPUT81), .ZN(n545) );
  NAND2_X1 U637 ( .A1(KEYINPUT80), .A2(n543), .ZN(n544) );
  NAND2_X1 U638 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U639 ( .A1(n546), .A2(KEYINPUT47), .ZN(n547) );
  INV_X1 U640 ( .A(KEYINPUT6), .ZN(n549) );
  INV_X1 U641 ( .A(n550), .ZN(n551) );
  XNOR2_X1 U642 ( .A(n553), .B(KEYINPUT36), .ZN(n554) );
  NAND2_X1 U643 ( .A1(n554), .A2(n698), .ZN(n555) );
  INV_X1 U644 ( .A(n557), .ZN(n558) );
  XNOR2_X2 U645 ( .A(n561), .B(n560), .ZN(n715) );
  INV_X1 U646 ( .A(KEYINPUT38), .ZN(n562) );
  XNOR2_X1 U647 ( .A(n562), .B(n582), .ZN(n711) );
  AND2_X1 U648 ( .A1(n711), .A2(n575), .ZN(n563) );
  NOR2_X1 U649 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U650 ( .A1(n733), .A2(n567), .ZN(n569) );
  XOR2_X1 U651 ( .A(KEYINPUT42), .B(KEYINPUT115), .Z(n568) );
  XNOR2_X1 U652 ( .A(n569), .B(n568), .ZN(n571) );
  XNOR2_X1 U653 ( .A(n571), .B(n570), .ZN(n767) );
  INV_X1 U654 ( .A(n711), .ZN(n713) );
  XNOR2_X1 U655 ( .A(KEYINPUT85), .B(KEYINPUT39), .ZN(n573) );
  XOR2_X1 U656 ( .A(KEYINPUT40), .B(n574), .Z(n769) );
  INV_X1 U657 ( .A(n575), .ZN(n717) );
  NOR2_X1 U658 ( .A1(n717), .A2(n576), .ZN(n577) );
  XNOR2_X1 U659 ( .A(n577), .B(KEYINPUT111), .ZN(n578) );
  NOR2_X1 U660 ( .A1(n578), .A2(n698), .ZN(n579) );
  XNOR2_X1 U661 ( .A(n579), .B(KEYINPUT112), .ZN(n580) );
  XNOR2_X1 U662 ( .A(KEYINPUT43), .B(n580), .ZN(n581) );
  NOR2_X1 U663 ( .A1(n582), .A2(n581), .ZN(n695) );
  NAND2_X1 U664 ( .A1(n583), .A2(n691), .ZN(n694) );
  INV_X1 U665 ( .A(n694), .ZN(n584) );
  INV_X1 U666 ( .A(n587), .ZN(n589) );
  INV_X1 U667 ( .A(G953), .ZN(n588) );
  NOR2_X1 U668 ( .A1(G898), .A2(n588), .ZN(n752) );
  NAND2_X1 U669 ( .A1(n589), .A2(n752), .ZN(n592) );
  INV_X1 U670 ( .A(n590), .ZN(n591) );
  NAND2_X1 U671 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U672 ( .A1(n594), .A2(n593), .ZN(n596) );
  INV_X1 U673 ( .A(KEYINPUT0), .ZN(n595) );
  NAND2_X1 U674 ( .A1(n697), .A2(n599), .ZN(n597) );
  INV_X1 U675 ( .A(n698), .ZN(n615) );
  NOR2_X1 U676 ( .A1(n597), .A2(n615), .ZN(n707) );
  NAND2_X1 U677 ( .A1(n605), .A2(n707), .ZN(n598) );
  XNOR2_X2 U678 ( .A(n598), .B(KEYINPUT31), .ZN(n692) );
  NOR2_X1 U679 ( .A1(n600), .A2(n599), .ZN(n601) );
  AND2_X1 U680 ( .A1(n605), .A2(n601), .ZN(n679) );
  NOR2_X1 U681 ( .A1(n692), .A2(n679), .ZN(n602) );
  NOR2_X1 U682 ( .A1(n712), .A2(n602), .ZN(n603) );
  XNOR2_X1 U683 ( .A(n603), .B(KEYINPUT105), .ZN(n613) );
  XNOR2_X2 U684 ( .A(n604), .B(KEYINPUT33), .ZN(n732) );
  NAND2_X1 U685 ( .A1(n605), .A2(n732), .ZN(n608) );
  XNOR2_X1 U686 ( .A(KEYINPUT77), .B(KEYINPUT34), .ZN(n606) );
  XNOR2_X1 U687 ( .A(n606), .B(KEYINPUT74), .ZN(n607) );
  XNOR2_X1 U688 ( .A(n608), .B(n607), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n609), .A2(n361), .ZN(n610) );
  XNOR2_X2 U690 ( .A(n610), .B(KEYINPUT35), .ZN(n625) );
  NAND2_X1 U691 ( .A1(n625), .A2(KEYINPUT44), .ZN(n611) );
  NAND2_X1 U692 ( .A1(n611), .A2(KEYINPUT87), .ZN(n612) );
  AND2_X1 U693 ( .A1(n613), .A2(n612), .ZN(n616) );
  XOR2_X1 U694 ( .A(n622), .B(KEYINPUT107), .Z(n702) );
  XNOR2_X1 U695 ( .A(n617), .B(KEYINPUT78), .ZN(n618) );
  XNOR2_X1 U696 ( .A(n620), .B(KEYINPUT32), .ZN(n768) );
  AND2_X1 U697 ( .A1(n622), .A2(n700), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n615), .A2(n623), .ZN(n624) );
  NOR2_X1 U699 ( .A1(n621), .A2(n624), .ZN(n682) );
  NOR2_X1 U700 ( .A1(n768), .A2(n682), .ZN(n631) );
  BUF_X2 U701 ( .A(n625), .Z(n635) );
  NAND2_X1 U702 ( .A1(n635), .A2(KEYINPUT67), .ZN(n629) );
  INV_X1 U703 ( .A(n635), .ZN(n627) );
  NOR2_X1 U704 ( .A1(KEYINPUT44), .A2(KEYINPUT67), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n632) );
  OR2_X1 U708 ( .A1(n682), .A2(KEYINPUT67), .ZN(n634) );
  NOR2_X1 U709 ( .A1(n768), .A2(n634), .ZN(n638) );
  INV_X1 U710 ( .A(KEYINPUT87), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n635), .A2(n636), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U713 ( .A1(n639), .A2(KEYINPUT44), .ZN(n640) );
  INV_X1 U714 ( .A(n642), .ZN(n643) );
  NAND2_X1 U715 ( .A1(n643), .A2(KEYINPUT2), .ZN(n644) );
  NAND2_X1 U716 ( .A1(n421), .A2(n744), .ZN(n645) );
  AND2_X2 U717 ( .A1(n646), .A2(n729), .ZN(n665) );
  NAND2_X1 U718 ( .A1(n665), .A2(G472), .ZN(n649) );
  XNOR2_X1 U719 ( .A(n647), .B(KEYINPUT62), .ZN(n648) );
  XNOR2_X1 U720 ( .A(n649), .B(n648), .ZN(n650) );
  INV_X1 U721 ( .A(n650), .ZN(n651) );
  INV_X1 U722 ( .A(n671), .ZN(n743) );
  NAND2_X1 U723 ( .A1(n651), .A2(n671), .ZN(n652) );
  XNOR2_X1 U724 ( .A(n652), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U725 ( .A(n653), .B(G101), .ZN(G3) );
  XOR2_X1 U726 ( .A(n625), .B(G122), .Z(G24) );
  NAND2_X1 U727 ( .A1(n665), .A2(G475), .ZN(n657) );
  XOR2_X1 U728 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n654) );
  XNOR2_X1 U729 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U731 ( .A(n659), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U732 ( .A1(n739), .A2(G469), .ZN(n663) );
  XOR2_X1 U733 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n661) );
  XOR2_X1 U734 ( .A(n661), .B(n660), .Z(n662) );
  XNOR2_X1 U735 ( .A(n663), .B(n662), .ZN(n664) );
  NOR2_X1 U736 ( .A1(n664), .A2(n743), .ZN(G54) );
  NAND2_X1 U737 ( .A1(n665), .A2(G210), .ZN(n670) );
  XOR2_X1 U738 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n667) );
  XNOR2_X1 U739 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U740 ( .A(n670), .B(n669), .ZN(n672) );
  NAND2_X1 U741 ( .A1(n672), .A2(n671), .ZN(n674) );
  XOR2_X1 U742 ( .A(KEYINPUT124), .B(KEYINPUT56), .Z(n673) );
  XNOR2_X1 U743 ( .A(n674), .B(n673), .ZN(G51) );
  NAND2_X1 U744 ( .A1(n679), .A2(n689), .ZN(n675) );
  XNOR2_X1 U745 ( .A(n675), .B(G104), .ZN(G6) );
  XOR2_X1 U746 ( .A(KEYINPUT27), .B(KEYINPUT119), .Z(n677) );
  XNOR2_X1 U747 ( .A(G107), .B(KEYINPUT118), .ZN(n676) );
  XNOR2_X1 U748 ( .A(n677), .B(n676), .ZN(n678) );
  XOR2_X1 U749 ( .A(KEYINPUT26), .B(n678), .Z(n681) );
  NAND2_X1 U750 ( .A1(n679), .A2(n691), .ZN(n680) );
  XNOR2_X1 U751 ( .A(n681), .B(n680), .ZN(G9) );
  XOR2_X1 U752 ( .A(G110), .B(n682), .Z(n683) );
  XNOR2_X1 U753 ( .A(KEYINPUT120), .B(n683), .ZN(G12) );
  XOR2_X1 U754 ( .A(G128), .B(KEYINPUT29), .Z(n685) );
  NAND2_X1 U755 ( .A1(n691), .A2(n686), .ZN(n684) );
  XNOR2_X1 U756 ( .A(n685), .B(n684), .ZN(G30) );
  XOR2_X1 U757 ( .A(G146), .B(KEYINPUT121), .Z(n688) );
  NAND2_X1 U758 ( .A1(n686), .A2(n689), .ZN(n687) );
  XNOR2_X1 U759 ( .A(n688), .B(n687), .ZN(G48) );
  NAND2_X1 U760 ( .A1(n692), .A2(n689), .ZN(n690) );
  XNOR2_X1 U761 ( .A(n690), .B(G113), .ZN(G15) );
  NAND2_X1 U762 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U763 ( .A(n693), .B(G116), .ZN(G18) );
  XNOR2_X1 U764 ( .A(G134), .B(n694), .ZN(G36) );
  XOR2_X1 U765 ( .A(G140), .B(n695), .Z(n696) );
  XNOR2_X1 U766 ( .A(KEYINPUT122), .B(n696), .ZN(G42) );
  NOR2_X1 U767 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U768 ( .A(KEYINPUT50), .B(n699), .Z(n701) );
  NAND2_X1 U769 ( .A1(n701), .A2(n700), .ZN(n706) );
  NAND2_X1 U770 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U771 ( .A(KEYINPUT49), .B(n704), .ZN(n705) );
  NOR2_X1 U772 ( .A1(n706), .A2(n705), .ZN(n708) );
  XNOR2_X1 U773 ( .A(KEYINPUT51), .B(n359), .ZN(n709) );
  NAND2_X1 U774 ( .A1(n709), .A2(n733), .ZN(n710) );
  XNOR2_X1 U775 ( .A(n710), .B(KEYINPUT123), .ZN(n723) );
  AND2_X1 U776 ( .A1(n711), .A2(n715), .ZN(n719) );
  NOR2_X1 U777 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U778 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U779 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U780 ( .A1(n719), .A2(n718), .ZN(n721) );
  INV_X1 U781 ( .A(n732), .ZN(n720) );
  NOR2_X1 U782 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U783 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U784 ( .A(n724), .B(KEYINPUT52), .ZN(n725) );
  NOR2_X1 U785 ( .A1(n726), .A2(n725), .ZN(n731) );
  NAND2_X1 U786 ( .A1(n727), .A2(n388), .ZN(n728) );
  NAND2_X1 U787 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U788 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U789 ( .A(n735), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U790 ( .A1(n739), .A2(G478), .ZN(n737) );
  XNOR2_X1 U791 ( .A(n737), .B(n736), .ZN(n738) );
  NOR2_X1 U792 ( .A1(n743), .A2(n738), .ZN(G63) );
  NAND2_X1 U793 ( .A1(n739), .A2(G217), .ZN(n741) );
  XNOR2_X1 U794 ( .A(n741), .B(n740), .ZN(n742) );
  NOR2_X1 U795 ( .A1(n743), .A2(n742), .ZN(G66) );
  INV_X1 U796 ( .A(n744), .ZN(n745) );
  NOR2_X1 U797 ( .A1(n745), .A2(G953), .ZN(n750) );
  NAND2_X1 U798 ( .A1(G224), .A2(G953), .ZN(n746) );
  XNOR2_X1 U799 ( .A(n746), .B(KEYINPUT126), .ZN(n747) );
  XNOR2_X1 U800 ( .A(KEYINPUT61), .B(n747), .ZN(n748) );
  AND2_X1 U801 ( .A1(n748), .A2(G898), .ZN(n749) );
  NOR2_X1 U802 ( .A1(n750), .A2(n749), .ZN(n754) );
  NOR2_X1 U803 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U804 ( .A(n754), .B(n753), .Z(G69) );
  XOR2_X1 U805 ( .A(n756), .B(n755), .Z(n759) );
  XOR2_X1 U806 ( .A(n759), .B(G227), .Z(n757) );
  NAND2_X1 U807 ( .A1(n757), .A2(G900), .ZN(n758) );
  NAND2_X1 U808 ( .A1(n758), .A2(G953), .ZN(n764) );
  NAND2_X1 U809 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U810 ( .A(KEYINPUT127), .B(n762), .Z(n763) );
  NAND2_X1 U811 ( .A1(n764), .A2(n763), .ZN(G72) );
  XNOR2_X1 U812 ( .A(G125), .B(n765), .ZN(n766) );
  XNOR2_X1 U813 ( .A(n766), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U814 ( .A(G137), .B(n767), .Z(G39) );
  XOR2_X1 U815 ( .A(n768), .B(G119), .Z(G21) );
  XOR2_X1 U816 ( .A(G131), .B(n769), .Z(G33) );
  XOR2_X1 U817 ( .A(G143), .B(n770), .Z(G45) );
endmodule

