//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n566, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n584, new_n585, new_n586, new_n587, new_n589,
    new_n590, new_n591, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n637,
    new_n640, new_n641, new_n643, new_n644, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1199, new_n1200;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT67), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(G2105), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n460), .A2(G101), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND4_X1  g041(.A1(new_n464), .A2(new_n466), .A3(G137), .A4(new_n461), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n469), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n468), .B1(new_n461), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n464), .A2(new_n466), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT68), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n474), .A2(new_n476), .A3(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G124), .ZN(new_n478));
  OR3_X1    g053(.A1(new_n477), .A2(KEYINPUT69), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g054(.A(KEYINPUT69), .B1(new_n477), .B2(new_n478), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n474), .A2(new_n476), .A3(new_n461), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n479), .A2(new_n480), .B1(G136), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(new_n461), .B2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND3_X1  g062(.A1(new_n461), .A2(G102), .A3(G2104), .ZN(new_n488));
  NAND2_X1  g063(.A1(G114), .A2(G2104), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n469), .B2(G126), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n488), .B1(new_n491), .B2(new_n461), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n461), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n469), .A2(KEYINPUT4), .A3(G138), .A4(new_n461), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n492), .A2(new_n497), .ZN(G164));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G543), .ZN(new_n502));
  AND2_X1   g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(G88), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(G50), .A3(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n505), .A2(KEYINPUT70), .A3(new_n506), .ZN(new_n510));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n500), .A2(new_n502), .ZN(new_n512));
  INV_X1    g087(.A(G62), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n509), .A2(new_n510), .B1(G651), .B2(new_n514), .ZN(G166));
  NAND2_X1  g090(.A1(new_n504), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G51), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n500), .B(new_n502), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G89), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n516), .A2(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n512), .A2(KEYINPUT71), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n500), .A2(new_n502), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n527), .A2(G63), .A3(G651), .ZN(new_n528));
  XOR2_X1   g103(.A(KEYINPUT72), .B(KEYINPUT7), .Z(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n523), .A2(new_n528), .A3(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  AND3_X1   g108(.A1(new_n500), .A2(new_n502), .A3(new_n525), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n525), .B1(new_n500), .B2(new_n502), .ZN(new_n535));
  OAI21_X1  g110(.A(G64), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G651), .ZN(new_n539));
  INV_X1    g114(.A(new_n516), .ZN(new_n540));
  XOR2_X1   g115(.A(KEYINPUT73), .B(G52), .Z(new_n541));
  INV_X1    g116(.A(new_n520), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n540), .A2(new_n541), .B1(new_n542), .B2(G90), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n539), .A2(KEYINPUT74), .A3(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n545));
  INV_X1    g120(.A(G651), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n546), .B1(new_n536), .B2(new_n537), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n540), .A2(new_n541), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n542), .A2(G90), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n545), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n544), .A2(new_n551), .ZN(G171));
  XNOR2_X1  g127(.A(KEYINPUT75), .B(G81), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n503), .A2(new_n504), .A3(new_n553), .ZN(new_n554));
  OAI211_X1 g129(.A(G43), .B(G543), .C1(new_n518), .C2(new_n519), .ZN(new_n555));
  AOI21_X1  g130(.A(KEYINPUT76), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  XOR2_X1   g131(.A(KEYINPUT75), .B(G81), .Z(new_n557));
  OAI211_X1 g132(.A(KEYINPUT76), .B(new_n555), .C1(new_n520), .C2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n527), .A2(G56), .ZN(new_n561));
  NAND2_X1  g136(.A1(G68), .A2(G543), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n546), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  AND3_X1   g140(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G36), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n566), .A2(new_n569), .ZN(G188));
  NAND3_X1  g145(.A1(new_n504), .A2(G53), .A3(G543), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(KEYINPUT77), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n573), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n504), .A2(new_n575), .A3(G53), .A4(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n542), .A2(G91), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G65), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n512), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n577), .A2(new_n578), .A3(new_n582), .ZN(G299));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n544), .A2(new_n551), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n584), .B1(new_n544), .B2(new_n551), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G301));
  NAND2_X1  g163(.A1(new_n514), .A2(G651), .ZN(new_n589));
  INV_X1    g164(.A(new_n510), .ZN(new_n590));
  AOI21_X1  g165(.A(KEYINPUT70), .B1(new_n505), .B2(new_n506), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(G303));
  OAI21_X1  g167(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n593));
  INV_X1    g168(.A(G49), .ZN(new_n594));
  INV_X1    g169(.A(G87), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n516), .A2(new_n594), .B1(new_n520), .B2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(G288));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G61), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n512), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G651), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n601), .A2(KEYINPUT79), .A3(G651), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n604), .A2(new_n605), .B1(G86), .B2(new_n542), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n540), .A2(G48), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(G305));
  INV_X1    g183(.A(G47), .ZN(new_n609));
  INV_X1    g184(.A(G85), .ZN(new_n610));
  OAI22_X1  g185(.A1(new_n516), .A2(new_n609), .B1(new_n520), .B2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n527), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(new_n546), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(KEYINPUT80), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n616), .B(new_n612), .C1(new_n613), .C2(new_n546), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n617), .ZN(G290));
  INV_X1    g193(.A(G66), .ZN(new_n619));
  INV_X1    g194(.A(G79), .ZN(new_n620));
  OAI22_X1  g195(.A1(new_n512), .A2(new_n619), .B1(new_n620), .B2(new_n499), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(KEYINPUT81), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT81), .ZN(new_n623));
  OAI221_X1 g198(.A(new_n623), .B1(new_n620), .B2(new_n499), .C1(new_n512), .C2(new_n619), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n622), .A2(G651), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n540), .A2(G54), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n542), .A2(KEYINPUT10), .A3(G92), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n628));
  INV_X1    g203(.A(G92), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n520), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n625), .A2(new_n626), .A3(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(G868), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n587), .B2(new_n633), .ZN(G284));
  OAI21_X1  g210(.A(new_n634), .B1(new_n587), .B2(new_n633), .ZN(G321));
  NAND2_X1  g211(.A1(G299), .A2(new_n633), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(G168), .B2(new_n633), .ZN(G297));
  XNOR2_X1  g213(.A(G297), .B(KEYINPUT82), .ZN(G280));
  INV_X1    g214(.A(new_n632), .ZN(new_n640));
  INV_X1    g215(.A(G559), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(new_n641), .B2(G860), .ZN(G148));
  OAI21_X1  g217(.A(new_n633), .B1(new_n560), .B2(new_n563), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n632), .A2(G559), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n643), .B1(new_n644), .B2(new_n633), .ZN(G323));
  XNOR2_X1  g220(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g221(.A1(new_n460), .A2(new_n462), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(new_n469), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT13), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2100), .ZN(new_n651));
  INV_X1    g226(.A(new_n477), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(G123), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n482), .A2(G135), .ZN(new_n654));
  NOR2_X1   g229(.A1(G99), .A2(G2105), .ZN(new_n655));
  OAI21_X1  g230(.A(G2104), .B1(new_n461), .B2(G111), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n653), .B(new_n654), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2096), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT83), .Z(G156));
  XNOR2_X1  g235(.A(KEYINPUT15), .B(G2435), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2438), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2427), .B(G2430), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT86), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n662), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(KEYINPUT14), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2451), .B(G2454), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2443), .B(G2446), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT85), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT84), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT16), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n668), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1341), .B(G1348), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(G14), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G401));
  XOR2_X1   g252(.A(G2067), .B(G2678), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT88), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2072), .B(G2078), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2084), .B(G2090), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT87), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n680), .B(KEYINPUT17), .Z(new_n685));
  OAI211_X1 g260(.A(new_n682), .B(new_n684), .C1(new_n679), .C2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT90), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n679), .A2(new_n684), .A3(new_n681), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n684), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n692), .A2(new_n685), .A3(new_n679), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n688), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G2096), .B(G2100), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(G227));
  INV_X1    g271(.A(KEYINPUT20), .ZN(new_n697));
  XOR2_X1   g272(.A(G1961), .B(G1966), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT91), .ZN(new_n699));
  XOR2_X1   g274(.A(G1956), .B(G2474), .Z(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1971), .B(G1976), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT19), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n697), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n699), .A2(new_n700), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n706), .A2(new_n703), .A3(new_n701), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n701), .A2(new_n697), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(new_n705), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n704), .B(new_n707), .C1(new_n709), .C2(new_n703), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G1996), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT92), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1991), .ZN(new_n714));
  XOR2_X1   g289(.A(G1981), .B(G1986), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT93), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n714), .B(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n711), .B(new_n717), .ZN(G229));
  NAND2_X1  g293(.A1(G168), .A2(G16), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G16), .B2(G21), .ZN(new_n720));
  INV_X1    g295(.A(G1966), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT104), .ZN(new_n723));
  INV_X1    g298(.A(G26), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n724), .A2(G29), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n652), .A2(G128), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n482), .A2(G140), .ZN(new_n727));
  OR2_X1    g302(.A1(G104), .A2(G2105), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n728), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n725), .B1(new_n730), .B2(G29), .ZN(new_n731));
  MUX2_X1   g306(.A(new_n725), .B(new_n731), .S(KEYINPUT28), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G2067), .ZN(new_n733));
  NOR2_X1   g308(.A1(G4), .A2(G16), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n640), .B2(G16), .ZN(new_n735));
  INV_X1    g310(.A(G1348), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n482), .A2(G141), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n652), .A2(G129), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT26), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n647), .A2(G105), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n738), .A2(new_n739), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G29), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G29), .B2(G32), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT27), .B(G1996), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n733), .B(new_n737), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  AND2_X1   g323(.A1(KEYINPUT96), .A2(G16), .ZN(new_n749));
  NOR2_X1   g324(.A1(KEYINPUT96), .A2(G16), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n564), .A2(new_n752), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n752), .A2(G19), .ZN(new_n754));
  OAI21_X1  g329(.A(KEYINPUT98), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(KEYINPUT98), .B2(new_n754), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1341), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n746), .A2(new_n747), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT103), .ZN(new_n759));
  NOR3_X1   g334(.A1(new_n748), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT99), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G29), .B2(G33), .ZN(new_n762));
  OR3_X1    g337(.A1(new_n761), .A2(G29), .A3(G33), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n482), .A2(G139), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT100), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT101), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G2105), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT25), .Z(new_n770));
  NAND3_X1  g345(.A1(new_n765), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(G29), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n762), .B(new_n763), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G2072), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT102), .Z(new_n776));
  NAND2_X1  g351(.A1(new_n772), .A2(G35), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G162), .B2(new_n772), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT105), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT29), .B(G2090), .Z(new_n780));
  XOR2_X1   g355(.A(new_n779), .B(new_n780), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n772), .A2(G27), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G164), .B2(new_n772), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(G2078), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(G2078), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n784), .B(new_n785), .C1(new_n720), .C2(new_n721), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n752), .A2(KEYINPUT23), .A3(G20), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT23), .ZN(new_n788));
  INV_X1    g363(.A(G20), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n751), .B2(new_n789), .ZN(new_n790));
  AND3_X1   g365(.A1(new_n577), .A2(new_n578), .A3(new_n582), .ZN(new_n791));
  INV_X1    g366(.A(G16), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n787), .B(new_n790), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1956), .ZN(new_n794));
  OR2_X1    g369(.A1(KEYINPUT24), .A2(G34), .ZN(new_n795));
  NAND2_X1  g370(.A1(KEYINPUT24), .A2(G34), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n795), .A2(new_n772), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G160), .B2(new_n772), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2084), .ZN(new_n799));
  INV_X1    g374(.A(G28), .ZN(new_n800));
  AOI21_X1  g375(.A(G29), .B1(new_n800), .B2(KEYINPUT30), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(KEYINPUT30), .B2(new_n800), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n657), .B2(new_n772), .ZN(new_n803));
  OR4_X1    g378(.A1(new_n786), .A2(new_n794), .A3(new_n799), .A4(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(G5), .A2(G16), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G171), .B2(G16), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1961), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n773), .A2(new_n774), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT31), .B(G11), .Z(new_n809));
  NOR4_X1   g384(.A1(new_n804), .A2(new_n807), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n760), .A2(new_n776), .A3(new_n781), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n752), .A2(G22), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G166), .B2(new_n752), .ZN(new_n813));
  MUX2_X1   g388(.A(new_n812), .B(new_n813), .S(KEYINPUT97), .Z(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(G1971), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n792), .A2(G6), .ZN(new_n816));
  INV_X1    g391(.A(G305), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(new_n792), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT32), .B(G1981), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n792), .A2(G23), .ZN(new_n821));
  INV_X1    g396(.A(G288), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n822), .B2(new_n792), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT33), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G1976), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n815), .A2(new_n820), .A3(new_n825), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n826), .A2(KEYINPUT34), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n772), .A2(G25), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n652), .A2(G119), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n482), .A2(G131), .ZN(new_n830));
  OR3_X1    g405(.A1(KEYINPUT95), .A2(G95), .A3(G2105), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n461), .A2(G107), .ZN(new_n832));
  OAI21_X1  g407(.A(KEYINPUT95), .B1(G95), .B2(G2105), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n831), .A2(new_n832), .A3(G2104), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n829), .A2(new_n830), .A3(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n828), .B1(new_n836), .B2(new_n772), .ZN(new_n837));
  MUX2_X1   g412(.A(new_n828), .B(new_n837), .S(KEYINPUT94), .Z(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT35), .B(G1991), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n826), .A2(KEYINPUT34), .ZN(new_n841));
  MUX2_X1   g416(.A(G24), .B(G290), .S(new_n751), .Z(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(G1986), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n842), .A2(G1986), .ZN(new_n844));
  AOI211_X1 g419(.A(new_n843), .B(new_n844), .C1(new_n839), .C2(new_n838), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n827), .A2(new_n840), .A3(new_n841), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT36), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n841), .A2(new_n845), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT36), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n848), .A2(new_n849), .A3(new_n840), .A4(new_n827), .ZN(new_n850));
  AOI211_X1 g425(.A(new_n723), .B(new_n811), .C1(new_n847), .C2(new_n850), .ZN(G311));
  AOI21_X1  g426(.A(new_n811), .B1(new_n847), .B2(new_n850), .ZN(new_n852));
  INV_X1    g427(.A(new_n723), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(G150));
  INV_X1    g429(.A(G55), .ZN(new_n855));
  INV_X1    g430(.A(G93), .ZN(new_n856));
  OAI22_X1  g431(.A1(new_n516), .A2(new_n855), .B1(new_n520), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n527), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n858), .B1(new_n859), .B2(new_n546), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(G860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT107), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT37), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n632), .A2(new_n641), .ZN(new_n864));
  XNOR2_X1  g439(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT106), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n560), .B2(new_n563), .ZN(new_n868));
  INV_X1    g443(.A(G56), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(new_n524), .B2(new_n526), .ZN(new_n870));
  INV_X1    g445(.A(new_n562), .ZN(new_n871));
  OAI21_X1  g446(.A(G651), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n872), .B(KEYINPUT106), .C1(new_n556), .C2(new_n559), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n868), .A2(new_n873), .A3(new_n860), .ZN(new_n874));
  INV_X1    g449(.A(new_n860), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n564), .A2(new_n875), .A3(KEYINPUT106), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n866), .B(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n863), .B1(new_n878), .B2(G860), .ZN(G145));
  XNOR2_X1  g454(.A(new_n657), .B(G160), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(G162), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n744), .A2(new_n730), .ZN(new_n882));
  INV_X1    g457(.A(new_n730), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n883), .A2(new_n743), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT108), .ZN(new_n885));
  NOR2_X1   g460(.A1(G164), .A2(new_n885), .ZN(new_n886));
  NOR3_X1   g461(.A1(new_n492), .A2(new_n497), .A3(KEYINPUT108), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n882), .A2(new_n884), .A3(new_n888), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n886), .A2(new_n887), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n744), .A2(new_n730), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n883), .A2(new_n743), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n771), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G142), .ZN(new_n895));
  NOR2_X1   g470(.A1(G106), .A2(G2105), .ZN(new_n896));
  OAI21_X1  g471(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n897));
  OAI22_X1  g472(.A1(new_n481), .A2(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n898), .B1(G130), .B2(new_n652), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(new_n649), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n835), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n888), .B1(new_n882), .B2(new_n884), .ZN(new_n902));
  INV_X1    g477(.A(new_n771), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n891), .A2(new_n892), .A3(new_n890), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n894), .A2(new_n901), .A3(KEYINPUT109), .A4(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n900), .B(new_n836), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n889), .A2(new_n893), .A3(new_n771), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n903), .B1(new_n902), .B2(new_n904), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n894), .A2(new_n901), .A3(new_n905), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n881), .B(new_n906), .C1(new_n912), .C2(KEYINPUT109), .ZN(new_n913));
  INV_X1    g488(.A(G37), .ZN(new_n914));
  INV_X1    g489(.A(new_n881), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n910), .A2(new_n911), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g493(.A1(new_n860), .A2(new_n633), .ZN(new_n919));
  NAND2_X1  g494(.A1(G166), .A2(G288), .ZN(new_n920));
  NAND2_X1  g495(.A1(G303), .A2(new_n822), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n817), .ZN(new_n923));
  NAND2_X1  g498(.A1(G290), .A2(KEYINPUT112), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT112), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n615), .A2(new_n925), .A3(new_n617), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n920), .A2(new_n921), .A3(G305), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n923), .A2(new_n924), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n920), .A2(new_n921), .A3(G305), .ZN(new_n929));
  AOI21_X1  g504(.A(G305), .B1(new_n920), .B2(new_n921), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n615), .A2(new_n925), .A3(new_n617), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n925), .B1(new_n615), .B2(new_n617), .ZN(new_n932));
  OAI22_X1  g507(.A1(new_n929), .A2(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n928), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT42), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n877), .B(new_n644), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n632), .A2(new_n791), .ZN(new_n937));
  NAND4_X1  g512(.A1(G299), .A2(new_n626), .A3(new_n625), .A4(new_n631), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n640), .A2(KEYINPUT110), .A3(G299), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n936), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(KEYINPUT41), .ZN(new_n944));
  AOI211_X1 g519(.A(KEYINPUT111), .B(KEYINPUT41), .C1(new_n937), .C2(new_n938), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n937), .A2(new_n938), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT41), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT111), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n944), .A2(new_n946), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n943), .B1(new_n936), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n935), .B(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n919), .B1(new_n953), .B2(new_n633), .ZN(G295));
  OAI21_X1  g529(.A(new_n919), .B1(new_n953), .B2(new_n633), .ZN(G331));
  INV_X1    g530(.A(new_n934), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n874), .A2(new_n876), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT74), .B1(new_n539), .B2(new_n543), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n547), .A2(new_n550), .A3(new_n545), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT78), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n544), .A2(new_n551), .A3(new_n584), .ZN(new_n961));
  AOI21_X1  g536(.A(G286), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(G171), .A2(G286), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n957), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(G168), .B1(new_n585), .B2(new_n586), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n966), .A2(new_n963), .A3(new_n877), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n951), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n965), .A2(new_n942), .A3(new_n967), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n956), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT114), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n948), .B1(new_n940), .B2(new_n941), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n974), .B1(new_n947), .B2(new_n948), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n973), .A2(new_n975), .A3(new_n945), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n966), .A2(new_n963), .A3(new_n877), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n877), .B1(new_n966), .B2(new_n963), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n965), .A2(new_n942), .A3(new_n967), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n981), .A2(KEYINPUT114), .A3(new_n956), .ZN(new_n982));
  AOI21_X1  g557(.A(G37), .B1(new_n972), .B2(new_n982), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n928), .A2(new_n933), .A3(KEYINPUT113), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT113), .B1(new_n928), .B2(new_n933), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n986), .A2(new_n980), .A3(new_n979), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT43), .B1(new_n983), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n948), .B1(new_n965), .B2(new_n967), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n947), .ZN(new_n990));
  INV_X1    g565(.A(new_n942), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n986), .B(new_n990), .C1(new_n991), .C2(new_n989), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT114), .B1(new_n981), .B2(new_n956), .ZN(new_n993));
  AOI211_X1 g568(.A(new_n971), .B(new_n934), .C1(new_n979), .C2(new_n980), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n914), .B(new_n992), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT43), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT44), .B1(new_n988), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n996), .B1(new_n983), .B2(new_n987), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n995), .A2(KEYINPUT43), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n998), .A2(new_n1002), .ZN(G397));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n468), .B(G40), .C1(new_n461), .C2(new_n470), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1004), .B(new_n1006), .C1(new_n888), .C2(G1384), .ZN(new_n1007));
  INV_X1    g582(.A(G1996), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1007), .A2(new_n1008), .A3(new_n744), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1007), .A2(G1996), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n1011), .A2(new_n1012), .B1(new_n744), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1007), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n730), .B(G2067), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT116), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n835), .A2(new_n839), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1019), .B(KEYINPUT126), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1014), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G2067), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n883), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1007), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n1013), .A2(KEYINPUT46), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1015), .B1(new_n743), .B2(new_n1016), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1013), .A2(KEYINPUT46), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  XOR2_X1   g603(.A(new_n1028), .B(KEYINPUT47), .Z(new_n1029));
  AND2_X1   g604(.A1(new_n835), .A2(new_n839), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1015), .B1(new_n1019), .B2(new_n1030), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1007), .A2(G1986), .A3(G290), .ZN(new_n1032));
  XOR2_X1   g607(.A(new_n1032), .B(KEYINPUT48), .Z(new_n1033));
  AND4_X1   g608(.A1(new_n1031), .A2(new_n1014), .A3(new_n1018), .A4(new_n1033), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n1024), .A2(new_n1029), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1384), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(new_n492), .B2(new_n497), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1037), .A2(new_n1005), .ZN(new_n1038));
  INV_X1    g613(.A(G8), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT49), .ZN(new_n1041));
  INV_X1    g616(.A(G1981), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n606), .A2(new_n1042), .A3(new_n607), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1042), .B1(new_n606), .B2(new_n607), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1041), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1045), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1047), .A2(KEYINPUT49), .A3(new_n1043), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1046), .A2(new_n1048), .A3(new_n1040), .ZN(new_n1049));
  INV_X1    g624(.A(G1976), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1049), .A2(new_n1050), .A3(new_n822), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1040), .B1(new_n1051), .B2(new_n1044), .ZN(new_n1052));
  NOR2_X1   g627(.A1(G166), .A2(new_n1039), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT55), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1053), .A2(KEYINPUT55), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1053), .A2(KEYINPUT118), .A3(KEYINPUT55), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  OAI211_X1 g634(.A(KEYINPUT45), .B(new_n1036), .C1(new_n886), .C2(new_n887), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1005), .B1(new_n1037), .B2(new_n1004), .ZN(new_n1061));
  AOI21_X1  g636(.A(G1971), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1037), .A2(KEYINPUT50), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT50), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1064), .B(new_n1036), .C1(new_n492), .C2(new_n497), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1063), .A2(new_n1006), .A3(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT117), .B(G2090), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1059), .B(G8), .C1(new_n1062), .C2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1040), .B1(new_n1050), .B2(G288), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT52), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT52), .B1(G288), .B2(new_n1050), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1040), .B(new_n1073), .C1(new_n1050), .C2(G288), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1049), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1070), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(G8), .B1(new_n1062), .B2(new_n1068), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1077), .A2(new_n1057), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n495), .A2(new_n496), .ZN(new_n1079));
  INV_X1    g654(.A(new_n488), .ZN(new_n1080));
  INV_X1    g655(.A(G126), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n489), .B1(new_n473), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1080), .B1(new_n1082), .B2(G2105), .ZN(new_n1083));
  AOI21_X1  g658(.A(G1384), .B1(new_n1079), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1006), .B1(new_n1084), .B2(KEYINPUT45), .ZN(new_n1085));
  OAI211_X1 g660(.A(KEYINPUT45), .B(new_n1036), .C1(new_n492), .C2(new_n497), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n721), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT119), .B(G2084), .Z(new_n1089));
  NAND4_X1  g664(.A1(new_n1063), .A2(new_n1006), .A3(new_n1065), .A4(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1039), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1091), .A2(G168), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1075), .A2(new_n1078), .A3(new_n1069), .A4(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT63), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1093), .A2(KEYINPUT120), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1094), .B1(new_n1093), .B2(KEYINPUT120), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1052), .B(new_n1076), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n1098));
  AND4_X1   g673(.A1(new_n1006), .A2(new_n1063), .A3(new_n1065), .A4(new_n1089), .ZN(new_n1099));
  AOI21_X1  g674(.A(G1966), .B1(new_n1061), .B2(new_n1086), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1088), .A2(KEYINPUT122), .A3(new_n1090), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1101), .A2(G168), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT51), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1104), .A2(new_n1039), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1103), .A2(KEYINPUT124), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT124), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1104), .B1(G168), .B2(new_n1039), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1108), .B1(new_n1091), .B2(G168), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1106), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1111));
  NOR2_X1   g686(.A1(G168), .A2(new_n1039), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT123), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1111), .A2(new_n1115), .A3(new_n1112), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT62), .B1(new_n1110), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1119), .B1(new_n1120), .B2(G2078), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1066), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1122), .A2(G1961), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1119), .A2(G2078), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1061), .A2(new_n1124), .A3(new_n1086), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1121), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n587), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1109), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1103), .A2(KEYINPUT124), .A3(new_n1105), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1129), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1118), .A2(new_n1128), .A3(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1060), .A2(new_n1008), .A3(new_n1061), .ZN(new_n1139));
  XOR2_X1   g714(.A(KEYINPUT58), .B(G1341), .Z(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n1037), .B2(new_n1005), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n564), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT59), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1142), .A2(new_n1145), .A3(new_n564), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1066), .A2(new_n736), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1038), .A2(new_n1022), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1150), .A2(new_n1151), .A3(new_n640), .ZN(new_n1152));
  XNOR2_X1  g727(.A(KEYINPUT56), .B(G2072), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1060), .A2(new_n1061), .A3(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n791), .B(KEYINPUT57), .ZN(new_n1155));
  INV_X1    g730(.A(G1956), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1066), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1154), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT121), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1152), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1158), .A2(KEYINPUT61), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n632), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1164), .B1(new_n1151), .B2(new_n1150), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1147), .A2(new_n1162), .A3(new_n1163), .A4(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1158), .A2(new_n640), .A3(new_n1150), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n1168), .A2(new_n1155), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1166), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1129), .A2(new_n1135), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1004), .B1(new_n888), .B2(G1384), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1172), .A2(new_n1006), .A3(new_n1060), .A4(new_n1124), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1121), .A2(new_n1173), .A3(new_n1123), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1127), .B1(new_n1174), .B2(new_n587), .ZN(new_n1175));
  XOR2_X1   g750(.A(KEYINPUT125), .B(KEYINPUT54), .Z(new_n1176));
  NAND4_X1  g751(.A1(new_n1121), .A2(G301), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n1177), .A2(KEYINPUT54), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1174), .A2(G171), .ZN(new_n1179));
  AOI22_X1  g754(.A1(new_n1175), .A2(new_n1176), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1170), .A2(new_n1171), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1138), .A2(new_n1181), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1075), .A2(new_n1078), .A3(new_n1069), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1097), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g759(.A(G290), .B(G1986), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(new_n1015), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1014), .A2(new_n1031), .A3(new_n1018), .A4(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1035), .B1(new_n1184), .B2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g763(.A1(G401), .A2(G229), .ZN(new_n1190));
  INV_X1    g764(.A(G319), .ZN(new_n1191));
  NOR2_X1   g765(.A1(G227), .A2(new_n1191), .ZN(new_n1192));
  XOR2_X1   g766(.A(new_n1192), .B(KEYINPUT127), .Z(new_n1193));
  NAND2_X1  g767(.A1(new_n917), .A2(new_n1193), .ZN(new_n1194));
  OAI211_X1 g768(.A(new_n914), .B(new_n987), .C1(new_n993), .C2(new_n994), .ZN(new_n1195));
  NAND2_X1  g769(.A1(new_n1195), .A2(KEYINPUT43), .ZN(new_n1196));
  NAND3_X1  g770(.A1(new_n983), .A2(new_n996), .A3(new_n992), .ZN(new_n1197));
  AOI211_X1 g771(.A(new_n1190), .B(new_n1194), .C1(new_n1196), .C2(new_n1197), .ZN(G308));
  AOI21_X1  g772(.A(new_n1194), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1199));
  INV_X1    g773(.A(new_n1190), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n1199), .A2(new_n1200), .ZN(G225));
endmodule


