

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U551 ( .A1(G2105), .A2(G2104), .ZN(n894) );
  XNOR2_X2 U552 ( .A(n672), .B(KEYINPUT32), .ZN(n696) );
  NAND2_X1 U553 ( .A1(n734), .A2(n736), .ZN(n663) );
  OR2_X1 U554 ( .A1(n525), .A2(n524), .ZN(n532) );
  BUF_X1 U555 ( .A(n713), .Z(n714) );
  AND2_X2 U556 ( .A1(n521), .A2(G2104), .ZN(n890) );
  NOR2_X1 U557 ( .A1(G2104), .A2(n521), .ZN(n713) );
  NOR2_X2 U558 ( .A1(n532), .A2(n531), .ZN(G160) );
  NOR2_X1 U559 ( .A1(n1006), .A2(n622), .ZN(n628) );
  XNOR2_X1 U560 ( .A(n642), .B(n641), .ZN(n649) );
  AND2_X1 U561 ( .A1(G160), .A2(G40), .ZN(n734) );
  NOR2_X1 U562 ( .A1(G164), .A2(G1384), .ZN(n736) );
  XOR2_X1 U563 ( .A(n673), .B(KEYINPUT104), .Z(n519) );
  NOR2_X1 U564 ( .A1(n682), .A2(n681), .ZN(n520) );
  NOR2_X1 U565 ( .A1(n663), .A2(n954), .ZN(n619) );
  INV_X1 U566 ( .A(KEYINPUT103), .ZN(n651) );
  INV_X1 U567 ( .A(KEYINPUT29), .ZN(n641) );
  INV_X1 U568 ( .A(KEYINPUT31), .ZN(n659) );
  INV_X1 U569 ( .A(KEYINPUT105), .ZN(n669) );
  XNOR2_X1 U570 ( .A(n670), .B(n669), .ZN(n671) );
  NAND2_X1 U571 ( .A1(n671), .A2(G8), .ZN(n672) );
  INV_X1 U572 ( .A(KEYINPUT107), .ZN(n693) );
  INV_X1 U573 ( .A(KEYINPUT12), .ZN(n602) );
  XNOR2_X1 U574 ( .A(n603), .B(n602), .ZN(n604) );
  INV_X1 U575 ( .A(KEYINPUT109), .ZN(n710) );
  INV_X1 U576 ( .A(KEYINPUT77), .ZN(n596) );
  XNOR2_X1 U577 ( .A(n597), .B(n596), .ZN(n598) );
  NOR2_X1 U578 ( .A1(G651), .A2(G543), .ZN(n798) );
  XOR2_X1 U579 ( .A(KEYINPUT15), .B(n600), .Z(n1022) );
  NOR2_X2 U580 ( .A1(G651), .A2(n570), .ZN(n799) );
  INV_X1 U581 ( .A(G2105), .ZN(n521) );
  NAND2_X1 U582 ( .A1(G125), .A2(n713), .ZN(n522) );
  XOR2_X1 U583 ( .A(n522), .B(KEYINPUT64), .Z(n525) );
  NAND2_X1 U584 ( .A1(G101), .A2(n890), .ZN(n523) );
  XNOR2_X1 U585 ( .A(KEYINPUT23), .B(n523), .ZN(n524) );
  NOR2_X1 U586 ( .A1(G2105), .A2(G2104), .ZN(n526) );
  XOR2_X1 U587 ( .A(KEYINPUT66), .B(n526), .Z(n527) );
  XNOR2_X1 U588 ( .A(KEYINPUT17), .B(n527), .ZN(n717) );
  NAND2_X1 U589 ( .A1(G137), .A2(n717), .ZN(n530) );
  NAND2_X1 U590 ( .A1(G113), .A2(n894), .ZN(n528) );
  XOR2_X1 U591 ( .A(KEYINPUT65), .B(n528), .Z(n529) );
  NAND2_X1 U592 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U593 ( .A1(G91), .A2(n798), .ZN(n534) );
  XOR2_X1 U594 ( .A(KEYINPUT0), .B(G543), .Z(n570) );
  XNOR2_X1 U595 ( .A(KEYINPUT67), .B(G651), .ZN(n535) );
  NOR2_X1 U596 ( .A1(n570), .A2(n535), .ZN(n804) );
  NAND2_X1 U597 ( .A1(G78), .A2(n804), .ZN(n533) );
  NAND2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n539) );
  NOR2_X1 U599 ( .A1(G543), .A2(n535), .ZN(n536) );
  XOR2_X1 U600 ( .A(KEYINPUT1), .B(n536), .Z(n802) );
  NAND2_X1 U601 ( .A1(G65), .A2(n802), .ZN(n537) );
  XNOR2_X1 U602 ( .A(KEYINPUT71), .B(n537), .ZN(n538) );
  NOR2_X1 U603 ( .A1(n539), .A2(n538), .ZN(n541) );
  NAND2_X1 U604 ( .A1(n799), .A2(G53), .ZN(n540) );
  NAND2_X1 U605 ( .A1(n541), .A2(n540), .ZN(G299) );
  NAND2_X1 U606 ( .A1(n799), .A2(G52), .ZN(n543) );
  NAND2_X1 U607 ( .A1(G64), .A2(n802), .ZN(n542) );
  NAND2_X1 U608 ( .A1(n543), .A2(n542), .ZN(n549) );
  NAND2_X1 U609 ( .A1(n798), .A2(G90), .ZN(n544) );
  XOR2_X1 U610 ( .A(KEYINPUT69), .B(n544), .Z(n546) );
  NAND2_X1 U611 ( .A1(G77), .A2(n804), .ZN(n545) );
  NAND2_X1 U612 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U613 ( .A(KEYINPUT9), .B(n547), .Z(n548) );
  NOR2_X1 U614 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U615 ( .A(KEYINPUT70), .B(n550), .ZN(G171) );
  NAND2_X1 U616 ( .A1(n798), .A2(G89), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n551), .B(KEYINPUT4), .ZN(n553) );
  NAND2_X1 U618 ( .A1(G76), .A2(n804), .ZN(n552) );
  NAND2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n554), .B(KEYINPUT5), .ZN(n561) );
  XNOR2_X1 U621 ( .A(KEYINPUT79), .B(KEYINPUT6), .ZN(n559) );
  NAND2_X1 U622 ( .A1(G63), .A2(n802), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n555), .B(KEYINPUT78), .ZN(n557) );
  NAND2_X1 U624 ( .A1(G51), .A2(n799), .ZN(n556) );
  NAND2_X1 U625 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n560) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(KEYINPUT7), .B(n562), .ZN(G168) );
  XOR2_X1 U629 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U630 ( .A1(n798), .A2(G88), .ZN(n564) );
  NAND2_X1 U631 ( .A1(G62), .A2(n802), .ZN(n563) );
  NAND2_X1 U632 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n799), .A2(G50), .ZN(n566) );
  NAND2_X1 U634 ( .A1(G75), .A2(n804), .ZN(n565) );
  NAND2_X1 U635 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U636 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U637 ( .A(KEYINPUT84), .B(n569), .Z(G303) );
  NAND2_X1 U638 ( .A1(G87), .A2(n570), .ZN(n572) );
  NAND2_X1 U639 ( .A1(G74), .A2(G651), .ZN(n571) );
  NAND2_X1 U640 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U641 ( .A1(n802), .A2(n573), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n799), .A2(G49), .ZN(n574) );
  NAND2_X1 U643 ( .A1(n575), .A2(n574), .ZN(G288) );
  NAND2_X1 U644 ( .A1(n804), .A2(G73), .ZN(n576) );
  XOR2_X1 U645 ( .A(KEYINPUT2), .B(n576), .Z(n581) );
  NAND2_X1 U646 ( .A1(n798), .A2(G86), .ZN(n578) );
  NAND2_X1 U647 ( .A1(G61), .A2(n802), .ZN(n577) );
  NAND2_X1 U648 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U649 ( .A(KEYINPUT83), .B(n579), .Z(n580) );
  NOR2_X1 U650 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U651 ( .A1(n799), .A2(G48), .ZN(n582) );
  NAND2_X1 U652 ( .A1(n583), .A2(n582), .ZN(G305) );
  NAND2_X1 U653 ( .A1(n798), .A2(G85), .ZN(n585) );
  NAND2_X1 U654 ( .A1(G60), .A2(n802), .ZN(n584) );
  NAND2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n799), .A2(G47), .ZN(n586) );
  XOR2_X1 U657 ( .A(KEYINPUT68), .B(n586), .Z(n587) );
  NOR2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n590) );
  NAND2_X1 U659 ( .A1(G72), .A2(n804), .ZN(n589) );
  NAND2_X1 U660 ( .A1(n590), .A2(n589), .ZN(G290) );
  NAND2_X1 U661 ( .A1(n798), .A2(G92), .ZN(n592) );
  NAND2_X1 U662 ( .A1(G66), .A2(n802), .ZN(n591) );
  NAND2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n599) );
  NAND2_X1 U664 ( .A1(n799), .A2(G54), .ZN(n593) );
  XNOR2_X1 U665 ( .A(n593), .B(KEYINPUT76), .ZN(n595) );
  NAND2_X1 U666 ( .A1(G79), .A2(n804), .ZN(n594) );
  NAND2_X1 U667 ( .A1(n595), .A2(n594), .ZN(n597) );
  NOR2_X1 U668 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U669 ( .A1(n802), .A2(G56), .ZN(n601) );
  XOR2_X1 U670 ( .A(KEYINPUT14), .B(n601), .Z(n609) );
  NAND2_X1 U671 ( .A1(G81), .A2(n798), .ZN(n603) );
  XNOR2_X1 U672 ( .A(n604), .B(KEYINPUT75), .ZN(n606) );
  NAND2_X1 U673 ( .A1(G68), .A2(n804), .ZN(n605) );
  NAND2_X1 U674 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U675 ( .A(KEYINPUT13), .B(n607), .Z(n608) );
  NOR2_X1 U676 ( .A1(n609), .A2(n608), .ZN(n611) );
  NAND2_X1 U677 ( .A1(n799), .A2(G43), .ZN(n610) );
  NAND2_X1 U678 ( .A1(n611), .A2(n610), .ZN(n1006) );
  NAND2_X1 U679 ( .A1(G102), .A2(n890), .ZN(n613) );
  NAND2_X1 U680 ( .A1(G114), .A2(n894), .ZN(n612) );
  AND2_X1 U681 ( .A1(n613), .A2(n612), .ZN(n616) );
  NAND2_X1 U682 ( .A1(G126), .A2(n713), .ZN(n614) );
  XOR2_X1 U683 ( .A(KEYINPUT89), .B(n614), .Z(n615) );
  AND2_X1 U684 ( .A1(n616), .A2(n615), .ZN(n618) );
  NAND2_X1 U685 ( .A1(n717), .A2(G138), .ZN(n617) );
  AND2_X1 U686 ( .A1(n618), .A2(n617), .ZN(G164) );
  INV_X1 U687 ( .A(G1996), .ZN(n954) );
  XOR2_X1 U688 ( .A(n619), .B(KEYINPUT26), .Z(n621) );
  NAND2_X1 U689 ( .A1(n663), .A2(G1341), .ZN(n620) );
  NAND2_X1 U690 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U691 ( .A1(n1022), .A2(n628), .ZN(n627) );
  AND2_X1 U692 ( .A1(n736), .A2(n734), .ZN(n644) );
  AND2_X1 U693 ( .A1(n644), .A2(G2067), .ZN(n623) );
  XOR2_X1 U694 ( .A(n623), .B(KEYINPUT102), .Z(n625) );
  NAND2_X1 U695 ( .A1(n663), .A2(G1348), .ZN(n624) );
  NAND2_X1 U696 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n627), .A2(n626), .ZN(n630) );
  OR2_X1 U698 ( .A1(n1022), .A2(n628), .ZN(n629) );
  NAND2_X1 U699 ( .A1(n630), .A2(n629), .ZN(n635) );
  INV_X1 U700 ( .A(G299), .ZN(n1012) );
  NAND2_X1 U701 ( .A1(n644), .A2(G2072), .ZN(n631) );
  XNOR2_X1 U702 ( .A(n631), .B(KEYINPUT27), .ZN(n633) );
  INV_X1 U703 ( .A(G1956), .ZN(n926) );
  NOR2_X1 U704 ( .A1(n926), .A2(n644), .ZN(n632) );
  NOR2_X1 U705 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U706 ( .A1(n1012), .A2(n636), .ZN(n634) );
  NAND2_X1 U707 ( .A1(n635), .A2(n634), .ZN(n640) );
  NOR2_X1 U708 ( .A1(n1012), .A2(n636), .ZN(n638) );
  XNOR2_X1 U709 ( .A(KEYINPUT101), .B(KEYINPUT28), .ZN(n637) );
  XNOR2_X1 U710 ( .A(n638), .B(n637), .ZN(n639) );
  NAND2_X1 U711 ( .A1(n640), .A2(n639), .ZN(n642) );
  NOR2_X1 U712 ( .A1(n644), .A2(G1961), .ZN(n643) );
  XNOR2_X1 U713 ( .A(n643), .B(KEYINPUT99), .ZN(n646) );
  XNOR2_X1 U714 ( .A(KEYINPUT25), .B(G2078), .ZN(n953) );
  NAND2_X1 U715 ( .A1(n644), .A2(n953), .ZN(n645) );
  NAND2_X1 U716 ( .A1(n646), .A2(n645), .ZN(n656) );
  NAND2_X1 U717 ( .A1(G171), .A2(n656), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n647), .B(KEYINPUT100), .ZN(n648) );
  NAND2_X1 U719 ( .A1(n649), .A2(n648), .ZN(n662) );
  NAND2_X1 U720 ( .A1(G8), .A2(n663), .ZN(n707) );
  NOR2_X1 U721 ( .A1(G1966), .A2(n707), .ZN(n674) );
  NOR2_X1 U722 ( .A1(n663), .A2(G2084), .ZN(n650) );
  XNOR2_X1 U723 ( .A(n650), .B(KEYINPUT98), .ZN(n675) );
  NOR2_X1 U724 ( .A1(n674), .A2(n675), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n652), .B(n651), .ZN(n653) );
  NAND2_X1 U726 ( .A1(n653), .A2(G8), .ZN(n654) );
  XNOR2_X1 U727 ( .A(n654), .B(KEYINPUT30), .ZN(n655) );
  NOR2_X1 U728 ( .A1(G168), .A2(n655), .ZN(n658) );
  NOR2_X1 U729 ( .A1(G171), .A2(n656), .ZN(n657) );
  NOR2_X1 U730 ( .A1(n658), .A2(n657), .ZN(n660) );
  XNOR2_X1 U731 ( .A(n660), .B(n659), .ZN(n661) );
  NAND2_X1 U732 ( .A1(n662), .A2(n661), .ZN(n673) );
  NAND2_X1 U733 ( .A1(n673), .A2(G286), .ZN(n668) );
  NOR2_X1 U734 ( .A1(G1971), .A2(n707), .ZN(n665) );
  NOR2_X1 U735 ( .A1(G2090), .A2(n663), .ZN(n664) );
  NOR2_X1 U736 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U737 ( .A1(G303), .A2(n666), .ZN(n667) );
  NAND2_X1 U738 ( .A1(n668), .A2(n667), .ZN(n670) );
  NOR2_X1 U739 ( .A1(n674), .A2(n519), .ZN(n677) );
  NAND2_X1 U740 ( .A1(n675), .A2(G8), .ZN(n676) );
  NAND2_X1 U741 ( .A1(n677), .A2(n676), .ZN(n697) );
  INV_X1 U742 ( .A(KEYINPUT33), .ZN(n678) );
  NAND2_X1 U743 ( .A1(G1976), .A2(G288), .ZN(n1015) );
  AND2_X1 U744 ( .A1(n678), .A2(n1015), .ZN(n683) );
  AND2_X1 U745 ( .A1(n697), .A2(n683), .ZN(n679) );
  NAND2_X1 U746 ( .A1(n696), .A2(n679), .ZN(n692) );
  NOR2_X1 U747 ( .A1(G1976), .A2(G288), .ZN(n685) );
  INV_X1 U748 ( .A(n707), .ZN(n681) );
  NAND2_X1 U749 ( .A1(n685), .A2(n681), .ZN(n680) );
  NAND2_X1 U750 ( .A1(n680), .A2(KEYINPUT33), .ZN(n688) );
  INV_X1 U751 ( .A(n688), .ZN(n682) );
  INV_X1 U752 ( .A(n683), .ZN(n687) );
  NOR2_X1 U753 ( .A1(G303), .A2(G1971), .ZN(n684) );
  NOR2_X1 U754 ( .A1(n685), .A2(n684), .ZN(n1016) );
  XNOR2_X1 U755 ( .A(KEYINPUT106), .B(n1016), .ZN(n686) );
  OR2_X1 U756 ( .A1(n687), .A2(n686), .ZN(n689) );
  AND2_X1 U757 ( .A1(n689), .A2(n688), .ZN(n690) );
  OR2_X1 U758 ( .A1(n520), .A2(n690), .ZN(n691) );
  NAND2_X1 U759 ( .A1(n692), .A2(n691), .ZN(n694) );
  XNOR2_X1 U760 ( .A(n694), .B(n693), .ZN(n695) );
  XOR2_X1 U761 ( .A(G1981), .B(G305), .Z(n1007) );
  NAND2_X1 U762 ( .A1(n695), .A2(n1007), .ZN(n703) );
  NAND2_X1 U763 ( .A1(n697), .A2(n696), .ZN(n700) );
  NOR2_X1 U764 ( .A1(G2090), .A2(G303), .ZN(n698) );
  NAND2_X1 U765 ( .A1(G8), .A2(n698), .ZN(n699) );
  NAND2_X1 U766 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U767 ( .A1(n701), .A2(n707), .ZN(n702) );
  NAND2_X1 U768 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U769 ( .A(n704), .B(KEYINPUT108), .ZN(n709) );
  NOR2_X1 U770 ( .A1(G1981), .A2(G305), .ZN(n705) );
  XOR2_X1 U771 ( .A(n705), .B(KEYINPUT24), .Z(n706) );
  NOR2_X1 U772 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U773 ( .A1(n709), .A2(n708), .ZN(n711) );
  XNOR2_X1 U774 ( .A(n711), .B(n710), .ZN(n752) );
  NAND2_X1 U775 ( .A1(G107), .A2(n894), .ZN(n712) );
  XNOR2_X1 U776 ( .A(n712), .B(KEYINPUT94), .ZN(n722) );
  NAND2_X1 U777 ( .A1(G119), .A2(n714), .ZN(n716) );
  NAND2_X1 U778 ( .A1(G95), .A2(n890), .ZN(n715) );
  NAND2_X1 U779 ( .A1(n716), .A2(n715), .ZN(n720) );
  BUF_X1 U780 ( .A(n717), .Z(n891) );
  NAND2_X1 U781 ( .A1(G131), .A2(n891), .ZN(n718) );
  XNOR2_X1 U782 ( .A(KEYINPUT95), .B(n718), .ZN(n719) );
  NOR2_X1 U783 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U784 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U785 ( .A(KEYINPUT96), .B(n723), .ZN(n873) );
  AND2_X1 U786 ( .A1(G1991), .A2(n873), .ZN(n733) );
  NAND2_X1 U787 ( .A1(G105), .A2(n890), .ZN(n724) );
  XNOR2_X1 U788 ( .A(n724), .B(KEYINPUT38), .ZN(n731) );
  NAND2_X1 U789 ( .A1(G129), .A2(n714), .ZN(n726) );
  NAND2_X1 U790 ( .A1(G141), .A2(n891), .ZN(n725) );
  NAND2_X1 U791 ( .A1(n726), .A2(n725), .ZN(n729) );
  NAND2_X1 U792 ( .A1(G117), .A2(n894), .ZN(n727) );
  XNOR2_X1 U793 ( .A(KEYINPUT97), .B(n727), .ZN(n728) );
  NOR2_X1 U794 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U795 ( .A1(n731), .A2(n730), .ZN(n885) );
  AND2_X1 U796 ( .A1(n885), .A2(G1996), .ZN(n732) );
  NOR2_X1 U797 ( .A1(n733), .A2(n732), .ZN(n989) );
  INV_X1 U798 ( .A(n734), .ZN(n735) );
  NOR2_X1 U799 ( .A1(n736), .A2(n735), .ZN(n767) );
  INV_X1 U800 ( .A(n767), .ZN(n737) );
  NOR2_X1 U801 ( .A1(n989), .A2(n737), .ZN(n758) );
  INV_X1 U802 ( .A(n758), .ZN(n750) );
  XNOR2_X1 U803 ( .A(G2067), .B(KEYINPUT37), .ZN(n765) );
  NAND2_X1 U804 ( .A1(n890), .A2(G104), .ZN(n738) );
  XOR2_X1 U805 ( .A(KEYINPUT91), .B(n738), .Z(n740) );
  NAND2_X1 U806 ( .A1(G140), .A2(n891), .ZN(n739) );
  NAND2_X1 U807 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U808 ( .A(KEYINPUT34), .B(n741), .ZN(n747) );
  NAND2_X1 U809 ( .A1(G128), .A2(n714), .ZN(n743) );
  NAND2_X1 U810 ( .A1(G116), .A2(n894), .ZN(n742) );
  NAND2_X1 U811 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U812 ( .A(KEYINPUT92), .B(n744), .Z(n745) );
  XNOR2_X1 U813 ( .A(KEYINPUT35), .B(n745), .ZN(n746) );
  NOR2_X1 U814 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U815 ( .A(n748), .B(KEYINPUT36), .Z(n749) );
  XNOR2_X1 U816 ( .A(KEYINPUT93), .B(n749), .ZN(n901) );
  NOR2_X1 U817 ( .A1(n765), .A2(n901), .ZN(n977) );
  NAND2_X1 U818 ( .A1(n767), .A2(n977), .ZN(n763) );
  NAND2_X1 U819 ( .A1(n750), .A2(n763), .ZN(n751) );
  NOR2_X1 U820 ( .A1(n752), .A2(n751), .ZN(n755) );
  XNOR2_X1 U821 ( .A(G1986), .B(KEYINPUT90), .ZN(n753) );
  XNOR2_X1 U822 ( .A(n753), .B(G290), .ZN(n1024) );
  NAND2_X1 U823 ( .A1(n1024), .A2(n767), .ZN(n754) );
  NAND2_X1 U824 ( .A1(n755), .A2(n754), .ZN(n770) );
  XOR2_X1 U825 ( .A(KEYINPUT39), .B(KEYINPUT111), .Z(n762) );
  NOR2_X1 U826 ( .A1(G1996), .A2(n885), .ZN(n991) );
  NOR2_X1 U827 ( .A1(G1986), .A2(G290), .ZN(n756) );
  NOR2_X1 U828 ( .A1(G1991), .A2(n873), .ZN(n987) );
  NOR2_X1 U829 ( .A1(n756), .A2(n987), .ZN(n757) );
  NOR2_X1 U830 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U831 ( .A(n759), .B(KEYINPUT110), .ZN(n760) );
  NOR2_X1 U832 ( .A1(n991), .A2(n760), .ZN(n761) );
  XNOR2_X1 U833 ( .A(n762), .B(n761), .ZN(n764) );
  NAND2_X1 U834 ( .A1(n764), .A2(n763), .ZN(n766) );
  NAND2_X1 U835 ( .A1(n765), .A2(n901), .ZN(n979) );
  NAND2_X1 U836 ( .A1(n766), .A2(n979), .ZN(n768) );
  NAND2_X1 U837 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U838 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U839 ( .A(n771), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U840 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U841 ( .A1(G123), .A2(n714), .ZN(n773) );
  XNOR2_X1 U842 ( .A(n773), .B(KEYINPUT18), .ZN(n780) );
  NAND2_X1 U843 ( .A1(G99), .A2(n890), .ZN(n775) );
  NAND2_X1 U844 ( .A1(G111), .A2(n894), .ZN(n774) );
  NAND2_X1 U845 ( .A1(n775), .A2(n774), .ZN(n778) );
  NAND2_X1 U846 ( .A1(G135), .A2(n891), .ZN(n776) );
  XNOR2_X1 U847 ( .A(KEYINPUT81), .B(n776), .ZN(n777) );
  NOR2_X1 U848 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U849 ( .A1(n780), .A2(n779), .ZN(n984) );
  XNOR2_X1 U850 ( .A(G2096), .B(n984), .ZN(n781) );
  OR2_X1 U851 ( .A1(G2100), .A2(n781), .ZN(G156) );
  INV_X1 U852 ( .A(G108), .ZN(G238) );
  INV_X1 U853 ( .A(G132), .ZN(G219) );
  NAND2_X1 U854 ( .A1(G7), .A2(G661), .ZN(n782) );
  XNOR2_X1 U855 ( .A(n782), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U856 ( .A(KEYINPUT74), .B(KEYINPUT11), .Z(n784) );
  XNOR2_X1 U857 ( .A(G223), .B(KEYINPUT73), .ZN(n837) );
  NAND2_X1 U858 ( .A1(G567), .A2(n837), .ZN(n783) );
  XNOR2_X1 U859 ( .A(n784), .B(n783), .ZN(G234) );
  INV_X1 U860 ( .A(G860), .ZN(n790) );
  OR2_X1 U861 ( .A1(n1006), .A2(n790), .ZN(G153) );
  INV_X1 U862 ( .A(G171), .ZN(G301) );
  NAND2_X1 U863 ( .A1(G301), .A2(G868), .ZN(n786) );
  INV_X1 U864 ( .A(n1022), .ZN(n905) );
  INV_X1 U865 ( .A(G868), .ZN(n787) );
  NAND2_X1 U866 ( .A1(n905), .A2(n787), .ZN(n785) );
  NAND2_X1 U867 ( .A1(n786), .A2(n785), .ZN(G284) );
  NOR2_X1 U868 ( .A1(G286), .A2(n787), .ZN(n789) );
  NOR2_X1 U869 ( .A1(G868), .A2(G299), .ZN(n788) );
  NOR2_X1 U870 ( .A1(n789), .A2(n788), .ZN(G297) );
  NAND2_X1 U871 ( .A1(G559), .A2(n790), .ZN(n791) );
  XNOR2_X1 U872 ( .A(KEYINPUT80), .B(n791), .ZN(n792) );
  NAND2_X1 U873 ( .A1(n792), .A2(n1022), .ZN(n793) );
  XNOR2_X1 U874 ( .A(KEYINPUT16), .B(n793), .ZN(G148) );
  NOR2_X1 U875 ( .A1(G868), .A2(n1006), .ZN(n796) );
  NAND2_X1 U876 ( .A1(n1022), .A2(G868), .ZN(n794) );
  NOR2_X1 U877 ( .A1(G559), .A2(n794), .ZN(n795) );
  NOR2_X1 U878 ( .A1(n796), .A2(n795), .ZN(G282) );
  NAND2_X1 U879 ( .A1(G559), .A2(n1022), .ZN(n797) );
  XNOR2_X1 U880 ( .A(n797), .B(n1006), .ZN(n817) );
  NOR2_X1 U881 ( .A1(n817), .A2(G860), .ZN(n809) );
  NAND2_X1 U882 ( .A1(G93), .A2(n798), .ZN(n801) );
  NAND2_X1 U883 ( .A1(G55), .A2(n799), .ZN(n800) );
  NAND2_X1 U884 ( .A1(n801), .A2(n800), .ZN(n808) );
  NAND2_X1 U885 ( .A1(G67), .A2(n802), .ZN(n803) );
  XNOR2_X1 U886 ( .A(n803), .B(KEYINPUT82), .ZN(n806) );
  NAND2_X1 U887 ( .A1(G80), .A2(n804), .ZN(n805) );
  NAND2_X1 U888 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U889 ( .A1(n808), .A2(n807), .ZN(n812) );
  XNOR2_X1 U890 ( .A(n809), .B(n812), .ZN(G145) );
  NOR2_X1 U891 ( .A1(G868), .A2(n812), .ZN(n810) );
  XNOR2_X1 U892 ( .A(n810), .B(KEYINPUT85), .ZN(n820) );
  XNOR2_X1 U893 ( .A(KEYINPUT19), .B(G290), .ZN(n811) );
  XNOR2_X1 U894 ( .A(n811), .B(G288), .ZN(n813) );
  XOR2_X1 U895 ( .A(n813), .B(n812), .Z(n815) );
  XNOR2_X1 U896 ( .A(n1012), .B(G303), .ZN(n814) );
  XNOR2_X1 U897 ( .A(n815), .B(n814), .ZN(n816) );
  XNOR2_X1 U898 ( .A(n816), .B(G305), .ZN(n907) );
  XNOR2_X1 U899 ( .A(n907), .B(n817), .ZN(n818) );
  NAND2_X1 U900 ( .A1(G868), .A2(n818), .ZN(n819) );
  NAND2_X1 U901 ( .A1(n820), .A2(n819), .ZN(G295) );
  NAND2_X1 U902 ( .A1(G2084), .A2(G2078), .ZN(n821) );
  XOR2_X1 U903 ( .A(KEYINPUT20), .B(n821), .Z(n822) );
  NAND2_X1 U904 ( .A1(G2090), .A2(n822), .ZN(n823) );
  XNOR2_X1 U905 ( .A(KEYINPUT21), .B(n823), .ZN(n824) );
  NAND2_X1 U906 ( .A1(n824), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U907 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U908 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  NOR2_X1 U909 ( .A1(G220), .A2(G219), .ZN(n825) );
  XOR2_X1 U910 ( .A(KEYINPUT22), .B(n825), .Z(n826) );
  NOR2_X1 U911 ( .A1(G218), .A2(n826), .ZN(n827) );
  NAND2_X1 U912 ( .A1(G96), .A2(n827), .ZN(n842) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n842), .ZN(n833) );
  NAND2_X1 U914 ( .A1(G69), .A2(G120), .ZN(n828) );
  XNOR2_X1 U915 ( .A(KEYINPUT86), .B(n828), .ZN(n829) );
  NOR2_X1 U916 ( .A1(G238), .A2(n829), .ZN(n830) );
  NAND2_X1 U917 ( .A1(G57), .A2(n830), .ZN(n841) );
  NAND2_X1 U918 ( .A1(G567), .A2(n841), .ZN(n831) );
  XOR2_X1 U919 ( .A(KEYINPUT87), .B(n831), .Z(n832) );
  NAND2_X1 U920 ( .A1(n833), .A2(n832), .ZN(n834) );
  XOR2_X1 U921 ( .A(KEYINPUT88), .B(n834), .Z(G319) );
  INV_X1 U922 ( .A(G319), .ZN(n836) );
  NAND2_X1 U923 ( .A1(G661), .A2(G483), .ZN(n835) );
  NOR2_X1 U924 ( .A1(n836), .A2(n835), .ZN(n840) );
  NAND2_X1 U925 ( .A1(n840), .A2(G36), .ZN(G176) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U928 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U930 ( .A1(n840), .A2(n839), .ZN(G188) );
  XOR2_X1 U931 ( .A(G120), .B(KEYINPUT112), .Z(G236) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  INV_X1 U934 ( .A(G69), .ZN(G235) );
  NOR2_X1 U935 ( .A1(n842), .A2(n841), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  XOR2_X1 U937 ( .A(G2474), .B(G1961), .Z(n844) );
  XNOR2_X1 U938 ( .A(G1996), .B(G1991), .ZN(n843) );
  XNOR2_X1 U939 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U940 ( .A(n845), .B(KEYINPUT114), .Z(n847) );
  XNOR2_X1 U941 ( .A(G1976), .B(G1971), .ZN(n846) );
  XNOR2_X1 U942 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U943 ( .A(G1956), .B(G1966), .Z(n849) );
  XNOR2_X1 U944 ( .A(G1986), .B(G1981), .ZN(n848) );
  XNOR2_X1 U945 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U946 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U947 ( .A(KEYINPUT41), .B(KEYINPUT113), .ZN(n852) );
  XNOR2_X1 U948 ( .A(n853), .B(n852), .ZN(G229) );
  XOR2_X1 U949 ( .A(G2100), .B(G2096), .Z(n855) );
  XNOR2_X1 U950 ( .A(KEYINPUT42), .B(G2678), .ZN(n854) );
  XNOR2_X1 U951 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U952 ( .A(KEYINPUT43), .B(G2090), .Z(n857) );
  XNOR2_X1 U953 ( .A(G2067), .B(G2072), .ZN(n856) );
  XNOR2_X1 U954 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U955 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U956 ( .A(G2084), .B(G2078), .ZN(n860) );
  XNOR2_X1 U957 ( .A(n861), .B(n860), .ZN(G227) );
  NAND2_X1 U958 ( .A1(G124), .A2(n714), .ZN(n862) );
  XOR2_X1 U959 ( .A(KEYINPUT115), .B(n862), .Z(n863) );
  XNOR2_X1 U960 ( .A(n863), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U961 ( .A1(G112), .A2(n894), .ZN(n864) );
  NAND2_X1 U962 ( .A1(n865), .A2(n864), .ZN(n869) );
  NAND2_X1 U963 ( .A1(G100), .A2(n890), .ZN(n867) );
  NAND2_X1 U964 ( .A1(G136), .A2(n891), .ZN(n866) );
  NAND2_X1 U965 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U966 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U967 ( .A(KEYINPUT116), .B(n870), .ZN(G162) );
  XOR2_X1 U968 ( .A(KEYINPUT118), .B(KEYINPUT46), .Z(n872) );
  XNOR2_X1 U969 ( .A(G164), .B(KEYINPUT48), .ZN(n871) );
  XNOR2_X1 U970 ( .A(n872), .B(n871), .ZN(n889) );
  XNOR2_X1 U971 ( .A(n873), .B(G162), .ZN(n874) );
  XNOR2_X1 U972 ( .A(n874), .B(n984), .ZN(n884) );
  NAND2_X1 U973 ( .A1(G130), .A2(n714), .ZN(n876) );
  NAND2_X1 U974 ( .A1(G118), .A2(n894), .ZN(n875) );
  NAND2_X1 U975 ( .A1(n876), .A2(n875), .ZN(n882) );
  NAND2_X1 U976 ( .A1(G106), .A2(n890), .ZN(n878) );
  NAND2_X1 U977 ( .A1(G142), .A2(n891), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U979 ( .A(KEYINPUT45), .B(n879), .ZN(n880) );
  XNOR2_X1 U980 ( .A(KEYINPUT117), .B(n880), .ZN(n881) );
  NOR2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U982 ( .A(n884), .B(n883), .Z(n887) );
  XOR2_X1 U983 ( .A(G160), .B(n885), .Z(n886) );
  XNOR2_X1 U984 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U985 ( .A(n889), .B(n888), .ZN(n903) );
  NAND2_X1 U986 ( .A1(G103), .A2(n890), .ZN(n893) );
  NAND2_X1 U987 ( .A1(G139), .A2(n891), .ZN(n892) );
  NAND2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n899) );
  NAND2_X1 U989 ( .A1(G127), .A2(n714), .ZN(n896) );
  NAND2_X1 U990 ( .A1(G115), .A2(n894), .ZN(n895) );
  NAND2_X1 U991 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U992 ( .A(KEYINPUT47), .B(n897), .Z(n898) );
  NOR2_X1 U993 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U994 ( .A(KEYINPUT119), .B(n900), .Z(n980) );
  XNOR2_X1 U995 ( .A(n901), .B(n980), .ZN(n902) );
  XNOR2_X1 U996 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U997 ( .A1(G37), .A2(n904), .ZN(G395) );
  XNOR2_X1 U998 ( .A(G286), .B(n905), .ZN(n906) );
  XNOR2_X1 U999 ( .A(n906), .B(n1006), .ZN(n909) );
  XOR2_X1 U1000 ( .A(G301), .B(n907), .Z(n908) );
  XNOR2_X1 U1001 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n910), .ZN(G397) );
  XOR2_X1 U1003 ( .A(G2451), .B(G2430), .Z(n912) );
  XNOR2_X1 U1004 ( .A(G2438), .B(G2443), .ZN(n911) );
  XNOR2_X1 U1005 ( .A(n912), .B(n911), .ZN(n918) );
  XOR2_X1 U1006 ( .A(G2435), .B(G2454), .Z(n914) );
  XNOR2_X1 U1007 ( .A(G1341), .B(G1348), .ZN(n913) );
  XNOR2_X1 U1008 ( .A(n914), .B(n913), .ZN(n916) );
  XOR2_X1 U1009 ( .A(G2446), .B(G2427), .Z(n915) );
  XNOR2_X1 U1010 ( .A(n916), .B(n915), .ZN(n917) );
  XOR2_X1 U1011 ( .A(n918), .B(n917), .Z(n919) );
  NAND2_X1 U1012 ( .A1(G14), .A2(n919), .ZN(n925) );
  NAND2_X1 U1013 ( .A1(n925), .A2(G319), .ZN(n922) );
  NOR2_X1 U1014 ( .A1(G229), .A2(G227), .ZN(n920) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n920), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(n922), .A2(n921), .ZN(n924) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1018 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G57), .ZN(G237) );
  INV_X1 U1021 ( .A(n925), .ZN(G401) );
  XOR2_X1 U1022 ( .A(G1981), .B(G6), .Z(n928) );
  XNOR2_X1 U1023 ( .A(n926), .B(G20), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n934) );
  XOR2_X1 U1025 ( .A(G1341), .B(G19), .Z(n932) );
  XOR2_X1 U1026 ( .A(KEYINPUT59), .B(G4), .Z(n929) );
  XNOR2_X1 U1027 ( .A(KEYINPUT125), .B(n929), .ZN(n930) );
  XNOR2_X1 U1028 ( .A(n930), .B(G1348), .ZN(n931) );
  NAND2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1031 ( .A(KEYINPUT60), .B(n935), .ZN(n939) );
  XNOR2_X1 U1032 ( .A(G1966), .B(G21), .ZN(n937) );
  XNOR2_X1 U1033 ( .A(G1961), .B(G5), .ZN(n936) );
  NOR2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(KEYINPUT126), .B(n940), .ZN(n948) );
  XOR2_X1 U1037 ( .A(G1986), .B(G24), .Z(n944) );
  XNOR2_X1 U1038 ( .A(G1976), .B(G23), .ZN(n942) );
  XNOR2_X1 U1039 ( .A(G1971), .B(G22), .ZN(n941) );
  NOR2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1042 ( .A(KEYINPUT127), .B(n945), .Z(n946) );
  XNOR2_X1 U1043 ( .A(KEYINPUT58), .B(n946), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1045 ( .A(KEYINPUT61), .B(n949), .Z(n951) );
  XNOR2_X1 U1046 ( .A(G16), .B(KEYINPUT124), .ZN(n950) );
  NOR2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n976) );
  INV_X1 U1048 ( .A(KEYINPUT55), .ZN(n1000) );
  XNOR2_X1 U1049 ( .A(G2090), .B(G35), .ZN(n967) );
  XOR2_X1 U1050 ( .A(G2072), .B(G33), .Z(n952) );
  NAND2_X1 U1051 ( .A1(n952), .A2(G28), .ZN(n964) );
  XNOR2_X1 U1052 ( .A(n953), .B(G27), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(KEYINPUT120), .B(G32), .ZN(n955) );
  XNOR2_X1 U1054 ( .A(n955), .B(n954), .ZN(n956) );
  NAND2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1056 ( .A(n958), .B(KEYINPUT121), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(G2067), .B(G26), .ZN(n960) );
  XNOR2_X1 U1058 ( .A(G1991), .B(G25), .ZN(n959) );
  NOR2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1062 ( .A(KEYINPUT53), .B(n965), .ZN(n966) );
  NOR2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n970) );
  XOR2_X1 U1064 ( .A(G2084), .B(G34), .Z(n968) );
  XNOR2_X1 U1065 ( .A(KEYINPUT54), .B(n968), .ZN(n969) );
  NAND2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1067 ( .A(n1000), .B(n971), .ZN(n973) );
  INV_X1 U1068 ( .A(G29), .ZN(n972) );
  NAND2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1070 ( .A1(G11), .A2(n974), .ZN(n975) );
  NOR2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n1004) );
  INV_X1 U1072 ( .A(n977), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n998) );
  XOR2_X1 U1074 ( .A(G2072), .B(n980), .Z(n982) );
  XOR2_X1 U1075 ( .A(G164), .B(G2078), .Z(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(KEYINPUT50), .B(n983), .ZN(n996) );
  XNOR2_X1 U1078 ( .A(G160), .B(G2084), .ZN(n985) );
  NAND2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n994) );
  XOR2_X1 U1082 ( .A(G2090), .B(G162), .Z(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1084 ( .A(n992), .B(KEYINPUT51), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(KEYINPUT52), .B(n999), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1090 ( .A1(n1002), .A2(G29), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1032) );
  XOR2_X1 U1092 ( .A(KEYINPUT56), .B(G16), .Z(n1030) );
  XOR2_X1 U1093 ( .A(G1341), .B(KEYINPUT123), .Z(n1005) );
  XNOR2_X1 U1094 ( .A(n1006), .B(n1005), .ZN(n1028) );
  XNOR2_X1 U1095 ( .A(G1961), .B(G171), .ZN(n1011) );
  XNOR2_X1 U1096 ( .A(G1966), .B(G168), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(n1009), .B(KEYINPUT57), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1021) );
  XNOR2_X1 U1100 ( .A(n1012), .B(G1956), .ZN(n1014) );
  NAND2_X1 U1101 ( .A1(G1971), .A2(G303), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1018) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1105 ( .A(KEYINPUT122), .B(n1019), .Z(n1020) );
  NOR2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1026) );
  XOR2_X1 U1107 ( .A(G1348), .B(n1022), .Z(n1023) );
  NOR2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1109 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1110 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1111 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1112 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1113 ( .A(n1033), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
  INV_X1 U1115 ( .A(G303), .ZN(G166) );
endmodule

